module BBGSharePredictorImp_BSD_c_NutShell(
    input [31:0] pc,
    input [31:0] train_pc,
    input  train_taken,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    input [15:0] train_ghr_rdata,
    output  taken,
    output  pht_wdata,
    output [8:0] pht_raddr,
    output [8:0] pht_waddr,
    output  ghr_wdata
);
wire [98:0] io_x;
wire [20:0] io_y;
assign io_x = { pc, train_pc, train_taken, pht_rdata, ghr_rdata, train_ghr_rdata };
assign { taken, pht_wdata, pht_raddr, pht_waddr, ghr_wdata } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[33] ? _GEN1 : _GEN0;
assign io_y[20] = _GEN2;
wire  _GEN3 = 1'b0;
wire  _GEN4 = 1'b1;
wire  _GEN5 = io_x[34] ? _GEN4 : _GEN3;
assign io_y[19] = _GEN5;
wire  _GEN6 = 1'b0;
wire  _GEN7 = 1'b1;
wire  _GEN8 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN9 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN10 = io_x[27] ? _GEN9 : _GEN8;
wire  _GEN11 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN12 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN13 = io_x[27] ? _GEN12 : _GEN11;
wire  _GEN14 = io_x[31] ? _GEN13 : _GEN10;
wire  _GEN15 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN16 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN17 = io_x[27] ? _GEN16 : _GEN15;
wire  _GEN18 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN19 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN20 = io_x[27] ? _GEN19 : _GEN18;
wire  _GEN21 = io_x[31] ? _GEN20 : _GEN17;
wire  _GEN22 = io_x[19] ? _GEN21 : _GEN14;
wire  _GEN23 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN24 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN25 = io_x[27] ? _GEN24 : _GEN23;
wire  _GEN26 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN27 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN28 = io_x[27] ? _GEN27 : _GEN26;
wire  _GEN29 = io_x[31] ? _GEN28 : _GEN25;
wire  _GEN30 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN31 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN32 = io_x[27] ? _GEN31 : _GEN30;
wire  _GEN33 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN34 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN35 = io_x[27] ? _GEN34 : _GEN33;
wire  _GEN36 = io_x[31] ? _GEN35 : _GEN32;
wire  _GEN37 = io_x[19] ? _GEN36 : _GEN29;
wire  _GEN38 = io_x[23] ? _GEN37 : _GEN22;
wire  _GEN39 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN40 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN41 = io_x[27] ? _GEN40 : _GEN39;
wire  _GEN42 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN43 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN44 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN45 = io_x[31] ? _GEN44 : _GEN41;
wire  _GEN46 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN47 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN48 = io_x[27] ? _GEN47 : _GEN46;
wire  _GEN49 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN50 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN51 = io_x[27] ? _GEN50 : _GEN49;
wire  _GEN52 = io_x[31] ? _GEN51 : _GEN48;
wire  _GEN53 = io_x[19] ? _GEN52 : _GEN45;
wire  _GEN54 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN55 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN56 = io_x[27] ? _GEN55 : _GEN54;
wire  _GEN57 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN58 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN59 = io_x[27] ? _GEN58 : _GEN57;
wire  _GEN60 = io_x[31] ? _GEN59 : _GEN56;
wire  _GEN61 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN62 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN63 = io_x[27] ? _GEN62 : _GEN61;
wire  _GEN64 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN65 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN66 = io_x[27] ? _GEN65 : _GEN64;
wire  _GEN67 = io_x[31] ? _GEN66 : _GEN63;
wire  _GEN68 = io_x[19] ? _GEN67 : _GEN60;
wire  _GEN69 = io_x[23] ? _GEN68 : _GEN53;
wire  _GEN70 = io_x[45] ? _GEN69 : _GEN38;
assign io_y[18] = _GEN70;
wire  _GEN71 = 1'b0;
wire  _GEN72 = 1'b1;
wire  _GEN73 = io_x[26] ? _GEN72 : _GEN71;
wire  _GEN74 = io_x[26] ? _GEN71 : _GEN72;
wire  _GEN75 = io_x[30] ? _GEN74 : _GEN73;
wire  _GEN76 = io_x[26] ? _GEN71 : _GEN72;
wire  _GEN77 = io_x[26] ? _GEN72 : _GEN71;
wire  _GEN78 = io_x[30] ? _GEN77 : _GEN76;
wire  _GEN79 = io_x[18] ? _GEN78 : _GEN75;
wire  _GEN80 = io_x[26] ? _GEN71 : _GEN72;
wire  _GEN81 = io_x[26] ? _GEN72 : _GEN71;
wire  _GEN82 = io_x[30] ? _GEN81 : _GEN80;
wire  _GEN83 = io_x[26] ? _GEN72 : _GEN71;
wire  _GEN84 = io_x[26] ? _GEN71 : _GEN72;
wire  _GEN85 = io_x[30] ? _GEN84 : _GEN83;
wire  _GEN86 = io_x[18] ? _GEN85 : _GEN82;
wire  _GEN87 = io_x[22] ? _GEN86 : _GEN79;
wire  _GEN88 = io_x[26] ? _GEN71 : _GEN72;
wire  _GEN89 = io_x[26] ? _GEN72 : _GEN71;
wire  _GEN90 = io_x[30] ? _GEN89 : _GEN88;
wire  _GEN91 = io_x[26] ? _GEN72 : _GEN71;
wire  _GEN92 = io_x[26] ? _GEN71 : _GEN72;
wire  _GEN93 = io_x[30] ? _GEN92 : _GEN91;
wire  _GEN94 = io_x[18] ? _GEN93 : _GEN90;
wire  _GEN95 = io_x[26] ? _GEN72 : _GEN71;
wire  _GEN96 = io_x[26] ? _GEN71 : _GEN72;
wire  _GEN97 = io_x[30] ? _GEN96 : _GEN95;
wire  _GEN98 = io_x[26] ? _GEN71 : _GEN72;
wire  _GEN99 = io_x[26] ? _GEN72 : _GEN71;
wire  _GEN100 = io_x[30] ? _GEN99 : _GEN98;
wire  _GEN101 = io_x[18] ? _GEN100 : _GEN97;
wire  _GEN102 = io_x[22] ? _GEN101 : _GEN94;
wire  _GEN103 = io_x[76] ? _GEN102 : _GEN87;
assign io_y[17] = _GEN103;
wire  _GEN104 = 1'b0;
wire  _GEN105 = 1'b1;
wire  _GEN106 = io_x[25] ? _GEN105 : _GEN104;
wire  _GEN107 = io_x[25] ? _GEN104 : _GEN105;
wire  _GEN108 = io_x[29] ? _GEN107 : _GEN106;
wire  _GEN109 = io_x[25] ? _GEN104 : _GEN105;
wire  _GEN110 = io_x[25] ? _GEN105 : _GEN104;
wire  _GEN111 = io_x[29] ? _GEN110 : _GEN109;
wire  _GEN112 = io_x[17] ? _GEN111 : _GEN108;
wire  _GEN113 = io_x[25] ? _GEN104 : _GEN105;
wire  _GEN114 = io_x[25] ? _GEN105 : _GEN104;
wire  _GEN115 = io_x[29] ? _GEN114 : _GEN113;
wire  _GEN116 = io_x[25] ? _GEN105 : _GEN104;
wire  _GEN117 = io_x[25] ? _GEN104 : _GEN105;
wire  _GEN118 = io_x[29] ? _GEN117 : _GEN116;
wire  _GEN119 = io_x[17] ? _GEN118 : _GEN115;
wire  _GEN120 = io_x[21] ? _GEN119 : _GEN112;
wire  _GEN121 = io_x[25] ? _GEN104 : _GEN105;
wire  _GEN122 = io_x[25] ? _GEN105 : _GEN104;
wire  _GEN123 = io_x[29] ? _GEN122 : _GEN121;
wire  _GEN124 = io_x[25] ? _GEN105 : _GEN104;
wire  _GEN125 = io_x[25] ? _GEN104 : _GEN105;
wire  _GEN126 = io_x[29] ? _GEN125 : _GEN124;
wire  _GEN127 = io_x[17] ? _GEN126 : _GEN123;
wire  _GEN128 = io_x[25] ? _GEN105 : _GEN104;
wire  _GEN129 = io_x[25] ? _GEN104 : _GEN105;
wire  _GEN130 = io_x[29] ? _GEN129 : _GEN128;
wire  _GEN131 = io_x[25] ? _GEN104 : _GEN105;
wire  _GEN132 = io_x[25] ? _GEN105 : _GEN104;
wire  _GEN133 = io_x[29] ? _GEN132 : _GEN131;
wire  _GEN134 = io_x[17] ? _GEN133 : _GEN130;
wire  _GEN135 = io_x[21] ? _GEN134 : _GEN127;
wire  _GEN136 = io_x[75] ? _GEN135 : _GEN120;
assign io_y[16] = _GEN136;
wire  _GEN137 = 1'b0;
wire  _GEN138 = 1'b1;
wire  _GEN139 = io_x[24] ? _GEN138 : _GEN137;
wire  _GEN140 = io_x[24] ? _GEN137 : _GEN138;
wire  _GEN141 = io_x[20] ? _GEN140 : _GEN139;
wire  _GEN142 = io_x[24] ? _GEN137 : _GEN138;
wire  _GEN143 = io_x[24] ? _GEN138 : _GEN137;
wire  _GEN144 = io_x[20] ? _GEN143 : _GEN142;
wire  _GEN145 = io_x[16] ? _GEN144 : _GEN141;
wire  _GEN146 = io_x[24] ? _GEN137 : _GEN138;
wire  _GEN147 = io_x[24] ? _GEN138 : _GEN137;
wire  _GEN148 = io_x[20] ? _GEN147 : _GEN146;
wire  _GEN149 = io_x[24] ? _GEN138 : _GEN137;
wire  _GEN150 = io_x[24] ? _GEN137 : _GEN138;
wire  _GEN151 = io_x[20] ? _GEN150 : _GEN149;
wire  _GEN152 = io_x[16] ? _GEN151 : _GEN148;
wire  _GEN153 = io_x[28] ? _GEN152 : _GEN145;
wire  _GEN154 = io_x[24] ? _GEN137 : _GEN138;
wire  _GEN155 = io_x[24] ? _GEN138 : _GEN137;
wire  _GEN156 = io_x[20] ? _GEN155 : _GEN154;
wire  _GEN157 = io_x[24] ? _GEN138 : _GEN137;
wire  _GEN158 = io_x[24] ? _GEN137 : _GEN138;
wire  _GEN159 = io_x[20] ? _GEN158 : _GEN157;
wire  _GEN160 = io_x[16] ? _GEN159 : _GEN156;
wire  _GEN161 = io_x[24] ? _GEN138 : _GEN137;
wire  _GEN162 = io_x[24] ? _GEN137 : _GEN138;
wire  _GEN163 = io_x[20] ? _GEN162 : _GEN161;
wire  _GEN164 = io_x[24] ? _GEN137 : _GEN138;
wire  _GEN165 = io_x[24] ? _GEN138 : _GEN137;
wire  _GEN166 = io_x[20] ? _GEN165 : _GEN164;
wire  _GEN167 = io_x[16] ? _GEN166 : _GEN163;
wire  _GEN168 = io_x[28] ? _GEN167 : _GEN160;
wire  _GEN169 = io_x[74] ? _GEN168 : _GEN153;
assign io_y[15] = _GEN169;
wire  _GEN170 = 1'b0;
wire  _GEN171 = 1'b1;
wire  _GEN172 = io_x[73] ? _GEN171 : _GEN170;
assign io_y[14] = _GEN172;
wire  _GEN173 = 1'b0;
wire  _GEN174 = 1'b1;
wire  _GEN175 = io_x[72] ? _GEN174 : _GEN173;
assign io_y[13] = _GEN175;
wire  _GEN176 = 1'b0;
wire  _GEN177 = 1'b1;
wire  _GEN178 = io_x[71] ? _GEN177 : _GEN176;
assign io_y[12] = _GEN178;
wire  _GEN179 = 1'b0;
wire  _GEN180 = 1'b1;
wire  _GEN181 = io_x[70] ? _GEN180 : _GEN179;
assign io_y[11] = _GEN181;
wire  _GEN182 = 1'b0;
wire  _GEN183 = 1'b1;
wire  _GEN184 = io_x[69] ? _GEN183 : _GEN182;
assign io_y[10] = _GEN184;
wire  _GEN185 = 1'b0;
wire  _GEN186 = 1'b1;
wire  _GEN187 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN188 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN189 = io_x[15] ? _GEN188 : _GEN187;
wire  _GEN190 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN191 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN192 = io_x[15] ? _GEN191 : _GEN190;
wire  _GEN193 = io_x[3] ? _GEN192 : _GEN189;
wire  _GEN194 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN195 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN196 = io_x[15] ? _GEN195 : _GEN194;
wire  _GEN197 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN198 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN199 = io_x[15] ? _GEN198 : _GEN197;
wire  _GEN200 = io_x[3] ? _GEN199 : _GEN196;
wire  _GEN201 = io_x[7] ? _GEN200 : _GEN193;
wire  _GEN202 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN203 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN204 = io_x[15] ? _GEN203 : _GEN202;
wire  _GEN205 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN206 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN207 = io_x[15] ? _GEN206 : _GEN205;
wire  _GEN208 = io_x[3] ? _GEN207 : _GEN204;
wire  _GEN209 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN210 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN211 = io_x[15] ? _GEN210 : _GEN209;
wire  _GEN212 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN213 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN214 = io_x[15] ? _GEN213 : _GEN212;
wire  _GEN215 = io_x[3] ? _GEN214 : _GEN211;
wire  _GEN216 = io_x[7] ? _GEN215 : _GEN208;
wire  _GEN217 = io_x[0] ? _GEN216 : _GEN201;
wire  _GEN218 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN219 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN220 = io_x[15] ? _GEN219 : _GEN218;
wire  _GEN221 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN222 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN223 = io_x[15] ? _GEN222 : _GEN221;
wire  _GEN224 = io_x[3] ? _GEN223 : _GEN220;
wire  _GEN225 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN226 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN227 = io_x[15] ? _GEN226 : _GEN225;
wire  _GEN228 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN229 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN230 = io_x[15] ? _GEN229 : _GEN228;
wire  _GEN231 = io_x[3] ? _GEN230 : _GEN227;
wire  _GEN232 = io_x[7] ? _GEN231 : _GEN224;
wire  _GEN233 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN234 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN235 = io_x[15] ? _GEN234 : _GEN233;
wire  _GEN236 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN237 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN238 = io_x[15] ? _GEN237 : _GEN236;
wire  _GEN239 = io_x[3] ? _GEN238 : _GEN235;
wire  _GEN240 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN241 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN242 = io_x[15] ? _GEN241 : _GEN240;
wire  _GEN243 = io_x[11] ? _GEN185 : _GEN186;
wire  _GEN244 = io_x[11] ? _GEN186 : _GEN185;
wire  _GEN245 = io_x[15] ? _GEN244 : _GEN243;
wire  _GEN246 = io_x[3] ? _GEN245 : _GEN242;
wire  _GEN247 = io_x[7] ? _GEN246 : _GEN239;
wire  _GEN248 = io_x[0] ? _GEN247 : _GEN232;
wire  _GEN249 = io_x[45] ? _GEN248 : _GEN217;
assign io_y[9] = _GEN249;
wire  _GEN250 = 1'b0;
wire  _GEN251 = 1'b1;
wire  _GEN252 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN253 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN254 = io_x[14] ? _GEN253 : _GEN252;
wire  _GEN255 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN256 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN257 = io_x[14] ? _GEN256 : _GEN255;
wire  _GEN258 = io_x[2] ? _GEN257 : _GEN254;
wire  _GEN259 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN260 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN261 = io_x[14] ? _GEN260 : _GEN259;
wire  _GEN262 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN263 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN264 = io_x[14] ? _GEN263 : _GEN262;
wire  _GEN265 = io_x[2] ? _GEN264 : _GEN261;
wire  _GEN266 = io_x[10] ? _GEN265 : _GEN258;
wire  _GEN267 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN268 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN269 = io_x[14] ? _GEN268 : _GEN267;
wire  _GEN270 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN271 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN272 = io_x[14] ? _GEN271 : _GEN270;
wire  _GEN273 = io_x[2] ? _GEN272 : _GEN269;
wire  _GEN274 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN275 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN276 = io_x[14] ? _GEN275 : _GEN274;
wire  _GEN277 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN278 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN279 = io_x[14] ? _GEN278 : _GEN277;
wire  _GEN280 = io_x[2] ? _GEN279 : _GEN276;
wire  _GEN281 = io_x[10] ? _GEN280 : _GEN273;
wire  _GEN282 = io_x[0] ? _GEN281 : _GEN266;
wire  _GEN283 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN284 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN285 = io_x[14] ? _GEN284 : _GEN283;
wire  _GEN286 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN287 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN288 = io_x[14] ? _GEN287 : _GEN286;
wire  _GEN289 = io_x[2] ? _GEN288 : _GEN285;
wire  _GEN290 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN291 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN292 = io_x[14] ? _GEN291 : _GEN290;
wire  _GEN293 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN294 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN295 = io_x[14] ? _GEN294 : _GEN293;
wire  _GEN296 = io_x[2] ? _GEN295 : _GEN292;
wire  _GEN297 = io_x[10] ? _GEN296 : _GEN289;
wire  _GEN298 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN299 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN300 = io_x[14] ? _GEN299 : _GEN298;
wire  _GEN301 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN302 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN303 = io_x[14] ? _GEN302 : _GEN301;
wire  _GEN304 = io_x[2] ? _GEN303 : _GEN300;
wire  _GEN305 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN306 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN307 = io_x[14] ? _GEN306 : _GEN305;
wire  _GEN308 = io_x[6] ? _GEN250 : _GEN251;
wire  _GEN309 = io_x[6] ? _GEN251 : _GEN250;
wire  _GEN310 = io_x[14] ? _GEN309 : _GEN308;
wire  _GEN311 = io_x[2] ? _GEN310 : _GEN307;
wire  _GEN312 = io_x[10] ? _GEN311 : _GEN304;
wire  _GEN313 = io_x[0] ? _GEN312 : _GEN297;
wire  _GEN314 = io_x[44] ? _GEN313 : _GEN282;
assign io_y[8] = _GEN314;
wire  _GEN315 = 1'b0;
wire  _GEN316 = 1'b1;
wire  _GEN317 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN318 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN319 = io_x[13] ? _GEN318 : _GEN317;
wire  _GEN320 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN321 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN322 = io_x[13] ? _GEN321 : _GEN320;
wire  _GEN323 = io_x[1] ? _GEN322 : _GEN319;
wire  _GEN324 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN325 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN326 = io_x[13] ? _GEN325 : _GEN324;
wire  _GEN327 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN328 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN329 = io_x[13] ? _GEN328 : _GEN327;
wire  _GEN330 = io_x[1] ? _GEN329 : _GEN326;
wire  _GEN331 = io_x[5] ? _GEN330 : _GEN323;
wire  _GEN332 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN333 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN334 = io_x[13] ? _GEN333 : _GEN332;
wire  _GEN335 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN336 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN337 = io_x[13] ? _GEN336 : _GEN335;
wire  _GEN338 = io_x[1] ? _GEN337 : _GEN334;
wire  _GEN339 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN340 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN341 = io_x[13] ? _GEN340 : _GEN339;
wire  _GEN342 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN343 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN344 = io_x[13] ? _GEN343 : _GEN342;
wire  _GEN345 = io_x[1] ? _GEN344 : _GEN341;
wire  _GEN346 = io_x[5] ? _GEN345 : _GEN338;
wire  _GEN347 = io_x[0] ? _GEN346 : _GEN331;
wire  _GEN348 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN349 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN350 = io_x[13] ? _GEN349 : _GEN348;
wire  _GEN351 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN352 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN353 = io_x[13] ? _GEN352 : _GEN351;
wire  _GEN354 = io_x[1] ? _GEN353 : _GEN350;
wire  _GEN355 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN356 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN357 = io_x[13] ? _GEN356 : _GEN355;
wire  _GEN358 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN359 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN360 = io_x[13] ? _GEN359 : _GEN358;
wire  _GEN361 = io_x[1] ? _GEN360 : _GEN357;
wire  _GEN362 = io_x[5] ? _GEN361 : _GEN354;
wire  _GEN363 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN364 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN365 = io_x[13] ? _GEN364 : _GEN363;
wire  _GEN366 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN367 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN368 = io_x[13] ? _GEN367 : _GEN366;
wire  _GEN369 = io_x[1] ? _GEN368 : _GEN365;
wire  _GEN370 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN371 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN372 = io_x[13] ? _GEN371 : _GEN370;
wire  _GEN373 = io_x[9] ? _GEN315 : _GEN316;
wire  _GEN374 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN375 = io_x[13] ? _GEN374 : _GEN373;
wire  _GEN376 = io_x[1] ? _GEN375 : _GEN372;
wire  _GEN377 = io_x[5] ? _GEN376 : _GEN369;
wire  _GEN378 = io_x[0] ? _GEN377 : _GEN362;
wire  _GEN379 = io_x[43] ? _GEN378 : _GEN347;
assign io_y[7] = _GEN379;
wire  _GEN380 = 1'b0;
wire  _GEN381 = 1'b1;
wire  _GEN382 = io_x[8] ? _GEN381 : _GEN380;
wire  _GEN383 = io_x[8] ? _GEN380 : _GEN381;
wire  _GEN384 = io_x[12] ? _GEN383 : _GEN382;
wire  _GEN385 = io_x[8] ? _GEN380 : _GEN381;
wire  _GEN386 = io_x[8] ? _GEN381 : _GEN380;
wire  _GEN387 = io_x[12] ? _GEN386 : _GEN385;
wire  _GEN388 = io_x[4] ? _GEN387 : _GEN384;
wire  _GEN389 = io_x[8] ? _GEN380 : _GEN381;
wire  _GEN390 = io_x[8] ? _GEN381 : _GEN380;
wire  _GEN391 = io_x[12] ? _GEN390 : _GEN389;
wire  _GEN392 = io_x[8] ? _GEN381 : _GEN380;
wire  _GEN393 = io_x[8] ? _GEN380 : _GEN381;
wire  _GEN394 = io_x[12] ? _GEN393 : _GEN392;
wire  _GEN395 = io_x[4] ? _GEN394 : _GEN391;
wire  _GEN396 = io_x[0] ? _GEN395 : _GEN388;
wire  _GEN397 = io_x[8] ? _GEN380 : _GEN381;
wire  _GEN398 = io_x[8] ? _GEN381 : _GEN380;
wire  _GEN399 = io_x[12] ? _GEN398 : _GEN397;
wire  _GEN400 = io_x[8] ? _GEN381 : _GEN380;
wire  _GEN401 = io_x[8] ? _GEN380 : _GEN381;
wire  _GEN402 = io_x[12] ? _GEN401 : _GEN400;
wire  _GEN403 = io_x[4] ? _GEN402 : _GEN399;
wire  _GEN404 = io_x[8] ? _GEN381 : _GEN380;
wire  _GEN405 = io_x[8] ? _GEN380 : _GEN381;
wire  _GEN406 = io_x[12] ? _GEN405 : _GEN404;
wire  _GEN407 = io_x[8] ? _GEN380 : _GEN381;
wire  _GEN408 = io_x[8] ? _GEN381 : _GEN380;
wire  _GEN409 = io_x[12] ? _GEN408 : _GEN407;
wire  _GEN410 = io_x[4] ? _GEN409 : _GEN406;
wire  _GEN411 = io_x[0] ? _GEN410 : _GEN403;
wire  _GEN412 = io_x[42] ? _GEN411 : _GEN396;
assign io_y[6] = _GEN412;
wire  _GEN413 = 1'b0;
wire  _GEN414 = 1'b1;
wire  _GEN415 = io_x[41] ? _GEN414 : _GEN413;
assign io_y[5] = _GEN415;
wire  _GEN416 = 1'b0;
wire  _GEN417 = 1'b1;
wire  _GEN418 = io_x[40] ? _GEN417 : _GEN416;
assign io_y[4] = _GEN418;
wire  _GEN419 = 1'b0;
wire  _GEN420 = 1'b1;
wire  _GEN421 = io_x[39] ? _GEN420 : _GEN419;
assign io_y[3] = _GEN421;
wire  _GEN422 = 1'b0;
wire  _GEN423 = 1'b1;
wire  _GEN424 = io_x[38] ? _GEN423 : _GEN422;
assign io_y[2] = _GEN424;
wire  _GEN425 = 1'b0;
wire  _GEN426 = 1'b1;
wire  _GEN427 = io_x[37] ? _GEN426 : _GEN425;
assign io_y[1] = _GEN427;
wire  _GEN428 = 1'b0;
wire  _GEN429 = 1'b1;
wire  _GEN430 = io_x[34] ? _GEN429 : _GEN428;
assign io_y[0] = _GEN430;
endmodule
