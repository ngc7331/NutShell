module BBGSharePredictorImp_BSD_c_NutShell_split(
    input [31:0] pc,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    output  taken,
    output [8:0] pht_raddr,
    input [31:0] train_pc,
    input  train_taken,
    input [15:0] train_ghr_rdata,
    output  pht_wdata,
    output [8:0] pht_waddr,
    output  ghr_wdata
);

BBGSharePredictorImp_BSD_NutShell_pred _pred(
    .pc        (pc),
    .pht_rdata (pht_rdata),
    .ghr_rdata (ghr_rdata),
    .taken     (taken),
    .pht_raddr (pht_raddr)
);

BBGSharePredictorImp_BSD_NutShell_train _train(
    .train_pc        (train_pc),
    .train_taken     (train_taken),
    .train_ghr_rdata (train_ghr_rdata),
    .pht_wdata       (pht_wdata),
    .pht_waddr       (pht_waddr),
    .ghr_wdata       (ghr_wdata)
);
endmodule
module BBGSharePredictorImp_BSD_NutShell_pred(
    input [31:0] pc,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    output  taken,
    output [8:0] pht_raddr
);
wire [49:0] io_x;
wire [9:0] io_y;
assign io_x = { pc, pht_rdata, ghr_rdata };
assign { taken, pht_raddr } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[17] ? _GEN1 : _GEN0;
assign io_y[9] = _GEN2;
wire  _GEN3 = 1'b0;
wire  _GEN4 = 1'b1;
wire  _GEN5 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN6 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN7 = io_x[15] ? _GEN6 : _GEN5;
wire  _GEN8 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN9 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN10 = io_x[15] ? _GEN9 : _GEN8;
wire  _GEN11 = io_x[3] ? _GEN10 : _GEN7;
wire  _GEN12 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN13 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN14 = io_x[15] ? _GEN13 : _GEN12;
wire  _GEN15 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN16 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN17 = io_x[15] ? _GEN16 : _GEN15;
wire  _GEN18 = io_x[3] ? _GEN17 : _GEN14;
wire  _GEN19 = io_x[7] ? _GEN18 : _GEN11;
wire  _GEN20 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN21 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN22 = io_x[15] ? _GEN21 : _GEN20;
wire  _GEN23 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN24 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN25 = io_x[15] ? _GEN24 : _GEN23;
wire  _GEN26 = io_x[3] ? _GEN25 : _GEN22;
wire  _GEN27 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN28 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN29 = io_x[15] ? _GEN28 : _GEN27;
wire  _GEN30 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN31 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN32 = io_x[15] ? _GEN31 : _GEN30;
wire  _GEN33 = io_x[3] ? _GEN32 : _GEN29;
wire  _GEN34 = io_x[7] ? _GEN33 : _GEN26;
wire  _GEN35 = io_x[28] ? _GEN34 : _GEN19;
assign io_y[8] = _GEN35;
wire  _GEN36 = 1'b0;
wire  _GEN37 = 1'b1;
wire  _GEN38 = io_x[10] ? _GEN37 : _GEN36;
wire  _GEN39 = io_x[10] ? _GEN36 : _GEN37;
wire  _GEN40 = io_x[14] ? _GEN39 : _GEN38;
wire  _GEN41 = io_x[10] ? _GEN36 : _GEN37;
wire  _GEN42 = io_x[10] ? _GEN37 : _GEN36;
wire  _GEN43 = io_x[14] ? _GEN42 : _GEN41;
wire  _GEN44 = io_x[2] ? _GEN43 : _GEN40;
wire  _GEN45 = io_x[10] ? _GEN36 : _GEN37;
wire  _GEN46 = io_x[10] ? _GEN37 : _GEN36;
wire  _GEN47 = io_x[14] ? _GEN46 : _GEN45;
wire  _GEN48 = io_x[10] ? _GEN37 : _GEN36;
wire  _GEN49 = io_x[10] ? _GEN36 : _GEN37;
wire  _GEN50 = io_x[14] ? _GEN49 : _GEN48;
wire  _GEN51 = io_x[2] ? _GEN50 : _GEN47;
wire  _GEN52 = io_x[6] ? _GEN51 : _GEN44;
wire  _GEN53 = io_x[10] ? _GEN36 : _GEN37;
wire  _GEN54 = io_x[10] ? _GEN37 : _GEN36;
wire  _GEN55 = io_x[14] ? _GEN54 : _GEN53;
wire  _GEN56 = io_x[10] ? _GEN37 : _GEN36;
wire  _GEN57 = io_x[10] ? _GEN36 : _GEN37;
wire  _GEN58 = io_x[14] ? _GEN57 : _GEN56;
wire  _GEN59 = io_x[2] ? _GEN58 : _GEN55;
wire  _GEN60 = io_x[10] ? _GEN37 : _GEN36;
wire  _GEN61 = io_x[10] ? _GEN36 : _GEN37;
wire  _GEN62 = io_x[14] ? _GEN61 : _GEN60;
wire  _GEN63 = io_x[10] ? _GEN36 : _GEN37;
wire  _GEN64 = io_x[10] ? _GEN37 : _GEN36;
wire  _GEN65 = io_x[14] ? _GEN64 : _GEN63;
wire  _GEN66 = io_x[2] ? _GEN65 : _GEN62;
wire  _GEN67 = io_x[6] ? _GEN66 : _GEN59;
wire  _GEN68 = io_x[27] ? _GEN67 : _GEN52;
assign io_y[7] = _GEN68;
wire  _GEN69 = 1'b0;
wire  _GEN70 = 1'b1;
wire  _GEN71 = io_x[9] ? _GEN70 : _GEN69;
wire  _GEN72 = io_x[9] ? _GEN69 : _GEN70;
wire  _GEN73 = io_x[13] ? _GEN72 : _GEN71;
wire  _GEN74 = io_x[9] ? _GEN69 : _GEN70;
wire  _GEN75 = io_x[9] ? _GEN70 : _GEN69;
wire  _GEN76 = io_x[13] ? _GEN75 : _GEN74;
wire  _GEN77 = io_x[1] ? _GEN76 : _GEN73;
wire  _GEN78 = io_x[9] ? _GEN69 : _GEN70;
wire  _GEN79 = io_x[9] ? _GEN70 : _GEN69;
wire  _GEN80 = io_x[13] ? _GEN79 : _GEN78;
wire  _GEN81 = io_x[9] ? _GEN70 : _GEN69;
wire  _GEN82 = io_x[9] ? _GEN69 : _GEN70;
wire  _GEN83 = io_x[13] ? _GEN82 : _GEN81;
wire  _GEN84 = io_x[1] ? _GEN83 : _GEN80;
wire  _GEN85 = io_x[5] ? _GEN84 : _GEN77;
wire  _GEN86 = io_x[9] ? _GEN69 : _GEN70;
wire  _GEN87 = io_x[9] ? _GEN70 : _GEN69;
wire  _GEN88 = io_x[13] ? _GEN87 : _GEN86;
wire  _GEN89 = io_x[9] ? _GEN70 : _GEN69;
wire  _GEN90 = io_x[9] ? _GEN69 : _GEN70;
wire  _GEN91 = io_x[13] ? _GEN90 : _GEN89;
wire  _GEN92 = io_x[1] ? _GEN91 : _GEN88;
wire  _GEN93 = io_x[9] ? _GEN70 : _GEN69;
wire  _GEN94 = io_x[9] ? _GEN69 : _GEN70;
wire  _GEN95 = io_x[13] ? _GEN94 : _GEN93;
wire  _GEN96 = io_x[9] ? _GEN69 : _GEN70;
wire  _GEN97 = io_x[9] ? _GEN70 : _GEN69;
wire  _GEN98 = io_x[13] ? _GEN97 : _GEN96;
wire  _GEN99 = io_x[1] ? _GEN98 : _GEN95;
wire  _GEN100 = io_x[5] ? _GEN99 : _GEN92;
wire  _GEN101 = io_x[26] ? _GEN100 : _GEN85;
assign io_y[6] = _GEN101;
wire  _GEN102 = 1'b0;
wire  _GEN103 = 1'b1;
wire  _GEN104 = io_x[8] ? _GEN103 : _GEN102;
wire  _GEN105 = io_x[8] ? _GEN102 : _GEN103;
wire  _GEN106 = io_x[4] ? _GEN105 : _GEN104;
wire  _GEN107 = io_x[8] ? _GEN102 : _GEN103;
wire  _GEN108 = io_x[8] ? _GEN103 : _GEN102;
wire  _GEN109 = io_x[4] ? _GEN108 : _GEN107;
wire  _GEN110 = io_x[0] ? _GEN109 : _GEN106;
wire  _GEN111 = io_x[8] ? _GEN102 : _GEN103;
wire  _GEN112 = io_x[8] ? _GEN103 : _GEN102;
wire  _GEN113 = io_x[4] ? _GEN112 : _GEN111;
wire  _GEN114 = io_x[8] ? _GEN103 : _GEN102;
wire  _GEN115 = io_x[8] ? _GEN102 : _GEN103;
wire  _GEN116 = io_x[4] ? _GEN115 : _GEN114;
wire  _GEN117 = io_x[0] ? _GEN116 : _GEN113;
wire  _GEN118 = io_x[12] ? _GEN117 : _GEN110;
wire  _GEN119 = io_x[8] ? _GEN102 : _GEN103;
wire  _GEN120 = io_x[8] ? _GEN103 : _GEN102;
wire  _GEN121 = io_x[4] ? _GEN120 : _GEN119;
wire  _GEN122 = io_x[8] ? _GEN103 : _GEN102;
wire  _GEN123 = io_x[8] ? _GEN102 : _GEN103;
wire  _GEN124 = io_x[4] ? _GEN123 : _GEN122;
wire  _GEN125 = io_x[0] ? _GEN124 : _GEN121;
wire  _GEN126 = io_x[8] ? _GEN103 : _GEN102;
wire  _GEN127 = io_x[8] ? _GEN102 : _GEN103;
wire  _GEN128 = io_x[4] ? _GEN127 : _GEN126;
wire  _GEN129 = io_x[8] ? _GEN102 : _GEN103;
wire  _GEN130 = io_x[8] ? _GEN103 : _GEN102;
wire  _GEN131 = io_x[4] ? _GEN130 : _GEN129;
wire  _GEN132 = io_x[0] ? _GEN131 : _GEN128;
wire  _GEN133 = io_x[12] ? _GEN132 : _GEN125;
wire  _GEN134 = io_x[25] ? _GEN133 : _GEN118;
assign io_y[5] = _GEN134;
wire  _GEN135 = 1'b0;
wire  _GEN136 = 1'b1;
wire  _GEN137 = io_x[24] ? _GEN136 : _GEN135;
assign io_y[4] = _GEN137;
wire  _GEN138 = 1'b0;
wire  _GEN139 = 1'b1;
wire  _GEN140 = io_x[23] ? _GEN139 : _GEN138;
assign io_y[3] = _GEN140;
wire  _GEN141 = 1'b0;
wire  _GEN142 = 1'b1;
wire  _GEN143 = io_x[22] ? _GEN142 : _GEN141;
assign io_y[2] = _GEN143;
wire  _GEN144 = 1'b0;
wire  _GEN145 = 1'b1;
wire  _GEN146 = io_x[21] ? _GEN145 : _GEN144;
assign io_y[1] = _GEN146;
wire  _GEN147 = 1'b0;
wire  _GEN148 = 1'b1;
wire  _GEN149 = io_x[20] ? _GEN148 : _GEN147;
assign io_y[0] = _GEN149;
endmodule
module BBGSharePredictorImp_BSD_NutShell_train(
    input [31:0] train_pc,
    input  train_taken,
    input [15:0] train_ghr_rdata,
    output  pht_wdata,
    output [8:0] pht_waddr,
    output  ghr_wdata
);
wire [48:0] io_x;
wire [10:0] io_y;
assign io_x = { train_pc, train_taken, train_ghr_rdata };
assign { pht_wdata, pht_waddr, ghr_wdata } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[16] ? _GEN1 : _GEN0;
assign io_y[10] = _GEN2;
wire  _GEN3 = 1'b0;
wire  _GEN4 = 1'b1;
wire  _GEN5 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN6 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN7 = io_x[15] ? _GEN6 : _GEN5;
wire  _GEN8 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN9 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN10 = io_x[15] ? _GEN9 : _GEN8;
wire  _GEN11 = io_x[3] ? _GEN10 : _GEN7;
wire  _GEN12 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN13 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN14 = io_x[15] ? _GEN13 : _GEN12;
wire  _GEN15 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN16 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN17 = io_x[15] ? _GEN16 : _GEN15;
wire  _GEN18 = io_x[3] ? _GEN17 : _GEN14;
wire  _GEN19 = io_x[7] ? _GEN18 : _GEN11;
wire  _GEN20 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN21 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN22 = io_x[15] ? _GEN21 : _GEN20;
wire  _GEN23 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN24 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN25 = io_x[15] ? _GEN24 : _GEN23;
wire  _GEN26 = io_x[3] ? _GEN25 : _GEN22;
wire  _GEN27 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN28 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN29 = io_x[15] ? _GEN28 : _GEN27;
wire  _GEN30 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN31 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN32 = io_x[15] ? _GEN31 : _GEN30;
wire  _GEN33 = io_x[3] ? _GEN32 : _GEN29;
wire  _GEN34 = io_x[7] ? _GEN33 : _GEN26;
wire  _GEN35 = io_x[0] ? _GEN34 : _GEN19;
wire  _GEN36 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN37 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN38 = io_x[15] ? _GEN37 : _GEN36;
wire  _GEN39 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN40 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN41 = io_x[15] ? _GEN40 : _GEN39;
wire  _GEN42 = io_x[3] ? _GEN41 : _GEN38;
wire  _GEN43 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN44 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN45 = io_x[15] ? _GEN44 : _GEN43;
wire  _GEN46 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN47 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN48 = io_x[15] ? _GEN47 : _GEN46;
wire  _GEN49 = io_x[3] ? _GEN48 : _GEN45;
wire  _GEN50 = io_x[7] ? _GEN49 : _GEN42;
wire  _GEN51 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN52 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN53 = io_x[15] ? _GEN52 : _GEN51;
wire  _GEN54 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN55 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN56 = io_x[15] ? _GEN55 : _GEN54;
wire  _GEN57 = io_x[3] ? _GEN56 : _GEN53;
wire  _GEN58 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN59 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN60 = io_x[15] ? _GEN59 : _GEN58;
wire  _GEN61 = io_x[11] ? _GEN3 : _GEN4;
wire  _GEN62 = io_x[11] ? _GEN4 : _GEN3;
wire  _GEN63 = io_x[15] ? _GEN62 : _GEN61;
wire  _GEN64 = io_x[3] ? _GEN63 : _GEN60;
wire  _GEN65 = io_x[7] ? _GEN64 : _GEN57;
wire  _GEN66 = io_x[0] ? _GEN65 : _GEN50;
wire  _GEN67 = io_x[27] ? _GEN66 : _GEN35;
assign io_y[9] = _GEN67;
wire  _GEN68 = 1'b0;
wire  _GEN69 = 1'b1;
wire  _GEN70 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN71 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN72 = io_x[14] ? _GEN71 : _GEN70;
wire  _GEN73 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN74 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN75 = io_x[14] ? _GEN74 : _GEN73;
wire  _GEN76 = io_x[2] ? _GEN75 : _GEN72;
wire  _GEN77 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN78 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN79 = io_x[14] ? _GEN78 : _GEN77;
wire  _GEN80 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN81 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN82 = io_x[14] ? _GEN81 : _GEN80;
wire  _GEN83 = io_x[2] ? _GEN82 : _GEN79;
wire  _GEN84 = io_x[10] ? _GEN83 : _GEN76;
wire  _GEN85 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN86 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN87 = io_x[14] ? _GEN86 : _GEN85;
wire  _GEN88 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN89 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN90 = io_x[14] ? _GEN89 : _GEN88;
wire  _GEN91 = io_x[2] ? _GEN90 : _GEN87;
wire  _GEN92 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN93 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN94 = io_x[14] ? _GEN93 : _GEN92;
wire  _GEN95 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN96 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN97 = io_x[14] ? _GEN96 : _GEN95;
wire  _GEN98 = io_x[2] ? _GEN97 : _GEN94;
wire  _GEN99 = io_x[10] ? _GEN98 : _GEN91;
wire  _GEN100 = io_x[0] ? _GEN99 : _GEN84;
wire  _GEN101 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN102 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN103 = io_x[14] ? _GEN102 : _GEN101;
wire  _GEN104 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN105 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN106 = io_x[14] ? _GEN105 : _GEN104;
wire  _GEN107 = io_x[2] ? _GEN106 : _GEN103;
wire  _GEN108 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN109 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN110 = io_x[14] ? _GEN109 : _GEN108;
wire  _GEN111 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN112 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN113 = io_x[14] ? _GEN112 : _GEN111;
wire  _GEN114 = io_x[2] ? _GEN113 : _GEN110;
wire  _GEN115 = io_x[10] ? _GEN114 : _GEN107;
wire  _GEN116 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN117 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN118 = io_x[14] ? _GEN117 : _GEN116;
wire  _GEN119 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN120 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN121 = io_x[14] ? _GEN120 : _GEN119;
wire  _GEN122 = io_x[2] ? _GEN121 : _GEN118;
wire  _GEN123 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN124 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN125 = io_x[14] ? _GEN124 : _GEN123;
wire  _GEN126 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN127 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN128 = io_x[14] ? _GEN127 : _GEN126;
wire  _GEN129 = io_x[2] ? _GEN128 : _GEN125;
wire  _GEN130 = io_x[10] ? _GEN129 : _GEN122;
wire  _GEN131 = io_x[0] ? _GEN130 : _GEN115;
wire  _GEN132 = io_x[26] ? _GEN131 : _GEN100;
assign io_y[8] = _GEN132;
wire  _GEN133 = 1'b0;
wire  _GEN134 = 1'b1;
wire  _GEN135 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN136 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN137 = io_x[13] ? _GEN136 : _GEN135;
wire  _GEN138 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN139 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN140 = io_x[13] ? _GEN139 : _GEN138;
wire  _GEN141 = io_x[1] ? _GEN140 : _GEN137;
wire  _GEN142 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN143 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN144 = io_x[13] ? _GEN143 : _GEN142;
wire  _GEN145 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN146 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN147 = io_x[13] ? _GEN146 : _GEN145;
wire  _GEN148 = io_x[1] ? _GEN147 : _GEN144;
wire  _GEN149 = io_x[5] ? _GEN148 : _GEN141;
wire  _GEN150 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN151 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN152 = io_x[13] ? _GEN151 : _GEN150;
wire  _GEN153 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN154 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN155 = io_x[13] ? _GEN154 : _GEN153;
wire  _GEN156 = io_x[1] ? _GEN155 : _GEN152;
wire  _GEN157 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN158 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN159 = io_x[13] ? _GEN158 : _GEN157;
wire  _GEN160 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN161 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN162 = io_x[13] ? _GEN161 : _GEN160;
wire  _GEN163 = io_x[1] ? _GEN162 : _GEN159;
wire  _GEN164 = io_x[5] ? _GEN163 : _GEN156;
wire  _GEN165 = io_x[0] ? _GEN164 : _GEN149;
wire  _GEN166 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN167 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN168 = io_x[13] ? _GEN167 : _GEN166;
wire  _GEN169 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN170 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN171 = io_x[13] ? _GEN170 : _GEN169;
wire  _GEN172 = io_x[1] ? _GEN171 : _GEN168;
wire  _GEN173 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN174 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN175 = io_x[13] ? _GEN174 : _GEN173;
wire  _GEN176 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN177 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN178 = io_x[13] ? _GEN177 : _GEN176;
wire  _GEN179 = io_x[1] ? _GEN178 : _GEN175;
wire  _GEN180 = io_x[5] ? _GEN179 : _GEN172;
wire  _GEN181 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN182 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN183 = io_x[13] ? _GEN182 : _GEN181;
wire  _GEN184 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN185 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN186 = io_x[13] ? _GEN185 : _GEN184;
wire  _GEN187 = io_x[1] ? _GEN186 : _GEN183;
wire  _GEN188 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN189 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN190 = io_x[13] ? _GEN189 : _GEN188;
wire  _GEN191 = io_x[9] ? _GEN133 : _GEN134;
wire  _GEN192 = io_x[9] ? _GEN134 : _GEN133;
wire  _GEN193 = io_x[13] ? _GEN192 : _GEN191;
wire  _GEN194 = io_x[1] ? _GEN193 : _GEN190;
wire  _GEN195 = io_x[5] ? _GEN194 : _GEN187;
wire  _GEN196 = io_x[0] ? _GEN195 : _GEN180;
wire  _GEN197 = io_x[25] ? _GEN196 : _GEN165;
assign io_y[7] = _GEN197;
wire  _GEN198 = 1'b0;
wire  _GEN199 = 1'b1;
wire  _GEN200 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN201 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN202 = io_x[12] ? _GEN201 : _GEN200;
wire  _GEN203 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN204 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN205 = io_x[12] ? _GEN204 : _GEN203;
wire  _GEN206 = io_x[4] ? _GEN205 : _GEN202;
wire  _GEN207 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN208 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN209 = io_x[12] ? _GEN208 : _GEN207;
wire  _GEN210 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN211 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN212 = io_x[12] ? _GEN211 : _GEN210;
wire  _GEN213 = io_x[4] ? _GEN212 : _GEN209;
wire  _GEN214 = io_x[0] ? _GEN213 : _GEN206;
wire  _GEN215 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN216 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN217 = io_x[12] ? _GEN216 : _GEN215;
wire  _GEN218 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN219 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN220 = io_x[12] ? _GEN219 : _GEN218;
wire  _GEN221 = io_x[4] ? _GEN220 : _GEN217;
wire  _GEN222 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN223 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN224 = io_x[12] ? _GEN223 : _GEN222;
wire  _GEN225 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN226 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN227 = io_x[12] ? _GEN226 : _GEN225;
wire  _GEN228 = io_x[4] ? _GEN227 : _GEN224;
wire  _GEN229 = io_x[0] ? _GEN228 : _GEN221;
wire  _GEN230 = io_x[24] ? _GEN229 : _GEN214;
assign io_y[6] = _GEN230;
wire  _GEN231 = 1'b0;
wire  _GEN232 = 1'b1;
wire  _GEN233 = io_x[23] ? _GEN232 : _GEN231;
assign io_y[5] = _GEN233;
wire  _GEN234 = 1'b0;
wire  _GEN235 = 1'b1;
wire  _GEN236 = io_x[22] ? _GEN235 : _GEN234;
assign io_y[4] = _GEN236;
wire  _GEN237 = 1'b0;
wire  _GEN238 = 1'b1;
wire  _GEN239 = io_x[21] ? _GEN238 : _GEN237;
assign io_y[3] = _GEN239;
wire  _GEN240 = 1'b0;
wire  _GEN241 = 1'b1;
wire  _GEN242 = io_x[20] ? _GEN241 : _GEN240;
assign io_y[2] = _GEN242;
wire  _GEN243 = 1'b0;
wire  _GEN244 = 1'b1;
wire  _GEN245 = io_x[19] ? _GEN244 : _GEN243;
assign io_y[1] = _GEN245;
wire  _GEN246 = 1'b0;
wire  _GEN247 = 1'b1;
wire  _GEN248 = io_x[16] ? _GEN247 : _GEN246;
assign io_y[0] = _GEN248;
endmodule
