module BBGSharePredictorImp_BSD_sim_split(
    input [31:0] pc,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    output  taken,
    output [8:0] pht_raddr,
    input [31:0] train_pc,
    input  train_taken,
    input [15:0] train_ghr_rdata,
    output  pht_wdata,
    output [8:0] pht_waddr,
    output  ghr_wdata
);

sim_GShare_pred _pred(
    .pc        (pc),
    .pht_rdata (pht_rdata),
    .ghr_rdata (ghr_rdata),
    .taken     (taken),
    .pht_raddr (pht_raddr)
);

sim_GShare_train _train(
    .train_pc        (train_pc),
    .train_taken     (train_taken),
    .train_ghr_rdata (train_ghr_rdata),
    .pht_wdata       (pht_wdata),
    .pht_waddr       (pht_waddr),
    .ghr_wdata       (ghr_wdata)
);

endmodule

module sim_GShare_pred(
    input [31:0] pc,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    output  taken,
    output [8:0] pht_raddr
);
wire [49:0] io_x;
wire [9:0] io_y;
assign io_x = { pc, pht_rdata, ghr_rdata };
assign { taken, pht_raddr } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN3 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN4 = io_x[6] ? _GEN3 : _GEN2;
wire  _GEN5 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN6 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN7 = io_x[6] ? _GEN6 : _GEN5;
wire  _GEN8 = io_x[12] ? _GEN7 : _GEN4;
wire  _GEN9 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN10 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN11 = io_x[6] ? _GEN10 : _GEN9;
wire  _GEN12 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN13 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN14 = io_x[6] ? _GEN13 : _GEN12;
wire  _GEN15 = io_x[12] ? _GEN14 : _GEN11;
wire  _GEN16 = io_x[32] ? _GEN15 : _GEN8;
wire  _GEN17 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN18 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN19 = io_x[6] ? _GEN18 : _GEN17;
wire  _GEN20 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN21 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN22 = io_x[6] ? _GEN21 : _GEN20;
wire  _GEN23 = io_x[12] ? _GEN22 : _GEN19;
wire  _GEN24 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN25 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN26 = io_x[6] ? _GEN25 : _GEN24;
wire  _GEN27 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN28 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN29 = io_x[6] ? _GEN28 : _GEN27;
wire  _GEN30 = io_x[12] ? _GEN29 : _GEN26;
wire  _GEN31 = io_x[32] ? _GEN30 : _GEN23;
wire  _GEN32 = io_x[2] ? _GEN31 : _GEN16;
wire  _GEN33 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN34 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN35 = io_x[6] ? _GEN34 : _GEN33;
wire  _GEN36 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN37 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN38 = io_x[6] ? _GEN37 : _GEN36;
wire  _GEN39 = io_x[12] ? _GEN38 : _GEN35;
wire  _GEN40 = 1'b1;
wire  _GEN41 = io_x[32] ? _GEN40 : _GEN39;
wire  _GEN42 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN43 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN44 = io_x[6] ? _GEN43 : _GEN42;
wire  _GEN45 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN46 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN47 = io_x[6] ? _GEN46 : _GEN45;
wire  _GEN48 = io_x[12] ? _GEN47 : _GEN44;
wire  _GEN49 = io_x[32] ? _GEN40 : _GEN48;
wire  _GEN50 = io_x[2] ? _GEN49 : _GEN41;
wire  _GEN51 = io_x[31] ? _GEN50 : _GEN32;
wire  _GEN52 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN53 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN54 = io_x[6] ? _GEN53 : _GEN52;
wire  _GEN55 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN56 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN57 = io_x[6] ? _GEN56 : _GEN55;
wire  _GEN58 = io_x[12] ? _GEN57 : _GEN54;
wire  _GEN59 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN60 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN61 = io_x[6] ? _GEN60 : _GEN59;
wire  _GEN62 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN63 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN64 = io_x[6] ? _GEN63 : _GEN62;
wire  _GEN65 = io_x[12] ? _GEN64 : _GEN61;
wire  _GEN66 = io_x[32] ? _GEN65 : _GEN58;
wire  _GEN67 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN68 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN69 = io_x[6] ? _GEN68 : _GEN67;
wire  _GEN70 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN71 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN72 = io_x[6] ? _GEN71 : _GEN70;
wire  _GEN73 = io_x[12] ? _GEN72 : _GEN69;
wire  _GEN74 = 1'b0;
wire  _GEN75 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN76 = io_x[6] ? _GEN75 : _GEN74;
wire  _GEN77 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN78 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN79 = io_x[6] ? _GEN78 : _GEN77;
wire  _GEN80 = io_x[12] ? _GEN79 : _GEN76;
wire  _GEN81 = io_x[32] ? _GEN80 : _GEN73;
wire  _GEN82 = io_x[2] ? _GEN81 : _GEN66;
wire  _GEN83 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN84 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN85 = io_x[6] ? _GEN84 : _GEN83;
wire  _GEN86 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN87 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN88 = io_x[6] ? _GEN87 : _GEN86;
wire  _GEN89 = io_x[12] ? _GEN88 : _GEN85;
wire  _GEN90 = io_x[32] ? _GEN40 : _GEN89;
wire  _GEN91 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN92 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN93 = io_x[6] ? _GEN92 : _GEN91;
wire  _GEN94 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN95 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN96 = io_x[6] ? _GEN95 : _GEN94;
wire  _GEN97 = io_x[12] ? _GEN96 : _GEN93;
wire  _GEN98 = io_x[32] ? _GEN40 : _GEN97;
wire  _GEN99 = io_x[2] ? _GEN98 : _GEN90;
wire  _GEN100 = io_x[31] ? _GEN99 : _GEN82;
wire  _GEN101 = io_x[4] ? _GEN100 : _GEN51;
wire  _GEN102 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN103 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN104 = io_x[6] ? _GEN103 : _GEN102;
wire  _GEN105 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN106 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN107 = io_x[6] ? _GEN106 : _GEN105;
wire  _GEN108 = io_x[12] ? _GEN107 : _GEN104;
wire  _GEN109 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN110 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN111 = io_x[6] ? _GEN110 : _GEN109;
wire  _GEN112 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN113 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN114 = io_x[6] ? _GEN113 : _GEN112;
wire  _GEN115 = io_x[12] ? _GEN114 : _GEN111;
wire  _GEN116 = io_x[32] ? _GEN115 : _GEN108;
wire  _GEN117 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN118 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN119 = io_x[6] ? _GEN118 : _GEN117;
wire  _GEN120 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN121 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN122 = io_x[6] ? _GEN121 : _GEN120;
wire  _GEN123 = io_x[12] ? _GEN122 : _GEN119;
wire  _GEN124 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN125 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN126 = io_x[6] ? _GEN125 : _GEN124;
wire  _GEN127 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN128 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN129 = io_x[6] ? _GEN128 : _GEN127;
wire  _GEN130 = io_x[12] ? _GEN129 : _GEN126;
wire  _GEN131 = io_x[32] ? _GEN130 : _GEN123;
wire  _GEN132 = io_x[2] ? _GEN131 : _GEN116;
wire  _GEN133 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN134 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN135 = io_x[6] ? _GEN134 : _GEN133;
wire  _GEN136 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN137 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN138 = io_x[6] ? _GEN137 : _GEN136;
wire  _GEN139 = io_x[12] ? _GEN138 : _GEN135;
wire  _GEN140 = io_x[32] ? _GEN40 : _GEN139;
wire  _GEN141 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN142 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN143 = io_x[6] ? _GEN142 : _GEN141;
wire  _GEN144 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN145 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN146 = io_x[6] ? _GEN145 : _GEN144;
wire  _GEN147 = io_x[12] ? _GEN146 : _GEN143;
wire  _GEN148 = io_x[32] ? _GEN40 : _GEN147;
wire  _GEN149 = io_x[2] ? _GEN148 : _GEN140;
wire  _GEN150 = io_x[31] ? _GEN149 : _GEN132;
wire  _GEN151 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN152 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN153 = io_x[6] ? _GEN152 : _GEN151;
wire  _GEN154 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN155 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN156 = io_x[6] ? _GEN155 : _GEN154;
wire  _GEN157 = io_x[12] ? _GEN156 : _GEN153;
wire  _GEN158 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN159 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN160 = io_x[6] ? _GEN159 : _GEN158;
wire  _GEN161 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN162 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN163 = io_x[6] ? _GEN162 : _GEN161;
wire  _GEN164 = io_x[12] ? _GEN163 : _GEN160;
wire  _GEN165 = io_x[32] ? _GEN164 : _GEN157;
wire  _GEN166 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN167 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN168 = io_x[6] ? _GEN167 : _GEN166;
wire  _GEN169 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN170 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN171 = io_x[6] ? _GEN170 : _GEN169;
wire  _GEN172 = io_x[12] ? _GEN171 : _GEN168;
wire  _GEN173 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN174 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN175 = io_x[6] ? _GEN174 : _GEN173;
wire  _GEN176 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN177 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN178 = io_x[6] ? _GEN177 : _GEN176;
wire  _GEN179 = io_x[12] ? _GEN178 : _GEN175;
wire  _GEN180 = io_x[32] ? _GEN179 : _GEN172;
wire  _GEN181 = io_x[2] ? _GEN180 : _GEN165;
wire  _GEN182 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN183 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN184 = io_x[6] ? _GEN183 : _GEN182;
wire  _GEN185 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN186 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN187 = io_x[6] ? _GEN186 : _GEN185;
wire  _GEN188 = io_x[12] ? _GEN187 : _GEN184;
wire  _GEN189 = io_x[32] ? _GEN40 : _GEN188;
wire  _GEN190 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN191 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN192 = io_x[6] ? _GEN191 : _GEN190;
wire  _GEN193 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN194 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN195 = io_x[6] ? _GEN194 : _GEN193;
wire  _GEN196 = io_x[12] ? _GEN195 : _GEN192;
wire  _GEN197 = io_x[32] ? _GEN40 : _GEN196;
wire  _GEN198 = io_x[2] ? _GEN197 : _GEN189;
wire  _GEN199 = io_x[31] ? _GEN198 : _GEN181;
wire  _GEN200 = io_x[4] ? _GEN199 : _GEN150;
wire  _GEN201 = io_x[0] ? _GEN200 : _GEN101;
assign io_y[9] = _GEN201;
wire  _GEN202 = 1'b0;
wire  _GEN203 = 1'b1;
wire  _GEN204 = 1'b1;
wire  _GEN205 = 1'b0;
wire  _GEN206 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN207 = 1'b0;
wire  _GEN208 = io_x[11] ? _GEN207 : _GEN206;
wire  _GEN209 = 1'b0;
wire  _GEN210 = io_x[3] ? _GEN209 : _GEN208;
wire  _GEN211 = io_x[7] ? _GEN210 : _GEN203;
wire  _GEN212 = io_x[2] ? _GEN211 : _GEN202;
wire  _GEN213 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN214 = 1'b1;
wire  _GEN215 = io_x[11] ? _GEN214 : _GEN213;
wire  _GEN216 = 1'b1;
wire  _GEN217 = io_x[3] ? _GEN216 : _GEN215;
wire  _GEN218 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN219 = io_x[11] ? _GEN218 : _GEN207;
wire  _GEN220 = io_x[3] ? _GEN219 : _GEN216;
wire  _GEN221 = io_x[7] ? _GEN220 : _GEN217;
wire  _GEN222 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN223 = io_x[11] ? _GEN222 : _GEN214;
wire  _GEN224 = io_x[3] ? _GEN223 : _GEN216;
wire  _GEN225 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN226 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN227 = io_x[11] ? _GEN226 : _GEN225;
wire  _GEN228 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN229 = io_x[3] ? _GEN228 : _GEN227;
wire  _GEN230 = io_x[7] ? _GEN229 : _GEN224;
wire  _GEN231 = io_x[2] ? _GEN230 : _GEN221;
wire  _GEN232 = io_x[17] ? _GEN231 : _GEN212;
wire  _GEN233 = 1'b1;
wire  _GEN234 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN235 = io_x[11] ? _GEN234 : _GEN214;
wire  _GEN236 = io_x[3] ? _GEN216 : _GEN235;
wire  _GEN237 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN238 = io_x[3] ? _GEN216 : _GEN237;
wire  _GEN239 = io_x[7] ? _GEN238 : _GEN236;
wire  _GEN240 = io_x[2] ? _GEN239 : _GEN233;
wire  _GEN241 = 1'b0;
wire  _GEN242 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN243 = io_x[11] ? _GEN242 : _GEN214;
wire  _GEN244 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN245 = io_x[11] ? _GEN244 : _GEN214;
wire  _GEN246 = io_x[3] ? _GEN245 : _GEN243;
wire  _GEN247 = io_x[7] ? _GEN246 : _GEN241;
wire  _GEN248 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN249 = io_x[11] ? _GEN248 : _GEN207;
wire  _GEN250 = io_x[3] ? _GEN216 : _GEN249;
wire  _GEN251 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN252 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN253 = io_x[11] ? _GEN252 : _GEN251;
wire  _GEN254 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN255 = io_x[11] ? _GEN254 : _GEN207;
wire  _GEN256 = io_x[3] ? _GEN255 : _GEN253;
wire  _GEN257 = io_x[7] ? _GEN256 : _GEN250;
wire  _GEN258 = io_x[2] ? _GEN257 : _GEN247;
wire  _GEN259 = io_x[17] ? _GEN258 : _GEN240;
wire  _GEN260 = io_x[15] ? _GEN259 : _GEN232;
wire  _GEN261 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN262 = io_x[11] ? _GEN261 : _GEN214;
wire  _GEN263 = io_x[3] ? _GEN209 : _GEN262;
wire  _GEN264 = io_x[7] ? _GEN263 : _GEN241;
wire  _GEN265 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN266 = io_x[3] ? _GEN209 : _GEN265;
wire  _GEN267 = io_x[7] ? _GEN266 : _GEN203;
wire  _GEN268 = io_x[2] ? _GEN267 : _GEN264;
wire  _GEN269 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN270 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN271 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN272 = io_x[11] ? _GEN271 : _GEN214;
wire  _GEN273 = io_x[3] ? _GEN272 : _GEN270;
wire  _GEN274 = io_x[7] ? _GEN273 : _GEN241;
wire  _GEN275 = io_x[2] ? _GEN274 : _GEN269;
wire  _GEN276 = io_x[17] ? _GEN275 : _GEN268;
wire  _GEN277 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN278 = io_x[11] ? _GEN214 : _GEN277;
wire  _GEN279 = io_x[3] ? _GEN278 : _GEN216;
wire  _GEN280 = io_x[7] ? _GEN279 : _GEN203;
wire  _GEN281 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN282 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN283 = io_x[3] ? _GEN282 : _GEN216;
wire  _GEN284 = io_x[7] ? _GEN283 : _GEN281;
wire  _GEN285 = io_x[2] ? _GEN284 : _GEN280;
wire  _GEN286 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN287 = io_x[3] ? _GEN286 : _GEN216;
wire  _GEN288 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN289 = io_x[11] ? _GEN214 : _GEN288;
wire  _GEN290 = io_x[3] ? _GEN289 : _GEN216;
wire  _GEN291 = io_x[7] ? _GEN290 : _GEN287;
wire  _GEN292 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN293 = io_x[3] ? _GEN216 : _GEN292;
wire  _GEN294 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN295 = io_x[11] ? _GEN294 : _GEN214;
wire  _GEN296 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN297 = io_x[11] ? _GEN296 : _GEN207;
wire  _GEN298 = io_x[3] ? _GEN297 : _GEN295;
wire  _GEN299 = io_x[7] ? _GEN298 : _GEN293;
wire  _GEN300 = io_x[2] ? _GEN299 : _GEN291;
wire  _GEN301 = io_x[17] ? _GEN300 : _GEN285;
wire  _GEN302 = io_x[15] ? _GEN301 : _GEN276;
wire  _GEN303 = io_x[12] ? _GEN302 : _GEN260;
wire  _GEN304 = io_x[7] ? _GEN203 : _GEN241;
wire  _GEN305 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN306 = io_x[3] ? _GEN305 : _GEN209;
wire  _GEN307 = io_x[7] ? _GEN306 : _GEN203;
wire  _GEN308 = io_x[2] ? _GEN307 : _GEN304;
wire  _GEN309 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN310 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN311 = io_x[3] ? _GEN310 : _GEN216;
wire  _GEN312 = io_x[7] ? _GEN311 : _GEN309;
wire  _GEN313 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN314 = io_x[11] ? _GEN313 : _GEN214;
wire  _GEN315 = io_x[3] ? _GEN314 : _GEN216;
wire  _GEN316 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN317 = io_x[11] ? _GEN316 : _GEN214;
wire  _GEN318 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN319 = io_x[3] ? _GEN318 : _GEN317;
wire  _GEN320 = io_x[7] ? _GEN319 : _GEN315;
wire  _GEN321 = io_x[2] ? _GEN320 : _GEN312;
wire  _GEN322 = io_x[17] ? _GEN321 : _GEN308;
wire  _GEN323 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN324 = io_x[3] ? _GEN216 : _GEN323;
wire  _GEN325 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN326 = io_x[11] ? _GEN325 : _GEN207;
wire  _GEN327 = io_x[3] ? _GEN326 : _GEN209;
wire  _GEN328 = io_x[7] ? _GEN327 : _GEN324;
wire  _GEN329 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN330 = io_x[11] ? _GEN214 : _GEN329;
wire  _GEN331 = io_x[3] ? _GEN330 : _GEN216;
wire  _GEN332 = io_x[7] ? _GEN331 : _GEN241;
wire  _GEN333 = io_x[2] ? _GEN332 : _GEN328;
wire  _GEN334 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN335 = io_x[11] ? _GEN214 : _GEN334;
wire  _GEN336 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN337 = io_x[11] ? _GEN336 : _GEN214;
wire  _GEN338 = io_x[3] ? _GEN337 : _GEN335;
wire  _GEN339 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN340 = io_x[3] ? _GEN339 : _GEN216;
wire  _GEN341 = io_x[7] ? _GEN340 : _GEN338;
wire  _GEN342 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN343 = io_x[11] ? _GEN342 : _GEN214;
wire  _GEN344 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN345 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN346 = io_x[11] ? _GEN345 : _GEN344;
wire  _GEN347 = io_x[3] ? _GEN346 : _GEN343;
wire  _GEN348 = io_x[7] ? _GEN347 : _GEN203;
wire  _GEN349 = io_x[2] ? _GEN348 : _GEN341;
wire  _GEN350 = io_x[17] ? _GEN349 : _GEN333;
wire  _GEN351 = io_x[15] ? _GEN350 : _GEN322;
wire  _GEN352 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN353 = io_x[11] ? _GEN214 : _GEN352;
wire  _GEN354 = io_x[3] ? _GEN353 : _GEN216;
wire  _GEN355 = io_x[7] ? _GEN354 : _GEN203;
wire  _GEN356 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN357 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN358 = io_x[11] ? _GEN357 : _GEN207;
wire  _GEN359 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN360 = io_x[11] ? _GEN359 : _GEN214;
wire  _GEN361 = io_x[3] ? _GEN360 : _GEN358;
wire  _GEN362 = io_x[7] ? _GEN361 : _GEN356;
wire  _GEN363 = io_x[2] ? _GEN362 : _GEN355;
wire  _GEN364 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN365 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN366 = io_x[11] ? _GEN207 : _GEN365;
wire  _GEN367 = io_x[3] ? _GEN366 : _GEN216;
wire  _GEN368 = io_x[7] ? _GEN367 : _GEN364;
wire  _GEN369 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN370 = io_x[11] ? _GEN207 : _GEN369;
wire  _GEN371 = io_x[3] ? _GEN370 : _GEN209;
wire  _GEN372 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN373 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN374 = io_x[3] ? _GEN373 : _GEN372;
wire  _GEN375 = io_x[7] ? _GEN374 : _GEN371;
wire  _GEN376 = io_x[2] ? _GEN375 : _GEN368;
wire  _GEN377 = io_x[17] ? _GEN376 : _GEN363;
wire  _GEN378 = io_x[7] ? _GEN203 : _GEN241;
wire  _GEN379 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN380 = io_x[11] ? _GEN379 : _GEN207;
wire  _GEN381 = io_x[3] ? _GEN380 : _GEN216;
wire  _GEN382 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN383 = io_x[11] ? _GEN382 : _GEN214;
wire  _GEN384 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN385 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN386 = io_x[11] ? _GEN385 : _GEN384;
wire  _GEN387 = io_x[3] ? _GEN386 : _GEN383;
wire  _GEN388 = io_x[7] ? _GEN387 : _GEN381;
wire  _GEN389 = io_x[2] ? _GEN388 : _GEN378;
wire  _GEN390 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN391 = io_x[3] ? _GEN390 : _GEN216;
wire  _GEN392 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN393 = io_x[11] ? _GEN392 : _GEN214;
wire  _GEN394 = io_x[3] ? _GEN393 : _GEN216;
wire  _GEN395 = io_x[7] ? _GEN394 : _GEN391;
wire  _GEN396 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN397 = io_x[11] ? _GEN396 : _GEN214;
wire  _GEN398 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN399 = io_x[11] ? _GEN207 : _GEN398;
wire  _GEN400 = io_x[3] ? _GEN399 : _GEN397;
wire  _GEN401 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN402 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN403 = io_x[11] ? _GEN402 : _GEN401;
wire  _GEN404 = io_x[3] ? _GEN403 : _GEN209;
wire  _GEN405 = io_x[7] ? _GEN404 : _GEN400;
wire  _GEN406 = io_x[2] ? _GEN405 : _GEN395;
wire  _GEN407 = io_x[17] ? _GEN406 : _GEN389;
wire  _GEN408 = io_x[15] ? _GEN407 : _GEN377;
wire  _GEN409 = io_x[12] ? _GEN408 : _GEN351;
wire  _GEN410 = io_x[10] ? _GEN409 : _GEN303;
wire  _GEN411 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN412 = io_x[11] ? _GEN411 : _GEN214;
wire  _GEN413 = io_x[3] ? _GEN216 : _GEN412;
wire  _GEN414 = io_x[7] ? _GEN413 : _GEN203;
wire  _GEN415 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN416 = io_x[11] ? _GEN415 : _GEN214;
wire  _GEN417 = io_x[3] ? _GEN209 : _GEN416;
wire  _GEN418 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN419 = io_x[11] ? _GEN418 : _GEN214;
wire  _GEN420 = io_x[3] ? _GEN209 : _GEN419;
wire  _GEN421 = io_x[7] ? _GEN420 : _GEN417;
wire  _GEN422 = io_x[2] ? _GEN421 : _GEN414;
wire  _GEN423 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN424 = io_x[11] ? _GEN423 : _GEN214;
wire  _GEN425 = io_x[3] ? _GEN216 : _GEN424;
wire  _GEN426 = io_x[7] ? _GEN425 : _GEN203;
wire  _GEN427 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN428 = io_x[3] ? _GEN209 : _GEN427;
wire  _GEN429 = io_x[7] ? _GEN428 : _GEN241;
wire  _GEN430 = io_x[2] ? _GEN429 : _GEN426;
wire  _GEN431 = io_x[17] ? _GEN430 : _GEN422;
wire  _GEN432 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN433 = io_x[3] ? _GEN216 : _GEN432;
wire  _GEN434 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN435 = io_x[11] ? _GEN434 : _GEN214;
wire  _GEN436 = io_x[3] ? _GEN216 : _GEN435;
wire  _GEN437 = io_x[7] ? _GEN436 : _GEN433;
wire  _GEN438 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN439 = io_x[11] ? _GEN438 : _GEN207;
wire  _GEN440 = io_x[3] ? _GEN216 : _GEN439;
wire  _GEN441 = io_x[7] ? _GEN440 : _GEN241;
wire  _GEN442 = io_x[2] ? _GEN441 : _GEN437;
wire  _GEN443 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN444 = io_x[11] ? _GEN443 : _GEN207;
wire  _GEN445 = io_x[3] ? _GEN216 : _GEN444;
wire  _GEN446 = io_x[7] ? _GEN445 : _GEN203;
wire  _GEN447 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN448 = io_x[11] ? _GEN447 : _GEN207;
wire  _GEN449 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN450 = io_x[11] ? _GEN207 : _GEN449;
wire  _GEN451 = io_x[3] ? _GEN450 : _GEN448;
wire  _GEN452 = io_x[7] ? _GEN203 : _GEN451;
wire  _GEN453 = io_x[2] ? _GEN452 : _GEN446;
wire  _GEN454 = io_x[17] ? _GEN453 : _GEN442;
wire  _GEN455 = io_x[15] ? _GEN454 : _GEN431;
wire  _GEN456 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN457 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN458 = io_x[11] ? _GEN457 : _GEN214;
wire  _GEN459 = io_x[3] ? _GEN458 : _GEN456;
wire  _GEN460 = io_x[7] ? _GEN459 : _GEN203;
wire  _GEN461 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN462 = io_x[11] ? _GEN461 : _GEN207;
wire  _GEN463 = io_x[3] ? _GEN216 : _GEN462;
wire  _GEN464 = io_x[7] ? _GEN203 : _GEN463;
wire  _GEN465 = io_x[2] ? _GEN464 : _GEN460;
wire  _GEN466 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN467 = io_x[11] ? _GEN466 : _GEN214;
wire  _GEN468 = io_x[3] ? _GEN467 : _GEN216;
wire  _GEN469 = io_x[7] ? _GEN468 : _GEN241;
wire  _GEN470 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN471 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN472 = io_x[11] ? _GEN471 : _GEN470;
wire  _GEN473 = io_x[3] ? _GEN216 : _GEN472;
wire  _GEN474 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN475 = io_x[11] ? _GEN474 : _GEN214;
wire  _GEN476 = io_x[3] ? _GEN475 : _GEN216;
wire  _GEN477 = io_x[7] ? _GEN476 : _GEN473;
wire  _GEN478 = io_x[2] ? _GEN477 : _GEN469;
wire  _GEN479 = io_x[17] ? _GEN478 : _GEN465;
wire  _GEN480 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN481 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN482 = io_x[3] ? _GEN481 : _GEN480;
wire  _GEN483 = io_x[7] ? _GEN482 : _GEN203;
wire  _GEN484 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN485 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN486 = io_x[11] ? _GEN485 : _GEN484;
wire  _GEN487 = io_x[3] ? _GEN486 : _GEN209;
wire  _GEN488 = io_x[7] ? _GEN487 : _GEN203;
wire  _GEN489 = io_x[2] ? _GEN488 : _GEN483;
wire  _GEN490 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN491 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN492 = io_x[11] ? _GEN491 : _GEN207;
wire  _GEN493 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN494 = io_x[11] ? _GEN493 : _GEN207;
wire  _GEN495 = io_x[3] ? _GEN494 : _GEN492;
wire  _GEN496 = io_x[7] ? _GEN495 : _GEN490;
wire  _GEN497 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN498 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN499 = io_x[11] ? _GEN498 : _GEN497;
wire  _GEN500 = io_x[3] ? _GEN499 : _GEN209;
wire  _GEN501 = io_x[7] ? _GEN500 : _GEN241;
wire  _GEN502 = io_x[2] ? _GEN501 : _GEN496;
wire  _GEN503 = io_x[17] ? _GEN502 : _GEN489;
wire  _GEN504 = io_x[15] ? _GEN503 : _GEN479;
wire  _GEN505 = io_x[12] ? _GEN504 : _GEN455;
wire  _GEN506 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN507 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN508 = io_x[11] ? _GEN507 : _GEN214;
wire  _GEN509 = io_x[3] ? _GEN508 : _GEN506;
wire  _GEN510 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN511 = io_x[3] ? _GEN216 : _GEN510;
wire  _GEN512 = io_x[7] ? _GEN511 : _GEN509;
wire  _GEN513 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN514 = io_x[3] ? _GEN216 : _GEN513;
wire  _GEN515 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN516 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN517 = io_x[11] ? _GEN516 : _GEN515;
wire  _GEN518 = io_x[3] ? _GEN216 : _GEN517;
wire  _GEN519 = io_x[7] ? _GEN518 : _GEN514;
wire  _GEN520 = io_x[2] ? _GEN519 : _GEN512;
wire  _GEN521 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN522 = io_x[11] ? _GEN214 : _GEN521;
wire  _GEN523 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN524 = io_x[3] ? _GEN523 : _GEN522;
wire  _GEN525 = io_x[7] ? _GEN524 : _GEN241;
wire  _GEN526 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN527 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN528 = io_x[11] ? _GEN527 : _GEN214;
wire  _GEN529 = io_x[3] ? _GEN528 : _GEN209;
wire  _GEN530 = io_x[7] ? _GEN529 : _GEN526;
wire  _GEN531 = io_x[2] ? _GEN530 : _GEN525;
wire  _GEN532 = io_x[17] ? _GEN531 : _GEN520;
wire  _GEN533 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN534 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN535 = io_x[11] ? _GEN214 : _GEN534;
wire  _GEN536 = io_x[3] ? _GEN535 : _GEN216;
wire  _GEN537 = io_x[7] ? _GEN536 : _GEN533;
wire  _GEN538 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN539 = io_x[11] ? _GEN207 : _GEN538;
wire  _GEN540 = io_x[3] ? _GEN539 : _GEN216;
wire  _GEN541 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN542 = io_x[11] ? _GEN207 : _GEN541;
wire  _GEN543 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN544 = io_x[3] ? _GEN543 : _GEN542;
wire  _GEN545 = io_x[7] ? _GEN544 : _GEN540;
wire  _GEN546 = io_x[2] ? _GEN545 : _GEN537;
wire  _GEN547 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN548 = io_x[11] ? _GEN547 : _GEN207;
wire  _GEN549 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN550 = io_x[11] ? _GEN549 : _GEN207;
wire  _GEN551 = io_x[3] ? _GEN550 : _GEN548;
wire  _GEN552 = io_x[7] ? _GEN551 : _GEN203;
wire  _GEN553 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN554 = io_x[11] ? _GEN214 : _GEN553;
wire  _GEN555 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN556 = io_x[11] ? _GEN214 : _GEN555;
wire  _GEN557 = io_x[3] ? _GEN556 : _GEN554;
wire  _GEN558 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN559 = io_x[11] ? _GEN558 : _GEN207;
wire  _GEN560 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN561 = io_x[11] ? _GEN560 : _GEN214;
wire  _GEN562 = io_x[3] ? _GEN561 : _GEN559;
wire  _GEN563 = io_x[7] ? _GEN562 : _GEN557;
wire  _GEN564 = io_x[2] ? _GEN563 : _GEN552;
wire  _GEN565 = io_x[17] ? _GEN564 : _GEN546;
wire  _GEN566 = io_x[15] ? _GEN565 : _GEN532;
wire  _GEN567 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN568 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN569 = io_x[3] ? _GEN216 : _GEN568;
wire  _GEN570 = io_x[7] ? _GEN569 : _GEN567;
wire  _GEN571 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN572 = io_x[11] ? _GEN571 : _GEN207;
wire  _GEN573 = io_x[3] ? _GEN572 : _GEN209;
wire  _GEN574 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN575 = io_x[7] ? _GEN574 : _GEN573;
wire  _GEN576 = io_x[2] ? _GEN575 : _GEN570;
wire  _GEN577 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN578 = io_x[11] ? _GEN577 : _GEN207;
wire  _GEN579 = io_x[3] ? _GEN216 : _GEN578;
wire  _GEN580 = io_x[7] ? _GEN579 : _GEN241;
wire  _GEN581 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN582 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN583 = io_x[11] ? _GEN214 : _GEN582;
wire  _GEN584 = io_x[3] ? _GEN583 : _GEN581;
wire  _GEN585 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN586 = io_x[7] ? _GEN585 : _GEN584;
wire  _GEN587 = io_x[2] ? _GEN586 : _GEN580;
wire  _GEN588 = io_x[17] ? _GEN587 : _GEN576;
wire  _GEN589 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN590 = io_x[11] ? _GEN214 : _GEN589;
wire  _GEN591 = io_x[3] ? _GEN590 : _GEN209;
wire  _GEN592 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN593 = io_x[11] ? _GEN592 : _GEN214;
wire  _GEN594 = io_x[3] ? _GEN209 : _GEN593;
wire  _GEN595 = io_x[7] ? _GEN594 : _GEN591;
wire  _GEN596 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN597 = io_x[3] ? _GEN209 : _GEN596;
wire  _GEN598 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN599 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN600 = io_x[11] ? _GEN599 : _GEN598;
wire  _GEN601 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN602 = io_x[3] ? _GEN601 : _GEN600;
wire  _GEN603 = io_x[7] ? _GEN602 : _GEN597;
wire  _GEN604 = io_x[2] ? _GEN603 : _GEN595;
wire  _GEN605 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN606 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN607 = io_x[11] ? _GEN606 : _GEN214;
wire  _GEN608 = io_x[3] ? _GEN607 : _GEN605;
wire  _GEN609 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN610 = io_x[11] ? _GEN609 : _GEN214;
wire  _GEN611 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN612 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN613 = io_x[11] ? _GEN612 : _GEN611;
wire  _GEN614 = io_x[3] ? _GEN613 : _GEN610;
wire  _GEN615 = io_x[7] ? _GEN614 : _GEN608;
wire  _GEN616 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN617 = io_x[11] ? _GEN214 : _GEN616;
wire  _GEN618 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN619 = io_x[11] ? _GEN618 : _GEN214;
wire  _GEN620 = io_x[3] ? _GEN619 : _GEN617;
wire  _GEN621 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN622 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN623 = io_x[11] ? _GEN622 : _GEN621;
wire  _GEN624 = io_x[3] ? _GEN623 : _GEN216;
wire  _GEN625 = io_x[7] ? _GEN624 : _GEN620;
wire  _GEN626 = io_x[2] ? _GEN625 : _GEN615;
wire  _GEN627 = io_x[17] ? _GEN626 : _GEN604;
wire  _GEN628 = io_x[15] ? _GEN627 : _GEN588;
wire  _GEN629 = io_x[12] ? _GEN628 : _GEN566;
wire  _GEN630 = io_x[10] ? _GEN629 : _GEN505;
wire  _GEN631 = io_x[4] ? _GEN630 : _GEN410;
wire  _GEN632 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN633 = io_x[3] ? _GEN632 : _GEN216;
wire  _GEN634 = io_x[7] ? _GEN633 : _GEN203;
wire  _GEN635 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN636 = io_x[3] ? _GEN635 : _GEN216;
wire  _GEN637 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN638 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN639 = io_x[3] ? _GEN638 : _GEN637;
wire  _GEN640 = io_x[7] ? _GEN639 : _GEN636;
wire  _GEN641 = io_x[2] ? _GEN640 : _GEN634;
wire  _GEN642 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN643 = io_x[11] ? _GEN642 : _GEN214;
wire  _GEN644 = io_x[3] ? _GEN216 : _GEN643;
wire  _GEN645 = io_x[7] ? _GEN241 : _GEN644;
wire  _GEN646 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN647 = io_x[11] ? _GEN646 : _GEN207;
wire  _GEN648 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN649 = io_x[3] ? _GEN648 : _GEN647;
wire  _GEN650 = io_x[7] ? _GEN649 : _GEN241;
wire  _GEN651 = io_x[2] ? _GEN650 : _GEN645;
wire  _GEN652 = io_x[17] ? _GEN651 : _GEN641;
wire  _GEN653 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN654 = io_x[7] ? _GEN203 : _GEN653;
wire  _GEN655 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN656 = io_x[7] ? _GEN655 : _GEN203;
wire  _GEN657 = io_x[2] ? _GEN656 : _GEN654;
wire  _GEN658 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN659 = io_x[11] ? _GEN658 : _GEN214;
wire  _GEN660 = io_x[3] ? _GEN659 : _GEN216;
wire  _GEN661 = io_x[7] ? _GEN660 : _GEN203;
wire  _GEN662 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN663 = io_x[11] ? _GEN662 : _GEN214;
wire  _GEN664 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN665 = io_x[11] ? _GEN664 : _GEN214;
wire  _GEN666 = io_x[3] ? _GEN665 : _GEN663;
wire  _GEN667 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN668 = io_x[11] ? _GEN667 : _GEN214;
wire  _GEN669 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN670 = io_x[3] ? _GEN669 : _GEN668;
wire  _GEN671 = io_x[7] ? _GEN670 : _GEN666;
wire  _GEN672 = io_x[2] ? _GEN671 : _GEN661;
wire  _GEN673 = io_x[17] ? _GEN672 : _GEN657;
wire  _GEN674 = io_x[15] ? _GEN673 : _GEN652;
wire  _GEN675 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN676 = io_x[11] ? _GEN675 : _GEN214;
wire  _GEN677 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN678 = io_x[11] ? _GEN677 : _GEN207;
wire  _GEN679 = io_x[3] ? _GEN678 : _GEN676;
wire  _GEN680 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN681 = io_x[11] ? _GEN680 : _GEN214;
wire  _GEN682 = io_x[3] ? _GEN209 : _GEN681;
wire  _GEN683 = io_x[7] ? _GEN682 : _GEN679;
wire  _GEN684 = io_x[2] ? _GEN683 : _GEN202;
wire  _GEN685 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN686 = io_x[7] ? _GEN203 : _GEN685;
wire  _GEN687 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN688 = io_x[11] ? _GEN687 : _GEN207;
wire  _GEN689 = io_x[3] ? _GEN688 : _GEN216;
wire  _GEN690 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN691 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN692 = io_x[11] ? _GEN691 : _GEN214;
wire  _GEN693 = io_x[3] ? _GEN692 : _GEN690;
wire  _GEN694 = io_x[7] ? _GEN693 : _GEN689;
wire  _GEN695 = io_x[2] ? _GEN694 : _GEN686;
wire  _GEN696 = io_x[17] ? _GEN695 : _GEN684;
wire  _GEN697 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN698 = io_x[11] ? _GEN214 : _GEN697;
wire  _GEN699 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN700 = io_x[3] ? _GEN699 : _GEN698;
wire  _GEN701 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN702 = io_x[7] ? _GEN701 : _GEN700;
wire  _GEN703 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN704 = io_x[11] ? _GEN207 : _GEN703;
wire  _GEN705 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN706 = io_x[11] ? _GEN214 : _GEN705;
wire  _GEN707 = io_x[3] ? _GEN706 : _GEN704;
wire  _GEN708 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN709 = io_x[11] ? _GEN708 : _GEN214;
wire  _GEN710 = io_x[3] ? _GEN209 : _GEN709;
wire  _GEN711 = io_x[7] ? _GEN710 : _GEN707;
wire  _GEN712 = io_x[2] ? _GEN711 : _GEN702;
wire  _GEN713 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN714 = io_x[11] ? _GEN214 : _GEN713;
wire  _GEN715 = io_x[3] ? _GEN714 : _GEN216;
wire  _GEN716 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN717 = io_x[11] ? _GEN214 : _GEN716;
wire  _GEN718 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN719 = io_x[3] ? _GEN718 : _GEN717;
wire  _GEN720 = io_x[7] ? _GEN719 : _GEN715;
wire  _GEN721 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN722 = io_x[11] ? _GEN214 : _GEN721;
wire  _GEN723 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN724 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN725 = io_x[11] ? _GEN724 : _GEN723;
wire  _GEN726 = io_x[3] ? _GEN725 : _GEN722;
wire  _GEN727 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN728 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN729 = io_x[11] ? _GEN728 : _GEN727;
wire  _GEN730 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN731 = io_x[11] ? _GEN730 : _GEN214;
wire  _GEN732 = io_x[3] ? _GEN731 : _GEN729;
wire  _GEN733 = io_x[7] ? _GEN732 : _GEN726;
wire  _GEN734 = io_x[2] ? _GEN733 : _GEN720;
wire  _GEN735 = io_x[17] ? _GEN734 : _GEN712;
wire  _GEN736 = io_x[15] ? _GEN735 : _GEN696;
wire  _GEN737 = io_x[12] ? _GEN736 : _GEN674;
wire  _GEN738 = io_x[7] ? _GEN203 : _GEN241;
wire  _GEN739 = io_x[2] ? _GEN233 : _GEN738;
wire  _GEN740 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN741 = io_x[3] ? _GEN209 : _GEN740;
wire  _GEN742 = io_x[7] ? _GEN203 : _GEN741;
wire  _GEN743 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN744 = io_x[11] ? _GEN207 : _GEN743;
wire  _GEN745 = io_x[3] ? _GEN209 : _GEN744;
wire  _GEN746 = io_x[7] ? _GEN203 : _GEN745;
wire  _GEN747 = io_x[2] ? _GEN746 : _GEN742;
wire  _GEN748 = io_x[17] ? _GEN747 : _GEN739;
wire  _GEN749 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN750 = io_x[11] ? _GEN207 : _GEN749;
wire  _GEN751 = io_x[3] ? _GEN750 : _GEN216;
wire  _GEN752 = io_x[7] ? _GEN241 : _GEN751;
wire  _GEN753 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN754 = io_x[11] ? _GEN753 : _GEN214;
wire  _GEN755 = io_x[3] ? _GEN216 : _GEN754;
wire  _GEN756 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN757 = io_x[11] ? _GEN756 : _GEN207;
wire  _GEN758 = io_x[3] ? _GEN757 : _GEN216;
wire  _GEN759 = io_x[7] ? _GEN758 : _GEN755;
wire  _GEN760 = io_x[2] ? _GEN759 : _GEN752;
wire  _GEN761 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN762 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN763 = io_x[11] ? _GEN762 : _GEN761;
wire  _GEN764 = io_x[3] ? _GEN763 : _GEN209;
wire  _GEN765 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN766 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN767 = io_x[11] ? _GEN766 : _GEN765;
wire  _GEN768 = io_x[3] ? _GEN767 : _GEN209;
wire  _GEN769 = io_x[7] ? _GEN768 : _GEN764;
wire  _GEN770 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN771 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN772 = io_x[11] ? _GEN771 : _GEN770;
wire  _GEN773 = io_x[3] ? _GEN772 : _GEN216;
wire  _GEN774 = io_x[7] ? _GEN773 : _GEN241;
wire  _GEN775 = io_x[2] ? _GEN774 : _GEN769;
wire  _GEN776 = io_x[17] ? _GEN775 : _GEN760;
wire  _GEN777 = io_x[15] ? _GEN776 : _GEN748;
wire  _GEN778 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN779 = io_x[11] ? _GEN214 : _GEN778;
wire  _GEN780 = io_x[3] ? _GEN779 : _GEN216;
wire  _GEN781 = io_x[7] ? _GEN241 : _GEN780;
wire  _GEN782 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN783 = io_x[11] ? _GEN782 : _GEN214;
wire  _GEN784 = io_x[3] ? _GEN209 : _GEN783;
wire  _GEN785 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN786 = io_x[11] ? _GEN785 : _GEN214;
wire  _GEN787 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN788 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN789 = io_x[11] ? _GEN788 : _GEN787;
wire  _GEN790 = io_x[3] ? _GEN789 : _GEN786;
wire  _GEN791 = io_x[7] ? _GEN790 : _GEN784;
wire  _GEN792 = io_x[2] ? _GEN791 : _GEN781;
wire  _GEN793 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN794 = io_x[11] ? _GEN214 : _GEN793;
wire  _GEN795 = io_x[3] ? _GEN794 : _GEN216;
wire  _GEN796 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN797 = io_x[11] ? _GEN796 : _GEN214;
wire  _GEN798 = io_x[3] ? _GEN797 : _GEN216;
wire  _GEN799 = io_x[7] ? _GEN798 : _GEN795;
wire  _GEN800 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN801 = io_x[3] ? _GEN209 : _GEN800;
wire  _GEN802 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN803 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN804 = io_x[11] ? _GEN803 : _GEN802;
wire  _GEN805 = io_x[3] ? _GEN804 : _GEN209;
wire  _GEN806 = io_x[7] ? _GEN805 : _GEN801;
wire  _GEN807 = io_x[2] ? _GEN806 : _GEN799;
wire  _GEN808 = io_x[17] ? _GEN807 : _GEN792;
wire  _GEN809 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN810 = io_x[11] ? _GEN809 : _GEN214;
wire  _GEN811 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN812 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN813 = io_x[11] ? _GEN812 : _GEN811;
wire  _GEN814 = io_x[3] ? _GEN813 : _GEN810;
wire  _GEN815 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN816 = io_x[11] ? _GEN815 : _GEN214;
wire  _GEN817 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN818 = io_x[3] ? _GEN817 : _GEN816;
wire  _GEN819 = io_x[7] ? _GEN818 : _GEN814;
wire  _GEN820 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN821 = io_x[3] ? _GEN216 : _GEN820;
wire  _GEN822 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN823 = io_x[11] ? _GEN822 : _GEN207;
wire  _GEN824 = io_x[3] ? _GEN823 : _GEN216;
wire  _GEN825 = io_x[7] ? _GEN824 : _GEN821;
wire  _GEN826 = io_x[2] ? _GEN825 : _GEN819;
wire  _GEN827 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN828 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN829 = io_x[11] ? _GEN828 : _GEN827;
wire  _GEN830 = io_x[3] ? _GEN829 : _GEN209;
wire  _GEN831 = io_x[11] ? _GEN815 : _GEN214;
wire  _GEN832 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN833 = io_x[11] ? _GEN832 : _GEN207;
wire  _GEN834 = io_x[3] ? _GEN833 : _GEN831;
wire  _GEN835 = io_x[7] ? _GEN834 : _GEN830;
wire  _GEN836 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN837 = io_x[11] ? _GEN207 : _GEN836;
wire  _GEN838 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN839 = io_x[11] ? _GEN838 : _GEN214;
wire  _GEN840 = io_x[3] ? _GEN839 : _GEN837;
wire  _GEN841 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN842 = io_x[11] ? _GEN841 : _GEN214;
wire  _GEN843 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN844 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN845 = io_x[11] ? _GEN844 : _GEN843;
wire  _GEN846 = io_x[3] ? _GEN845 : _GEN842;
wire  _GEN847 = io_x[7] ? _GEN846 : _GEN840;
wire  _GEN848 = io_x[2] ? _GEN847 : _GEN835;
wire  _GEN849 = io_x[17] ? _GEN848 : _GEN826;
wire  _GEN850 = io_x[15] ? _GEN849 : _GEN808;
wire  _GEN851 = io_x[12] ? _GEN850 : _GEN777;
wire  _GEN852 = io_x[10] ? _GEN851 : _GEN737;
wire  _GEN853 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN854 = io_x[11] ? _GEN853 : _GEN214;
wire  _GEN855 = io_x[3] ? _GEN854 : _GEN216;
wire  _GEN856 = io_x[7] ? _GEN855 : _GEN241;
wire  _GEN857 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN858 = io_x[11] ? _GEN857 : _GEN214;
wire  _GEN859 = io_x[3] ? _GEN216 : _GEN858;
wire  _GEN860 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN861 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN862 = io_x[11] ? _GEN861 : _GEN214;
wire  _GEN863 = io_x[3] ? _GEN862 : _GEN860;
wire  _GEN864 = io_x[7] ? _GEN863 : _GEN859;
wire  _GEN865 = io_x[2] ? _GEN864 : _GEN856;
wire  _GEN866 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN867 = io_x[11] ? _GEN866 : _GEN207;
wire  _GEN868 = io_x[3] ? _GEN216 : _GEN867;
wire  _GEN869 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN870 = io_x[11] ? _GEN869 : _GEN214;
wire  _GEN871 = io_x[3] ? _GEN870 : _GEN216;
wire  _GEN872 = io_x[7] ? _GEN871 : _GEN868;
wire  _GEN873 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN874 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN875 = io_x[11] ? _GEN874 : _GEN214;
wire  _GEN876 = io_x[3] ? _GEN875 : _GEN209;
wire  _GEN877 = io_x[7] ? _GEN876 : _GEN873;
wire  _GEN878 = io_x[2] ? _GEN877 : _GEN872;
wire  _GEN879 = io_x[17] ? _GEN878 : _GEN865;
wire  _GEN880 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN881 = io_x[3] ? _GEN209 : _GEN880;
wire  _GEN882 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN883 = io_x[3] ? _GEN216 : _GEN882;
wire  _GEN884 = io_x[7] ? _GEN883 : _GEN881;
wire  _GEN885 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN886 = io_x[11] ? _GEN885 : _GEN214;
wire  _GEN887 = io_x[3] ? _GEN216 : _GEN886;
wire  _GEN888 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN889 = io_x[7] ? _GEN888 : _GEN887;
wire  _GEN890 = io_x[2] ? _GEN889 : _GEN884;
wire  _GEN891 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN892 = io_x[11] ? _GEN891 : _GEN214;
wire  _GEN893 = io_x[3] ? _GEN209 : _GEN892;
wire  _GEN894 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN895 = io_x[11] ? _GEN894 : _GEN214;
wire  _GEN896 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN897 = io_x[11] ? _GEN896 : _GEN214;
wire  _GEN898 = io_x[3] ? _GEN897 : _GEN895;
wire  _GEN899 = io_x[7] ? _GEN898 : _GEN893;
wire  _GEN900 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN901 = io_x[11] ? _GEN900 : _GEN214;
wire  _GEN902 = io_x[3] ? _GEN216 : _GEN901;
wire  _GEN903 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN904 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN905 = io_x[11] ? _GEN904 : _GEN903;
wire  _GEN906 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN907 = io_x[11] ? _GEN906 : _GEN214;
wire  _GEN908 = io_x[3] ? _GEN907 : _GEN905;
wire  _GEN909 = io_x[7] ? _GEN908 : _GEN902;
wire  _GEN910 = io_x[2] ? _GEN909 : _GEN899;
wire  _GEN911 = io_x[17] ? _GEN910 : _GEN890;
wire  _GEN912 = io_x[15] ? _GEN911 : _GEN879;
wire  _GEN913 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN914 = io_x[3] ? _GEN913 : _GEN216;
wire  _GEN915 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN916 = io_x[11] ? _GEN915 : _GEN214;
wire  _GEN917 = io_x[3] ? _GEN216 : _GEN916;
wire  _GEN918 = io_x[7] ? _GEN917 : _GEN914;
wire  _GEN919 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN920 = io_x[11] ? _GEN919 : _GEN214;
wire  _GEN921 = io_x[3] ? _GEN920 : _GEN216;
wire  _GEN922 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN923 = io_x[3] ? _GEN922 : _GEN209;
wire  _GEN924 = io_x[7] ? _GEN923 : _GEN921;
wire  _GEN925 = io_x[2] ? _GEN924 : _GEN918;
wire  _GEN926 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN927 = io_x[3] ? _GEN926 : _GEN216;
wire  _GEN928 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN929 = io_x[11] ? _GEN928 : _GEN214;
wire  _GEN930 = io_x[3] ? _GEN929 : _GEN209;
wire  _GEN931 = io_x[7] ? _GEN930 : _GEN927;
wire  _GEN932 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN933 = io_x[11] ? _GEN932 : _GEN207;
wire  _GEN934 = io_x[3] ? _GEN933 : _GEN216;
wire  _GEN935 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN936 = io_x[11] ? _GEN935 : _GEN214;
wire  _GEN937 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN938 = io_x[11] ? _GEN937 : _GEN207;
wire  _GEN939 = io_x[3] ? _GEN938 : _GEN936;
wire  _GEN940 = io_x[7] ? _GEN939 : _GEN934;
wire  _GEN941 = io_x[2] ? _GEN940 : _GEN931;
wire  _GEN942 = io_x[17] ? _GEN941 : _GEN925;
wire  _GEN943 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN944 = io_x[11] ? _GEN214 : _GEN943;
wire  _GEN945 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN946 = io_x[3] ? _GEN945 : _GEN944;
wire  _GEN947 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN948 = io_x[11] ? _GEN947 : _GEN214;
wire  _GEN949 = io_x[3] ? _GEN209 : _GEN948;
wire  _GEN950 = io_x[7] ? _GEN949 : _GEN946;
wire  _GEN951 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN952 = io_x[11] ? _GEN207 : _GEN951;
wire  _GEN953 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN954 = io_x[11] ? _GEN953 : _GEN214;
wire  _GEN955 = io_x[3] ? _GEN954 : _GEN952;
wire  _GEN956 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN957 = io_x[11] ? _GEN207 : _GEN956;
wire  _GEN958 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN959 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN960 = io_x[11] ? _GEN959 : _GEN958;
wire  _GEN961 = io_x[3] ? _GEN960 : _GEN957;
wire  _GEN962 = io_x[7] ? _GEN961 : _GEN955;
wire  _GEN963 = io_x[2] ? _GEN962 : _GEN950;
wire  _GEN964 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN965 = io_x[11] ? _GEN214 : _GEN964;
wire  _GEN966 = io_x[3] ? _GEN965 : _GEN216;
wire  _GEN967 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN968 = io_x[11] ? _GEN967 : _GEN214;
wire  _GEN969 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN970 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN971 = io_x[11] ? _GEN970 : _GEN969;
wire  _GEN972 = io_x[3] ? _GEN971 : _GEN968;
wire  _GEN973 = io_x[7] ? _GEN972 : _GEN966;
wire  _GEN974 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN975 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN976 = io_x[11] ? _GEN975 : _GEN974;
wire  _GEN977 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN978 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN979 = io_x[11] ? _GEN978 : _GEN977;
wire  _GEN980 = io_x[3] ? _GEN979 : _GEN976;
wire  _GEN981 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN982 = io_x[11] ? _GEN981 : _GEN214;
wire  _GEN983 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN984 = io_x[11] ? _GEN983 : _GEN214;
wire  _GEN985 = io_x[3] ? _GEN984 : _GEN982;
wire  _GEN986 = io_x[7] ? _GEN985 : _GEN980;
wire  _GEN987 = io_x[2] ? _GEN986 : _GEN973;
wire  _GEN988 = io_x[17] ? _GEN987 : _GEN963;
wire  _GEN989 = io_x[15] ? _GEN988 : _GEN942;
wire  _GEN990 = io_x[12] ? _GEN989 : _GEN912;
wire  _GEN991 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN992 = io_x[11] ? _GEN991 : _GEN214;
wire  _GEN993 = io_x[3] ? _GEN992 : _GEN216;
wire  _GEN994 = io_x[7] ? _GEN993 : _GEN203;
wire  _GEN995 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN996 = io_x[11] ? _GEN995 : _GEN214;
wire  _GEN997 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN998 = io_x[11] ? _GEN997 : _GEN214;
wire  _GEN999 = io_x[3] ? _GEN998 : _GEN996;
wire  _GEN1000 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1001 = io_x[11] ? _GEN207 : _GEN1000;
wire  _GEN1002 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1003 = io_x[3] ? _GEN1002 : _GEN1001;
wire  _GEN1004 = io_x[7] ? _GEN1003 : _GEN999;
wire  _GEN1005 = io_x[2] ? _GEN1004 : _GEN994;
wire  _GEN1006 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1007 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1008 = io_x[11] ? _GEN1007 : _GEN1006;
wire  _GEN1009 = io_x[3] ? _GEN1008 : _GEN209;
wire  _GEN1010 = io_x[7] ? _GEN241 : _GEN1009;
wire  _GEN1011 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1012 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1013 = io_x[11] ? _GEN1012 : _GEN1011;
wire  _GEN1014 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1015 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1016 = io_x[11] ? _GEN1015 : _GEN1014;
wire  _GEN1017 = io_x[3] ? _GEN1016 : _GEN1013;
wire  _GEN1018 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1019 = io_x[11] ? _GEN207 : _GEN1018;
wire  _GEN1020 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1021 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1022 = io_x[11] ? _GEN1021 : _GEN1020;
wire  _GEN1023 = io_x[3] ? _GEN1022 : _GEN1019;
wire  _GEN1024 = io_x[7] ? _GEN1023 : _GEN1017;
wire  _GEN1025 = io_x[2] ? _GEN1024 : _GEN1010;
wire  _GEN1026 = io_x[17] ? _GEN1025 : _GEN1005;
wire  _GEN1027 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1028 = io_x[11] ? _GEN207 : _GEN1027;
wire  _GEN1029 = io_x[3] ? _GEN1028 : _GEN216;
wire  _GEN1030 = io_x[7] ? _GEN203 : _GEN1029;
wire  _GEN1031 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1032 = io_x[11] ? _GEN1031 : _GEN214;
wire  _GEN1033 = io_x[3] ? _GEN1032 : _GEN216;
wire  _GEN1034 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1035 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1036 = io_x[11] ? _GEN1035 : _GEN207;
wire  _GEN1037 = io_x[3] ? _GEN1036 : _GEN1034;
wire  _GEN1038 = io_x[7] ? _GEN1037 : _GEN1033;
wire  _GEN1039 = io_x[2] ? _GEN1038 : _GEN1030;
wire  _GEN1040 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1041 = io_x[11] ? _GEN1040 : _GEN214;
wire  _GEN1042 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1043 = io_x[11] ? _GEN207 : _GEN1042;
wire  _GEN1044 = io_x[3] ? _GEN1043 : _GEN1041;
wire  _GEN1045 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1046 = io_x[11] ? _GEN1045 : _GEN214;
wire  _GEN1047 = io_x[3] ? _GEN1046 : _GEN209;
wire  _GEN1048 = io_x[7] ? _GEN1047 : _GEN1044;
wire  _GEN1049 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1050 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1051 = io_x[11] ? _GEN1050 : _GEN1049;
wire  _GEN1052 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1053 = io_x[11] ? _GEN1052 : _GEN214;
wire  _GEN1054 = io_x[3] ? _GEN1053 : _GEN1051;
wire  _GEN1055 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1056 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1057 = io_x[11] ? _GEN1056 : _GEN1055;
wire  _GEN1058 = io_x[3] ? _GEN1057 : _GEN216;
wire  _GEN1059 = io_x[7] ? _GEN1058 : _GEN1054;
wire  _GEN1060 = io_x[2] ? _GEN1059 : _GEN1048;
wire  _GEN1061 = io_x[17] ? _GEN1060 : _GEN1039;
wire  _GEN1062 = io_x[15] ? _GEN1061 : _GEN1026;
wire  _GEN1063 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1064 = io_x[11] ? _GEN1063 : _GEN207;
wire  _GEN1065 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1066 = io_x[11] ? _GEN214 : _GEN1065;
wire  _GEN1067 = io_x[3] ? _GEN1066 : _GEN1064;
wire  _GEN1068 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1069 = io_x[11] ? _GEN1068 : _GEN214;
wire  _GEN1070 = io_x[3] ? _GEN216 : _GEN1069;
wire  _GEN1071 = io_x[7] ? _GEN1070 : _GEN1067;
wire  _GEN1072 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1073 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1074 = io_x[11] ? _GEN1073 : _GEN1072;
wire  _GEN1075 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1076 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1077 = io_x[11] ? _GEN1076 : _GEN1075;
wire  _GEN1078 = io_x[3] ? _GEN1077 : _GEN1074;
wire  _GEN1079 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1080 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1081 = io_x[11] ? _GEN1080 : _GEN1079;
wire  _GEN1082 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1083 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1084 = io_x[11] ? _GEN1083 : _GEN1082;
wire  _GEN1085 = io_x[3] ? _GEN1084 : _GEN1081;
wire  _GEN1086 = io_x[7] ? _GEN1085 : _GEN1078;
wire  _GEN1087 = io_x[2] ? _GEN1086 : _GEN1071;
wire  _GEN1088 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1089 = io_x[11] ? _GEN1088 : _GEN207;
wire  _GEN1090 = io_x[3] ? _GEN1089 : _GEN209;
wire  _GEN1091 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1092 = io_x[3] ? _GEN1091 : _GEN216;
wire  _GEN1093 = io_x[7] ? _GEN1092 : _GEN1090;
wire  _GEN1094 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1095 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1096 = io_x[11] ? _GEN1095 : _GEN1094;
wire  _GEN1097 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1098 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1099 = io_x[11] ? _GEN1098 : _GEN1097;
wire  _GEN1100 = io_x[3] ? _GEN1099 : _GEN1096;
wire  _GEN1101 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1102 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1103 = io_x[11] ? _GEN1102 : _GEN1101;
wire  _GEN1104 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1105 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1106 = io_x[11] ? _GEN1105 : _GEN1104;
wire  _GEN1107 = io_x[3] ? _GEN1106 : _GEN1103;
wire  _GEN1108 = io_x[7] ? _GEN1107 : _GEN1100;
wire  _GEN1109 = io_x[2] ? _GEN1108 : _GEN1093;
wire  _GEN1110 = io_x[17] ? _GEN1109 : _GEN1087;
wire  _GEN1111 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1112 = io_x[11] ? _GEN1111 : _GEN214;
wire  _GEN1113 = io_x[3] ? _GEN1112 : _GEN216;
wire  _GEN1114 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1115 = io_x[11] ? _GEN1114 : _GEN214;
wire  _GEN1116 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1117 = io_x[11] ? _GEN1116 : _GEN214;
wire  _GEN1118 = io_x[3] ? _GEN1117 : _GEN1115;
wire  _GEN1119 = io_x[7] ? _GEN1118 : _GEN1113;
wire  _GEN1120 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1121 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1122 = io_x[11] ? _GEN1121 : _GEN1120;
wire  _GEN1123 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1124 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1125 = io_x[11] ? _GEN1124 : _GEN1123;
wire  _GEN1126 = io_x[3] ? _GEN1125 : _GEN1122;
wire  _GEN1127 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1128 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1129 = io_x[11] ? _GEN1128 : _GEN1127;
wire  _GEN1130 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1131 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1132 = io_x[11] ? _GEN1131 : _GEN1130;
wire  _GEN1133 = io_x[3] ? _GEN1132 : _GEN1129;
wire  _GEN1134 = io_x[7] ? _GEN1133 : _GEN1126;
wire  _GEN1135 = io_x[2] ? _GEN1134 : _GEN1119;
wire  _GEN1136 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1137 = io_x[11] ? _GEN1136 : _GEN214;
wire  _GEN1138 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1139 = io_x[3] ? _GEN1138 : _GEN1137;
wire  _GEN1140 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1141 = io_x[11] ? _GEN1140 : _GEN207;
wire  _GEN1142 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1143 = io_x[11] ? _GEN1142 : _GEN214;
wire  _GEN1144 = io_x[3] ? _GEN1143 : _GEN1141;
wire  _GEN1145 = io_x[7] ? _GEN1144 : _GEN1139;
wire  _GEN1146 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1147 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1148 = io_x[11] ? _GEN1147 : _GEN1146;
wire  _GEN1149 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1150 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1151 = io_x[11] ? _GEN1150 : _GEN1149;
wire  _GEN1152 = io_x[3] ? _GEN1151 : _GEN1148;
wire  _GEN1153 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1154 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1155 = io_x[11] ? _GEN1154 : _GEN1153;
wire  _GEN1156 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1157 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1158 = io_x[11] ? _GEN1157 : _GEN1156;
wire  _GEN1159 = io_x[3] ? _GEN1158 : _GEN1155;
wire  _GEN1160 = io_x[7] ? _GEN1159 : _GEN1152;
wire  _GEN1161 = io_x[2] ? _GEN1160 : _GEN1145;
wire  _GEN1162 = io_x[17] ? _GEN1161 : _GEN1135;
wire  _GEN1163 = io_x[15] ? _GEN1162 : _GEN1110;
wire  _GEN1164 = io_x[12] ? _GEN1163 : _GEN1062;
wire  _GEN1165 = io_x[10] ? _GEN1164 : _GEN990;
wire  _GEN1166 = io_x[4] ? _GEN1165 : _GEN852;
wire  _GEN1167 = io_x[8] ? _GEN1166 : _GEN631;
wire  _GEN1168 = io_x[2] ? _GEN233 : _GEN202;
wire  _GEN1169 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1170 = io_x[11] ? _GEN1169 : _GEN214;
wire  _GEN1171 = io_x[3] ? _GEN1170 : _GEN216;
wire  _GEN1172 = io_x[7] ? _GEN1171 : _GEN241;
wire  _GEN1173 = io_x[2] ? _GEN233 : _GEN1172;
wire  _GEN1174 = io_x[17] ? _GEN1173 : _GEN1168;
wire  _GEN1175 = io_x[7] ? _GEN203 : _GEN241;
wire  _GEN1176 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1177 = io_x[11] ? _GEN1176 : _GEN214;
wire  _GEN1178 = io_x[3] ? _GEN1177 : _GEN209;
wire  _GEN1179 = io_x[7] ? _GEN1178 : _GEN203;
wire  _GEN1180 = io_x[2] ? _GEN1179 : _GEN1175;
wire  _GEN1181 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1182 = io_x[3] ? _GEN1181 : _GEN216;
wire  _GEN1183 = io_x[7] ? _GEN203 : _GEN1182;
wire  _GEN1184 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1185 = io_x[11] ? _GEN1184 : _GEN214;
wire  _GEN1186 = io_x[3] ? _GEN1185 : _GEN216;
wire  _GEN1187 = io_x[7] ? _GEN1186 : _GEN203;
wire  _GEN1188 = io_x[2] ? _GEN1187 : _GEN1183;
wire  _GEN1189 = io_x[17] ? _GEN1188 : _GEN1180;
wire  _GEN1190 = io_x[15] ? _GEN1189 : _GEN1174;
wire  _GEN1191 = io_x[7] ? _GEN203 : _GEN241;
wire  _GEN1192 = io_x[2] ? _GEN1191 : _GEN202;
wire  _GEN1193 = io_x[7] ? _GEN203 : _GEN241;
wire  _GEN1194 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1195 = io_x[3] ? _GEN1194 : _GEN216;
wire  _GEN1196 = io_x[7] ? _GEN1195 : _GEN203;
wire  _GEN1197 = io_x[2] ? _GEN1196 : _GEN1193;
wire  _GEN1198 = io_x[17] ? _GEN1197 : _GEN1192;
wire  _GEN1199 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1200 = io_x[3] ? _GEN1199 : _GEN216;
wire  _GEN1201 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1202 = io_x[3] ? _GEN1201 : _GEN216;
wire  _GEN1203 = io_x[7] ? _GEN1202 : _GEN1200;
wire  _GEN1204 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1205 = io_x[7] ? _GEN241 : _GEN1204;
wire  _GEN1206 = io_x[2] ? _GEN1205 : _GEN1203;
wire  _GEN1207 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1208 = io_x[3] ? _GEN1207 : _GEN216;
wire  _GEN1209 = io_x[7] ? _GEN203 : _GEN1208;
wire  _GEN1210 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1211 = io_x[7] ? _GEN241 : _GEN1210;
wire  _GEN1212 = io_x[2] ? _GEN1211 : _GEN1209;
wire  _GEN1213 = io_x[17] ? _GEN1212 : _GEN1206;
wire  _GEN1214 = io_x[15] ? _GEN1213 : _GEN1198;
wire  _GEN1215 = io_x[12] ? _GEN1214 : _GEN1190;
wire  _GEN1216 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1217 = io_x[3] ? _GEN1216 : _GEN216;
wire  _GEN1218 = io_x[7] ? _GEN1217 : _GEN241;
wire  _GEN1219 = io_x[2] ? _GEN1218 : _GEN233;
wire  _GEN1220 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1221 = io_x[3] ? _GEN1220 : _GEN216;
wire  _GEN1222 = io_x[7] ? _GEN1221 : _GEN203;
wire  _GEN1223 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1224 = io_x[11] ? _GEN1223 : _GEN207;
wire  _GEN1225 = io_x[3] ? _GEN1224 : _GEN216;
wire  _GEN1226 = io_x[7] ? _GEN1225 : _GEN241;
wire  _GEN1227 = io_x[2] ? _GEN1226 : _GEN1222;
wire  _GEN1228 = io_x[17] ? _GEN1227 : _GEN1219;
wire  _GEN1229 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1230 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1231 = io_x[11] ? _GEN1230 : _GEN1229;
wire  _GEN1232 = io_x[3] ? _GEN1231 : _GEN216;
wire  _GEN1233 = io_x[7] ? _GEN1232 : _GEN203;
wire  _GEN1234 = io_x[2] ? _GEN1233 : _GEN202;
wire  _GEN1235 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN1236 = io_x[7] ? _GEN1235 : _GEN203;
wire  _GEN1237 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1238 = io_x[3] ? _GEN216 : _GEN1237;
wire  _GEN1239 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1240 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1241 = io_x[11] ? _GEN1240 : _GEN214;
wire  _GEN1242 = io_x[3] ? _GEN1241 : _GEN1239;
wire  _GEN1243 = io_x[7] ? _GEN1242 : _GEN1238;
wire  _GEN1244 = io_x[2] ? _GEN1243 : _GEN1236;
wire  _GEN1245 = io_x[17] ? _GEN1244 : _GEN1234;
wire  _GEN1246 = io_x[15] ? _GEN1245 : _GEN1228;
wire  _GEN1247 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1248 = io_x[3] ? _GEN1247 : _GEN216;
wire  _GEN1249 = io_x[7] ? _GEN203 : _GEN1248;
wire  _GEN1250 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1251 = io_x[11] ? _GEN214 : _GEN1250;
wire  _GEN1252 = io_x[3] ? _GEN1251 : _GEN216;
wire  _GEN1253 = io_x[7] ? _GEN1252 : _GEN203;
wire  _GEN1254 = io_x[2] ? _GEN1253 : _GEN1249;
wire  _GEN1255 = io_x[2] ? _GEN202 : _GEN233;
wire  _GEN1256 = io_x[17] ? _GEN1255 : _GEN1254;
wire  _GEN1257 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1258 = io_x[7] ? _GEN1257 : _GEN203;
wire  _GEN1259 = io_x[2] ? _GEN1258 : _GEN233;
wire  _GEN1260 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1261 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1262 = io_x[11] ? _GEN214 : _GEN1261;
wire  _GEN1263 = io_x[3] ? _GEN1262 : _GEN216;
wire  _GEN1264 = io_x[7] ? _GEN1263 : _GEN1260;
wire  _GEN1265 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1266 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1267 = io_x[11] ? _GEN1266 : _GEN1265;
wire  _GEN1268 = io_x[3] ? _GEN1267 : _GEN216;
wire  _GEN1269 = io_x[7] ? _GEN1268 : _GEN203;
wire  _GEN1270 = io_x[2] ? _GEN1269 : _GEN1264;
wire  _GEN1271 = io_x[17] ? _GEN1270 : _GEN1259;
wire  _GEN1272 = io_x[15] ? _GEN1271 : _GEN1256;
wire  _GEN1273 = io_x[12] ? _GEN1272 : _GEN1246;
wire  _GEN1274 = io_x[10] ? _GEN1273 : _GEN1215;
wire  _GEN1275 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1276 = io_x[3] ? _GEN1275 : _GEN216;
wire  _GEN1277 = io_x[7] ? _GEN1276 : _GEN203;
wire  _GEN1278 = io_x[2] ? _GEN202 : _GEN1277;
wire  _GEN1279 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1280 = io_x[7] ? _GEN1279 : _GEN203;
wire  _GEN1281 = io_x[2] ? _GEN1280 : _GEN233;
wire  _GEN1282 = io_x[17] ? _GEN1281 : _GEN1278;
wire  _GEN1283 = 1'b0;
wire  _GEN1284 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1285 = io_x[11] ? _GEN1284 : _GEN214;
wire  _GEN1286 = io_x[3] ? _GEN1285 : _GEN209;
wire  _GEN1287 = io_x[7] ? _GEN1286 : _GEN241;
wire  _GEN1288 = io_x[2] ? _GEN1287 : _GEN233;
wire  _GEN1289 = io_x[17] ? _GEN1288 : _GEN1283;
wire  _GEN1290 = io_x[15] ? _GEN1289 : _GEN1282;
wire  _GEN1291 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1292 = io_x[3] ? _GEN216 : _GEN1291;
wire  _GEN1293 = io_x[7] ? _GEN1292 : _GEN203;
wire  _GEN1294 = io_x[2] ? _GEN233 : _GEN1293;
wire  _GEN1295 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1296 = io_x[3] ? _GEN209 : _GEN1295;
wire  _GEN1297 = io_x[7] ? _GEN1296 : _GEN203;
wire  _GEN1298 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN1299 = io_x[2] ? _GEN1298 : _GEN1297;
wire  _GEN1300 = io_x[17] ? _GEN1299 : _GEN1294;
wire  _GEN1301 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1302 = io_x[11] ? _GEN1301 : _GEN207;
wire  _GEN1303 = io_x[3] ? _GEN216 : _GEN1302;
wire  _GEN1304 = io_x[7] ? _GEN1303 : _GEN203;
wire  _GEN1305 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1306 = io_x[3] ? _GEN1305 : _GEN216;
wire  _GEN1307 = io_x[7] ? _GEN1306 : _GEN241;
wire  _GEN1308 = io_x[2] ? _GEN1307 : _GEN1304;
wire  _GEN1309 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1310 = io_x[3] ? _GEN216 : _GEN1309;
wire  _GEN1311 = io_x[7] ? _GEN1310 : _GEN203;
wire  _GEN1312 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1313 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1314 = io_x[11] ? _GEN1313 : _GEN1312;
wire  _GEN1315 = io_x[3] ? _GEN1314 : _GEN216;
wire  _GEN1316 = io_x[7] ? _GEN1315 : _GEN241;
wire  _GEN1317 = io_x[2] ? _GEN1316 : _GEN1311;
wire  _GEN1318 = io_x[17] ? _GEN1317 : _GEN1308;
wire  _GEN1319 = io_x[15] ? _GEN1318 : _GEN1300;
wire  _GEN1320 = io_x[12] ? _GEN1319 : _GEN1290;
wire  _GEN1321 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1322 = io_x[11] ? _GEN207 : _GEN1321;
wire  _GEN1323 = io_x[3] ? _GEN216 : _GEN1322;
wire  _GEN1324 = io_x[7] ? _GEN1323 : _GEN203;
wire  _GEN1325 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1326 = io_x[11] ? _GEN1325 : _GEN207;
wire  _GEN1327 = io_x[3] ? _GEN1326 : _GEN216;
wire  _GEN1328 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1329 = io_x[11] ? _GEN1328 : _GEN214;
wire  _GEN1330 = io_x[3] ? _GEN1329 : _GEN216;
wire  _GEN1331 = io_x[7] ? _GEN1330 : _GEN1327;
wire  _GEN1332 = io_x[2] ? _GEN1331 : _GEN1324;
wire  _GEN1333 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1334 = io_x[11] ? _GEN214 : _GEN1333;
wire  _GEN1335 = io_x[3] ? _GEN1334 : _GEN216;
wire  _GEN1336 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1337 = io_x[11] ? _GEN207 : _GEN1336;
wire  _GEN1338 = io_x[3] ? _GEN216 : _GEN1337;
wire  _GEN1339 = io_x[7] ? _GEN1338 : _GEN1335;
wire  _GEN1340 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1341 = io_x[11] ? _GEN1340 : _GEN214;
wire  _GEN1342 = io_x[3] ? _GEN1341 : _GEN216;
wire  _GEN1343 = io_x[7] ? _GEN203 : _GEN1342;
wire  _GEN1344 = io_x[2] ? _GEN1343 : _GEN1339;
wire  _GEN1345 = io_x[17] ? _GEN1344 : _GEN1332;
wire  _GEN1346 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN1347 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1348 = io_x[11] ? _GEN1347 : _GEN214;
wire  _GEN1349 = io_x[3] ? _GEN1348 : _GEN216;
wire  _GEN1350 = io_x[7] ? _GEN1349 : _GEN203;
wire  _GEN1351 = io_x[2] ? _GEN1350 : _GEN1346;
wire  _GEN1352 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1353 = io_x[3] ? _GEN209 : _GEN1352;
wire  _GEN1354 = io_x[7] ? _GEN1353 : _GEN203;
wire  _GEN1355 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1356 = io_x[11] ? _GEN1355 : _GEN214;
wire  _GEN1357 = io_x[3] ? _GEN1356 : _GEN216;
wire  _GEN1358 = io_x[7] ? _GEN1357 : _GEN203;
wire  _GEN1359 = io_x[2] ? _GEN1358 : _GEN1354;
wire  _GEN1360 = io_x[17] ? _GEN1359 : _GEN1351;
wire  _GEN1361 = io_x[15] ? _GEN1360 : _GEN1345;
wire  _GEN1362 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1363 = io_x[7] ? _GEN1362 : _GEN203;
wire  _GEN1364 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN1365 = io_x[2] ? _GEN1364 : _GEN1363;
wire  _GEN1366 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1367 = io_x[7] ? _GEN1366 : _GEN203;
wire  _GEN1368 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1369 = io_x[11] ? _GEN207 : _GEN1368;
wire  _GEN1370 = io_x[3] ? _GEN1369 : _GEN216;
wire  _GEN1371 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1372 = io_x[3] ? _GEN1371 : _GEN216;
wire  _GEN1373 = io_x[7] ? _GEN1372 : _GEN1370;
wire  _GEN1374 = io_x[2] ? _GEN1373 : _GEN1367;
wire  _GEN1375 = io_x[17] ? _GEN1374 : _GEN1365;
wire  _GEN1376 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN1377 = io_x[7] ? _GEN1376 : _GEN203;
wire  _GEN1378 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1379 = io_x[11] ? _GEN1378 : _GEN207;
wire  _GEN1380 = io_x[3] ? _GEN209 : _GEN1379;
wire  _GEN1381 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1382 = io_x[11] ? _GEN1381 : _GEN214;
wire  _GEN1383 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1384 = io_x[11] ? _GEN1383 : _GEN214;
wire  _GEN1385 = io_x[3] ? _GEN1384 : _GEN1382;
wire  _GEN1386 = io_x[7] ? _GEN1385 : _GEN1380;
wire  _GEN1387 = io_x[2] ? _GEN1386 : _GEN1377;
wire  _GEN1388 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN1389 = io_x[7] ? _GEN1388 : _GEN203;
wire  _GEN1390 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1391 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1392 = io_x[11] ? _GEN1391 : _GEN1390;
wire  _GEN1393 = io_x[3] ? _GEN1392 : _GEN216;
wire  _GEN1394 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1395 = io_x[11] ? _GEN1394 : _GEN214;
wire  _GEN1396 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1397 = io_x[11] ? _GEN1396 : _GEN214;
wire  _GEN1398 = io_x[3] ? _GEN1397 : _GEN1395;
wire  _GEN1399 = io_x[7] ? _GEN1398 : _GEN1393;
wire  _GEN1400 = io_x[2] ? _GEN1399 : _GEN1389;
wire  _GEN1401 = io_x[17] ? _GEN1400 : _GEN1387;
wire  _GEN1402 = io_x[15] ? _GEN1401 : _GEN1375;
wire  _GEN1403 = io_x[12] ? _GEN1402 : _GEN1361;
wire  _GEN1404 = io_x[10] ? _GEN1403 : _GEN1320;
wire  _GEN1405 = io_x[4] ? _GEN1404 : _GEN1274;
wire  _GEN1406 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1407 = io_x[11] ? _GEN1406 : _GEN214;
wire  _GEN1408 = io_x[3] ? _GEN1407 : _GEN209;
wire  _GEN1409 = io_x[7] ? _GEN203 : _GEN1408;
wire  _GEN1410 = io_x[2] ? _GEN1409 : _GEN233;
wire  _GEN1411 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1412 = io_x[3] ? _GEN209 : _GEN1411;
wire  _GEN1413 = io_x[7] ? _GEN203 : _GEN1412;
wire  _GEN1414 = io_x[2] ? _GEN1413 : _GEN202;
wire  _GEN1415 = io_x[17] ? _GEN1414 : _GEN1410;
wire  _GEN1416 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN1417 = io_x[2] ? _GEN1416 : _GEN202;
wire  _GEN1418 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1419 = io_x[11] ? _GEN1418 : _GEN214;
wire  _GEN1420 = io_x[3] ? _GEN1419 : _GEN216;
wire  _GEN1421 = io_x[7] ? _GEN1420 : _GEN241;
wire  _GEN1422 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1423 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1424 = io_x[11] ? _GEN1423 : _GEN214;
wire  _GEN1425 = io_x[3] ? _GEN1424 : _GEN1422;
wire  _GEN1426 = io_x[7] ? _GEN241 : _GEN1425;
wire  _GEN1427 = io_x[2] ? _GEN1426 : _GEN1421;
wire  _GEN1428 = io_x[17] ? _GEN1427 : _GEN1417;
wire  _GEN1429 = io_x[15] ? _GEN1428 : _GEN1415;
wire  _GEN1430 = io_x[2] ? _GEN202 : _GEN233;
wire  _GEN1431 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1432 = io_x[11] ? _GEN1431 : _GEN214;
wire  _GEN1433 = io_x[3] ? _GEN1432 : _GEN209;
wire  _GEN1434 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1435 = io_x[3] ? _GEN1434 : _GEN216;
wire  _GEN1436 = io_x[7] ? _GEN1435 : _GEN1433;
wire  _GEN1437 = io_x[2] ? _GEN1436 : _GEN233;
wire  _GEN1438 = io_x[17] ? _GEN1437 : _GEN1430;
wire  _GEN1439 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1440 = io_x[7] ? _GEN203 : _GEN1439;
wire  _GEN1441 = io_x[2] ? _GEN1440 : _GEN202;
wire  _GEN1442 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1443 = io_x[11] ? _GEN1442 : _GEN214;
wire  _GEN1444 = io_x[3] ? _GEN1443 : _GEN216;
wire  _GEN1445 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1446 = io_x[3] ? _GEN1445 : _GEN216;
wire  _GEN1447 = io_x[7] ? _GEN1446 : _GEN1444;
wire  _GEN1448 = io_x[2] ? _GEN1447 : _GEN233;
wire  _GEN1449 = io_x[17] ? _GEN1448 : _GEN1441;
wire  _GEN1450 = io_x[15] ? _GEN1449 : _GEN1438;
wire  _GEN1451 = io_x[12] ? _GEN1450 : _GEN1429;
wire  _GEN1452 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN1453 = io_x[7] ? _GEN241 : _GEN1452;
wire  _GEN1454 = io_x[2] ? _GEN1453 : _GEN202;
wire  _GEN1455 = io_x[17] ? _GEN1283 : _GEN1454;
wire  _GEN1456 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1457 = io_x[3] ? _GEN1456 : _GEN216;
wire  _GEN1458 = io_x[7] ? _GEN1457 : _GEN203;
wire  _GEN1459 = io_x[2] ? _GEN1458 : _GEN233;
wire  _GEN1460 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1461 = io_x[3] ? _GEN1460 : _GEN216;
wire  _GEN1462 = io_x[7] ? _GEN1461 : _GEN203;
wire  _GEN1463 = io_x[2] ? _GEN1462 : _GEN202;
wire  _GEN1464 = io_x[17] ? _GEN1463 : _GEN1459;
wire  _GEN1465 = io_x[15] ? _GEN1464 : _GEN1455;
wire  _GEN1466 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1467 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1468 = io_x[11] ? _GEN1467 : _GEN214;
wire  _GEN1469 = io_x[3] ? _GEN1468 : _GEN216;
wire  _GEN1470 = io_x[7] ? _GEN1469 : _GEN1466;
wire  _GEN1471 = io_x[2] ? _GEN1470 : _GEN233;
wire  _GEN1472 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1473 = io_x[3] ? _GEN216 : _GEN1472;
wire  _GEN1474 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1475 = io_x[11] ? _GEN1474 : _GEN214;
wire  _GEN1476 = io_x[3] ? _GEN1475 : _GEN216;
wire  _GEN1477 = io_x[7] ? _GEN1476 : _GEN1473;
wire  _GEN1478 = io_x[2] ? _GEN1477 : _GEN233;
wire  _GEN1479 = io_x[17] ? _GEN1478 : _GEN1471;
wire  _GEN1480 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1481 = io_x[11] ? _GEN1480 : _GEN214;
wire  _GEN1482 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1483 = io_x[11] ? _GEN1482 : _GEN214;
wire  _GEN1484 = io_x[3] ? _GEN1483 : _GEN1481;
wire  _GEN1485 = io_x[7] ? _GEN1484 : _GEN241;
wire  _GEN1486 = io_x[2] ? _GEN202 : _GEN1485;
wire  _GEN1487 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1488 = io_x[11] ? _GEN1487 : _GEN214;
wire  _GEN1489 = io_x[3] ? _GEN216 : _GEN1488;
wire  _GEN1490 = io_x[7] ? _GEN1489 : _GEN241;
wire  _GEN1491 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1492 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1493 = io_x[11] ? _GEN1492 : _GEN1491;
wire  _GEN1494 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1495 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1496 = io_x[11] ? _GEN1495 : _GEN1494;
wire  _GEN1497 = io_x[3] ? _GEN1496 : _GEN1493;
wire  _GEN1498 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1499 = io_x[11] ? _GEN1498 : _GEN214;
wire  _GEN1500 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1501 = io_x[11] ? _GEN1500 : _GEN214;
wire  _GEN1502 = io_x[3] ? _GEN1501 : _GEN1499;
wire  _GEN1503 = io_x[7] ? _GEN1502 : _GEN1497;
wire  _GEN1504 = io_x[2] ? _GEN1503 : _GEN1490;
wire  _GEN1505 = io_x[17] ? _GEN1504 : _GEN1486;
wire  _GEN1506 = io_x[15] ? _GEN1505 : _GEN1479;
wire  _GEN1507 = io_x[12] ? _GEN1506 : _GEN1465;
wire  _GEN1508 = io_x[10] ? _GEN1507 : _GEN1451;
wire  _GEN1509 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1510 = io_x[3] ? _GEN216 : _GEN1509;
wire  _GEN1511 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1512 = io_x[7] ? _GEN1511 : _GEN1510;
wire  _GEN1513 = io_x[2] ? _GEN233 : _GEN1512;
wire  _GEN1514 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1515 = io_x[3] ? _GEN216 : _GEN1514;
wire  _GEN1516 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1517 = io_x[7] ? _GEN1516 : _GEN1515;
wire  _GEN1518 = io_x[2] ? _GEN202 : _GEN1517;
wire  _GEN1519 = io_x[17] ? _GEN1518 : _GEN1513;
wire  _GEN1520 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1521 = io_x[7] ? _GEN203 : _GEN1520;
wire  _GEN1522 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1523 = io_x[11] ? _GEN1522 : _GEN214;
wire  _GEN1524 = io_x[3] ? _GEN1523 : _GEN216;
wire  _GEN1525 = io_x[7] ? _GEN1524 : _GEN203;
wire  _GEN1526 = io_x[2] ? _GEN1525 : _GEN1521;
wire  _GEN1527 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1528 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1529 = io_x[11] ? _GEN1528 : _GEN214;
wire  _GEN1530 = io_x[3] ? _GEN1529 : _GEN216;
wire  _GEN1531 = io_x[7] ? _GEN1530 : _GEN1527;
wire  _GEN1532 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1533 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1534 = io_x[11] ? _GEN1533 : _GEN1532;
wire  _GEN1535 = io_x[3] ? _GEN1534 : _GEN209;
wire  _GEN1536 = io_x[7] ? _GEN1535 : _GEN203;
wire  _GEN1537 = io_x[2] ? _GEN1536 : _GEN1531;
wire  _GEN1538 = io_x[17] ? _GEN1537 : _GEN1526;
wire  _GEN1539 = io_x[15] ? _GEN1538 : _GEN1519;
wire  _GEN1540 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1541 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1542 = io_x[11] ? _GEN207 : _GEN1541;
wire  _GEN1543 = io_x[3] ? _GEN1542 : _GEN1540;
wire  _GEN1544 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1545 = io_x[7] ? _GEN1544 : _GEN1543;
wire  _GEN1546 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1547 = io_x[3] ? _GEN1546 : _GEN209;
wire  _GEN1548 = io_x[7] ? _GEN1547 : _GEN241;
wire  _GEN1549 = io_x[2] ? _GEN1548 : _GEN1545;
wire  _GEN1550 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1551 = io_x[11] ? _GEN214 : _GEN1550;
wire  _GEN1552 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1553 = io_x[3] ? _GEN1552 : _GEN1551;
wire  _GEN1554 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1555 = io_x[11] ? _GEN1554 : _GEN207;
wire  _GEN1556 = io_x[3] ? _GEN1555 : _GEN209;
wire  _GEN1557 = io_x[7] ? _GEN1556 : _GEN1553;
wire  _GEN1558 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1559 = io_x[11] ? _GEN1558 : _GEN214;
wire  _GEN1560 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1561 = io_x[11] ? _GEN1560 : _GEN214;
wire  _GEN1562 = io_x[3] ? _GEN1561 : _GEN1559;
wire  _GEN1563 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1564 = io_x[7] ? _GEN1563 : _GEN1562;
wire  _GEN1565 = io_x[2] ? _GEN1564 : _GEN1557;
wire  _GEN1566 = io_x[17] ? _GEN1565 : _GEN1549;
wire  _GEN1567 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1568 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1569 = io_x[11] ? _GEN1568 : _GEN214;
wire  _GEN1570 = io_x[3] ? _GEN1569 : _GEN216;
wire  _GEN1571 = io_x[7] ? _GEN1570 : _GEN1567;
wire  _GEN1572 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1573 = io_x[11] ? _GEN214 : _GEN1572;
wire  _GEN1574 = io_x[3] ? _GEN1573 : _GEN209;
wire  _GEN1575 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1576 = io_x[11] ? _GEN1575 : _GEN214;
wire  _GEN1577 = io_x[3] ? _GEN1576 : _GEN216;
wire  _GEN1578 = io_x[7] ? _GEN1577 : _GEN1574;
wire  _GEN1579 = io_x[2] ? _GEN1578 : _GEN1571;
wire  _GEN1580 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1581 = io_x[3] ? _GEN1580 : _GEN209;
wire  _GEN1582 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1583 = io_x[11] ? _GEN1582 : _GEN214;
wire  _GEN1584 = io_x[3] ? _GEN1583 : _GEN216;
wire  _GEN1585 = io_x[7] ? _GEN1584 : _GEN1581;
wire  _GEN1586 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1587 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1588 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1589 = io_x[11] ? _GEN1588 : _GEN1587;
wire  _GEN1590 = io_x[3] ? _GEN1589 : _GEN216;
wire  _GEN1591 = io_x[7] ? _GEN1590 : _GEN1586;
wire  _GEN1592 = io_x[2] ? _GEN1591 : _GEN1585;
wire  _GEN1593 = io_x[17] ? _GEN1592 : _GEN1579;
wire  _GEN1594 = io_x[15] ? _GEN1593 : _GEN1566;
wire  _GEN1595 = io_x[12] ? _GEN1594 : _GEN1539;
wire  _GEN1596 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1597 = io_x[11] ? _GEN1596 : _GEN214;
wire  _GEN1598 = io_x[3] ? _GEN1597 : _GEN216;
wire  _GEN1599 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1600 = io_x[3] ? _GEN1599 : _GEN216;
wire  _GEN1601 = io_x[7] ? _GEN1600 : _GEN1598;
wire  _GEN1602 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1603 = io_x[11] ? _GEN214 : _GEN1602;
wire  _GEN1604 = io_x[3] ? _GEN1603 : _GEN216;
wire  _GEN1605 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1606 = io_x[11] ? _GEN1605 : _GEN214;
wire  _GEN1607 = io_x[3] ? _GEN1606 : _GEN216;
wire  _GEN1608 = io_x[7] ? _GEN1607 : _GEN1604;
wire  _GEN1609 = io_x[2] ? _GEN1608 : _GEN1601;
wire  _GEN1610 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1611 = io_x[3] ? _GEN209 : _GEN1610;
wire  _GEN1612 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1613 = io_x[11] ? _GEN1612 : _GEN214;
wire  _GEN1614 = io_x[3] ? _GEN1613 : _GEN216;
wire  _GEN1615 = io_x[7] ? _GEN1614 : _GEN1611;
wire  _GEN1616 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1617 = io_x[11] ? _GEN207 : _GEN1616;
wire  _GEN1618 = io_x[3] ? _GEN1617 : _GEN216;
wire  _GEN1619 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1620 = io_x[11] ? _GEN1619 : _GEN214;
wire  _GEN1621 = io_x[3] ? _GEN1620 : _GEN216;
wire  _GEN1622 = io_x[7] ? _GEN1621 : _GEN1618;
wire  _GEN1623 = io_x[2] ? _GEN1622 : _GEN1615;
wire  _GEN1624 = io_x[17] ? _GEN1623 : _GEN1609;
wire  _GEN1625 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1626 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1627 = io_x[11] ? _GEN1626 : _GEN214;
wire  _GEN1628 = io_x[3] ? _GEN1627 : _GEN1625;
wire  _GEN1629 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1630 = io_x[11] ? _GEN1629 : _GEN214;
wire  _GEN1631 = io_x[3] ? _GEN1630 : _GEN216;
wire  _GEN1632 = io_x[7] ? _GEN1631 : _GEN1628;
wire  _GEN1633 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1634 = io_x[11] ? _GEN1633 : _GEN214;
wire  _GEN1635 = io_x[3] ? _GEN209 : _GEN1634;
wire  _GEN1636 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1637 = io_x[11] ? _GEN1636 : _GEN214;
wire  _GEN1638 = io_x[3] ? _GEN1637 : _GEN209;
wire  _GEN1639 = io_x[7] ? _GEN1638 : _GEN1635;
wire  _GEN1640 = io_x[2] ? _GEN1639 : _GEN1632;
wire  _GEN1641 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1642 = io_x[11] ? _GEN1641 : _GEN214;
wire  _GEN1643 = io_x[3] ? _GEN1642 : _GEN209;
wire  _GEN1644 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1645 = io_x[11] ? _GEN1644 : _GEN214;
wire  _GEN1646 = io_x[3] ? _GEN1645 : _GEN216;
wire  _GEN1647 = io_x[7] ? _GEN1646 : _GEN1643;
wire  _GEN1648 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN1649 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1650 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1651 = io_x[11] ? _GEN1650 : _GEN1649;
wire  _GEN1652 = io_x[3] ? _GEN1651 : _GEN216;
wire  _GEN1653 = io_x[7] ? _GEN1652 : _GEN1648;
wire  _GEN1654 = io_x[2] ? _GEN1653 : _GEN1647;
wire  _GEN1655 = io_x[17] ? _GEN1654 : _GEN1640;
wire  _GEN1656 = io_x[15] ? _GEN1655 : _GEN1624;
wire  _GEN1657 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1658 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1659 = io_x[11] ? _GEN207 : _GEN1658;
wire  _GEN1660 = io_x[3] ? _GEN1659 : _GEN1657;
wire  _GEN1661 = io_x[7] ? _GEN1660 : _GEN241;
wire  _GEN1662 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1663 = io_x[11] ? _GEN214 : _GEN1662;
wire  _GEN1664 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1665 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1666 = io_x[11] ? _GEN1665 : _GEN1664;
wire  _GEN1667 = io_x[3] ? _GEN1666 : _GEN1663;
wire  _GEN1668 = io_x[7] ? _GEN1667 : _GEN203;
wire  _GEN1669 = io_x[2] ? _GEN1668 : _GEN1661;
wire  _GEN1670 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1671 = io_x[3] ? _GEN209 : _GEN1670;
wire  _GEN1672 = io_x[7] ? _GEN241 : _GEN1671;
wire  _GEN1673 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1674 = io_x[11] ? _GEN214 : _GEN1673;
wire  _GEN1675 = io_x[3] ? _GEN1674 : _GEN216;
wire  _GEN1676 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1677 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1678 = io_x[11] ? _GEN1677 : _GEN1676;
wire  _GEN1679 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1680 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1681 = io_x[11] ? _GEN1680 : _GEN1679;
wire  _GEN1682 = io_x[3] ? _GEN1681 : _GEN1678;
wire  _GEN1683 = io_x[7] ? _GEN1682 : _GEN1675;
wire  _GEN1684 = io_x[2] ? _GEN1683 : _GEN1672;
wire  _GEN1685 = io_x[17] ? _GEN1684 : _GEN1669;
wire  _GEN1686 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1687 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1688 = io_x[3] ? _GEN1687 : _GEN1686;
wire  _GEN1689 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1690 = io_x[11] ? _GEN1689 : _GEN207;
wire  _GEN1691 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1692 = io_x[11] ? _GEN1691 : _GEN214;
wire  _GEN1693 = io_x[3] ? _GEN1692 : _GEN1690;
wire  _GEN1694 = io_x[7] ? _GEN1693 : _GEN1688;
wire  _GEN1695 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1696 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1697 = io_x[11] ? _GEN1696 : _GEN1695;
wire  _GEN1698 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1699 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1700 = io_x[11] ? _GEN1699 : _GEN1698;
wire  _GEN1701 = io_x[3] ? _GEN1700 : _GEN1697;
wire  _GEN1702 = io_x[7] ? _GEN1701 : _GEN241;
wire  _GEN1703 = io_x[2] ? _GEN1702 : _GEN1694;
wire  _GEN1704 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1705 = io_x[11] ? _GEN1704 : _GEN214;
wire  _GEN1706 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1707 = io_x[3] ? _GEN1706 : _GEN1705;
wire  _GEN1708 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1709 = io_x[11] ? _GEN1708 : _GEN207;
wire  _GEN1710 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1711 = io_x[11] ? _GEN1710 : _GEN214;
wire  _GEN1712 = io_x[3] ? _GEN1711 : _GEN1709;
wire  _GEN1713 = io_x[7] ? _GEN1712 : _GEN1707;
wire  _GEN1714 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1715 = io_x[11] ? _GEN1714 : _GEN207;
wire  _GEN1716 = io_x[3] ? _GEN1715 : _GEN209;
wire  _GEN1717 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1718 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1719 = io_x[11] ? _GEN1718 : _GEN1717;
wire  _GEN1720 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1721 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1722 = io_x[11] ? _GEN1721 : _GEN1720;
wire  _GEN1723 = io_x[3] ? _GEN1722 : _GEN1719;
wire  _GEN1724 = io_x[7] ? _GEN1723 : _GEN1716;
wire  _GEN1725 = io_x[2] ? _GEN1724 : _GEN1713;
wire  _GEN1726 = io_x[17] ? _GEN1725 : _GEN1703;
wire  _GEN1727 = io_x[15] ? _GEN1726 : _GEN1685;
wire  _GEN1728 = io_x[12] ? _GEN1727 : _GEN1656;
wire  _GEN1729 = io_x[10] ? _GEN1728 : _GEN1595;
wire  _GEN1730 = io_x[4] ? _GEN1729 : _GEN1508;
wire  _GEN1731 = io_x[8] ? _GEN1730 : _GEN1405;
wire  _GEN1732 = io_x[29] ? _GEN1731 : _GEN1167;
wire  _GEN1733 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1734 = io_x[7] ? _GEN1733 : _GEN241;
wire  _GEN1735 = io_x[2] ? _GEN233 : _GEN1734;
wire  _GEN1736 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1737 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1738 = io_x[11] ? _GEN1737 : _GEN1736;
wire  _GEN1739 = io_x[3] ? _GEN1738 : _GEN209;
wire  _GEN1740 = io_x[7] ? _GEN1739 : _GEN203;
wire  _GEN1741 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1742 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1743 = io_x[11] ? _GEN1742 : _GEN1741;
wire  _GEN1744 = io_x[3] ? _GEN1743 : _GEN209;
wire  _GEN1745 = io_x[7] ? _GEN1744 : _GEN203;
wire  _GEN1746 = io_x[2] ? _GEN1745 : _GEN1740;
wire  _GEN1747 = io_x[17] ? _GEN1746 : _GEN1735;
wire  _GEN1748 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1749 = io_x[11] ? _GEN1748 : _GEN214;
wire  _GEN1750 = io_x[3] ? _GEN1749 : _GEN216;
wire  _GEN1751 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1752 = io_x[3] ? _GEN1751 : _GEN216;
wire  _GEN1753 = io_x[7] ? _GEN1752 : _GEN1750;
wire  _GEN1754 = io_x[2] ? _GEN233 : _GEN1753;
wire  _GEN1755 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN1756 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1757 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1758 = io_x[11] ? _GEN1757 : _GEN1756;
wire  _GEN1759 = io_x[3] ? _GEN1758 : _GEN216;
wire  _GEN1760 = io_x[7] ? _GEN1759 : _GEN1755;
wire  _GEN1761 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1762 = io_x[11] ? _GEN1761 : _GEN214;
wire  _GEN1763 = io_x[3] ? _GEN1762 : _GEN216;
wire  _GEN1764 = io_x[7] ? _GEN1763 : _GEN241;
wire  _GEN1765 = io_x[2] ? _GEN1764 : _GEN1760;
wire  _GEN1766 = io_x[17] ? _GEN1765 : _GEN1754;
wire  _GEN1767 = io_x[15] ? _GEN1766 : _GEN1747;
wire  _GEN1768 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN1769 = io_x[2] ? _GEN233 : _GEN1768;
wire  _GEN1770 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1771 = io_x[3] ? _GEN1770 : _GEN216;
wire  _GEN1772 = io_x[7] ? _GEN241 : _GEN1771;
wire  _GEN1773 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1774 = io_x[11] ? _GEN1773 : _GEN214;
wire  _GEN1775 = io_x[3] ? _GEN1774 : _GEN209;
wire  _GEN1776 = io_x[7] ? _GEN241 : _GEN1775;
wire  _GEN1777 = io_x[2] ? _GEN1776 : _GEN1772;
wire  _GEN1778 = io_x[17] ? _GEN1777 : _GEN1769;
wire  _GEN1779 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1780 = io_x[3] ? _GEN1779 : _GEN216;
wire  _GEN1781 = io_x[7] ? _GEN203 : _GEN1780;
wire  _GEN1782 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1783 = io_x[3] ? _GEN1782 : _GEN216;
wire  _GEN1784 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1785 = io_x[11] ? _GEN1784 : _GEN214;
wire  _GEN1786 = io_x[3] ? _GEN1785 : _GEN209;
wire  _GEN1787 = io_x[7] ? _GEN1786 : _GEN1783;
wire  _GEN1788 = io_x[2] ? _GEN1787 : _GEN1781;
wire  _GEN1789 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1790 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1791 = io_x[11] ? _GEN1790 : _GEN1789;
wire  _GEN1792 = io_x[3] ? _GEN1791 : _GEN209;
wire  _GEN1793 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1794 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1795 = io_x[11] ? _GEN1794 : _GEN1793;
wire  _GEN1796 = io_x[3] ? _GEN1795 : _GEN216;
wire  _GEN1797 = io_x[7] ? _GEN1796 : _GEN1792;
wire  _GEN1798 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1799 = io_x[11] ? _GEN1798 : _GEN207;
wire  _GEN1800 = io_x[3] ? _GEN1799 : _GEN216;
wire  _GEN1801 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1802 = io_x[11] ? _GEN1801 : _GEN214;
wire  _GEN1803 = io_x[3] ? _GEN1802 : _GEN216;
wire  _GEN1804 = io_x[7] ? _GEN1803 : _GEN1800;
wire  _GEN1805 = io_x[2] ? _GEN1804 : _GEN1797;
wire  _GEN1806 = io_x[17] ? _GEN1805 : _GEN1788;
wire  _GEN1807 = io_x[15] ? _GEN1806 : _GEN1778;
wire  _GEN1808 = io_x[12] ? _GEN1807 : _GEN1767;
wire  _GEN1809 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1810 = io_x[11] ? _GEN1809 : _GEN214;
wire  _GEN1811 = io_x[3] ? _GEN1810 : _GEN216;
wire  _GEN1812 = io_x[7] ? _GEN1811 : _GEN203;
wire  _GEN1813 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN1814 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN1815 = io_x[7] ? _GEN1814 : _GEN1813;
wire  _GEN1816 = io_x[2] ? _GEN1815 : _GEN1812;
wire  _GEN1817 = io_x[17] ? _GEN1816 : _GEN1283;
wire  _GEN1818 = io_x[2] ? _GEN202 : _GEN233;
wire  _GEN1819 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1820 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1821 = io_x[11] ? _GEN1820 : _GEN207;
wire  _GEN1822 = io_x[3] ? _GEN1821 : _GEN1819;
wire  _GEN1823 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1824 = io_x[11] ? _GEN1823 : _GEN214;
wire  _GEN1825 = io_x[3] ? _GEN1824 : _GEN216;
wire  _GEN1826 = io_x[7] ? _GEN1825 : _GEN1822;
wire  _GEN1827 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1828 = io_x[11] ? _GEN1827 : _GEN207;
wire  _GEN1829 = io_x[3] ? _GEN1828 : _GEN216;
wire  _GEN1830 = io_x[7] ? _GEN1829 : _GEN241;
wire  _GEN1831 = io_x[2] ? _GEN1830 : _GEN1826;
wire  _GEN1832 = io_x[17] ? _GEN1831 : _GEN1818;
wire  _GEN1833 = io_x[15] ? _GEN1832 : _GEN1817;
wire  _GEN1834 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1835 = io_x[11] ? _GEN214 : _GEN1834;
wire  _GEN1836 = io_x[3] ? _GEN1835 : _GEN209;
wire  _GEN1837 = io_x[7] ? _GEN203 : _GEN1836;
wire  _GEN1838 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1839 = io_x[3] ? _GEN1838 : _GEN216;
wire  _GEN1840 = io_x[7] ? _GEN1839 : _GEN241;
wire  _GEN1841 = io_x[2] ? _GEN1840 : _GEN1837;
wire  _GEN1842 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN1843 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1844 = io_x[11] ? _GEN214 : _GEN1843;
wire  _GEN1845 = io_x[3] ? _GEN1844 : _GEN216;
wire  _GEN1846 = io_x[7] ? _GEN1845 : _GEN1842;
wire  _GEN1847 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1848 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1849 = io_x[11] ? _GEN1848 : _GEN1847;
wire  _GEN1850 = io_x[3] ? _GEN1849 : _GEN209;
wire  _GEN1851 = io_x[7] ? _GEN1850 : _GEN203;
wire  _GEN1852 = io_x[2] ? _GEN1851 : _GEN1846;
wire  _GEN1853 = io_x[17] ? _GEN1852 : _GEN1841;
wire  _GEN1854 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN1855 = io_x[2] ? _GEN202 : _GEN1854;
wire  _GEN1856 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1857 = io_x[11] ? _GEN207 : _GEN1856;
wire  _GEN1858 = io_x[3] ? _GEN1857 : _GEN216;
wire  _GEN1859 = io_x[7] ? _GEN1858 : _GEN203;
wire  _GEN1860 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN1861 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1862 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1863 = io_x[11] ? _GEN1862 : _GEN207;
wire  _GEN1864 = io_x[3] ? _GEN1863 : _GEN1861;
wire  _GEN1865 = io_x[7] ? _GEN1864 : _GEN1860;
wire  _GEN1866 = io_x[2] ? _GEN1865 : _GEN1859;
wire  _GEN1867 = io_x[17] ? _GEN1866 : _GEN1855;
wire  _GEN1868 = io_x[15] ? _GEN1867 : _GEN1853;
wire  _GEN1869 = io_x[12] ? _GEN1868 : _GEN1833;
wire  _GEN1870 = io_x[10] ? _GEN1869 : _GEN1808;
wire  _GEN1871 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1872 = io_x[11] ? _GEN1871 : _GEN214;
wire  _GEN1873 = io_x[3] ? _GEN1872 : _GEN209;
wire  _GEN1874 = io_x[7] ? _GEN1873 : _GEN241;
wire  _GEN1875 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN1876 = io_x[7] ? _GEN1875 : _GEN203;
wire  _GEN1877 = io_x[2] ? _GEN1876 : _GEN1874;
wire  _GEN1878 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1879 = io_x[11] ? _GEN1878 : _GEN214;
wire  _GEN1880 = io_x[3] ? _GEN1879 : _GEN216;
wire  _GEN1881 = io_x[7] ? _GEN1880 : _GEN241;
wire  _GEN1882 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1883 = io_x[11] ? _GEN1882 : _GEN207;
wire  _GEN1884 = io_x[3] ? _GEN1883 : _GEN209;
wire  _GEN1885 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1886 = io_x[11] ? _GEN214 : _GEN1885;
wire  _GEN1887 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1888 = io_x[11] ? _GEN1887 : _GEN214;
wire  _GEN1889 = io_x[3] ? _GEN1888 : _GEN1886;
wire  _GEN1890 = io_x[7] ? _GEN1889 : _GEN1884;
wire  _GEN1891 = io_x[2] ? _GEN1890 : _GEN1881;
wire  _GEN1892 = io_x[17] ? _GEN1891 : _GEN1877;
wire  _GEN1893 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1894 = io_x[11] ? _GEN1893 : _GEN214;
wire  _GEN1895 = io_x[3] ? _GEN1894 : _GEN209;
wire  _GEN1896 = io_x[7] ? _GEN1895 : _GEN203;
wire  _GEN1897 = io_x[2] ? _GEN202 : _GEN1896;
wire  _GEN1898 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN1899 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1900 = io_x[11] ? _GEN1899 : _GEN214;
wire  _GEN1901 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1902 = io_x[11] ? _GEN1901 : _GEN214;
wire  _GEN1903 = io_x[3] ? _GEN1902 : _GEN1900;
wire  _GEN1904 = io_x[7] ? _GEN1903 : _GEN1898;
wire  _GEN1905 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1906 = io_x[11] ? _GEN214 : _GEN1905;
wire  _GEN1907 = io_x[3] ? _GEN1906 : _GEN209;
wire  _GEN1908 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1909 = io_x[11] ? _GEN1908 : _GEN214;
wire  _GEN1910 = io_x[3] ? _GEN1909 : _GEN209;
wire  _GEN1911 = io_x[7] ? _GEN1910 : _GEN1907;
wire  _GEN1912 = io_x[2] ? _GEN1911 : _GEN1904;
wire  _GEN1913 = io_x[17] ? _GEN1912 : _GEN1897;
wire  _GEN1914 = io_x[15] ? _GEN1913 : _GEN1892;
wire  _GEN1915 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN1916 = io_x[2] ? _GEN1915 : _GEN202;
wire  _GEN1917 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1918 = io_x[3] ? _GEN1917 : _GEN216;
wire  _GEN1919 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN1920 = io_x[7] ? _GEN1919 : _GEN1918;
wire  _GEN1921 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1922 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1923 = io_x[11] ? _GEN1922 : _GEN1921;
wire  _GEN1924 = io_x[3] ? _GEN1923 : _GEN216;
wire  _GEN1925 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1926 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1927 = io_x[11] ? _GEN1926 : _GEN1925;
wire  _GEN1928 = io_x[3] ? _GEN1927 : _GEN216;
wire  _GEN1929 = io_x[7] ? _GEN1928 : _GEN1924;
wire  _GEN1930 = io_x[2] ? _GEN1929 : _GEN1920;
wire  _GEN1931 = io_x[17] ? _GEN1930 : _GEN1916;
wire  _GEN1932 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1933 = io_x[3] ? _GEN209 : _GEN1932;
wire  _GEN1934 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1935 = io_x[11] ? _GEN1934 : _GEN214;
wire  _GEN1936 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1937 = io_x[3] ? _GEN1936 : _GEN1935;
wire  _GEN1938 = io_x[7] ? _GEN1937 : _GEN1933;
wire  _GEN1939 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1940 = io_x[11] ? _GEN1939 : _GEN214;
wire  _GEN1941 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1942 = io_x[11] ? _GEN214 : _GEN1941;
wire  _GEN1943 = io_x[3] ? _GEN1942 : _GEN1940;
wire  _GEN1944 = io_x[7] ? _GEN1943 : _GEN241;
wire  _GEN1945 = io_x[2] ? _GEN1944 : _GEN1938;
wire  _GEN1946 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1947 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1948 = io_x[11] ? _GEN214 : _GEN1947;
wire  _GEN1949 = io_x[3] ? _GEN1948 : _GEN1946;
wire  _GEN1950 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1951 = io_x[11] ? _GEN1950 : _GEN214;
wire  _GEN1952 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1953 = io_x[11] ? _GEN1952 : _GEN214;
wire  _GEN1954 = io_x[3] ? _GEN1953 : _GEN1951;
wire  _GEN1955 = io_x[7] ? _GEN1954 : _GEN1949;
wire  _GEN1956 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1957 = io_x[3] ? _GEN1956 : _GEN209;
wire  _GEN1958 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1959 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1960 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1961 = io_x[11] ? _GEN1960 : _GEN1959;
wire  _GEN1962 = io_x[3] ? _GEN1961 : _GEN1958;
wire  _GEN1963 = io_x[7] ? _GEN1962 : _GEN1957;
wire  _GEN1964 = io_x[2] ? _GEN1963 : _GEN1955;
wire  _GEN1965 = io_x[17] ? _GEN1964 : _GEN1945;
wire  _GEN1966 = io_x[15] ? _GEN1965 : _GEN1931;
wire  _GEN1967 = io_x[12] ? _GEN1966 : _GEN1914;
wire  _GEN1968 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1969 = io_x[11] ? _GEN1968 : _GEN207;
wire  _GEN1970 = io_x[3] ? _GEN216 : _GEN1969;
wire  _GEN1971 = io_x[7] ? _GEN1970 : _GEN241;
wire  _GEN1972 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1973 = io_x[11] ? _GEN207 : _GEN1972;
wire  _GEN1974 = io_x[3] ? _GEN1973 : _GEN209;
wire  _GEN1975 = io_x[7] ? _GEN1974 : _GEN203;
wire  _GEN1976 = io_x[2] ? _GEN1975 : _GEN1971;
wire  _GEN1977 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN1978 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1979 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1980 = io_x[11] ? _GEN1979 : _GEN1978;
wire  _GEN1981 = io_x[3] ? _GEN1980 : _GEN1977;
wire  _GEN1982 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN1983 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1984 = io_x[11] ? _GEN1983 : _GEN1982;
wire  _GEN1985 = io_x[3] ? _GEN216 : _GEN1984;
wire  _GEN1986 = io_x[7] ? _GEN1985 : _GEN1981;
wire  _GEN1987 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1988 = io_x[3] ? _GEN1987 : _GEN216;
wire  _GEN1989 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1990 = io_x[3] ? _GEN1989 : _GEN209;
wire  _GEN1991 = io_x[7] ? _GEN1990 : _GEN1988;
wire  _GEN1992 = io_x[2] ? _GEN1991 : _GEN1986;
wire  _GEN1993 = io_x[17] ? _GEN1992 : _GEN1976;
wire  _GEN1994 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN1995 = io_x[3] ? _GEN216 : _GEN1994;
wire  _GEN1996 = io_x[7] ? _GEN203 : _GEN1995;
wire  _GEN1997 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN1998 = io_x[11] ? _GEN1997 : _GEN214;
wire  _GEN1999 = io_x[3] ? _GEN216 : _GEN1998;
wire  _GEN2000 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2001 = io_x[11] ? _GEN2000 : _GEN214;
wire  _GEN2002 = io_x[3] ? _GEN2001 : _GEN216;
wire  _GEN2003 = io_x[7] ? _GEN2002 : _GEN1999;
wire  _GEN2004 = io_x[2] ? _GEN2003 : _GEN1996;
wire  _GEN2005 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2006 = io_x[3] ? _GEN216 : _GEN2005;
wire  _GEN2007 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2008 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2009 = io_x[11] ? _GEN2008 : _GEN2007;
wire  _GEN2010 = io_x[3] ? _GEN2009 : _GEN216;
wire  _GEN2011 = io_x[7] ? _GEN2010 : _GEN2006;
wire  _GEN2012 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2013 = io_x[11] ? _GEN2012 : _GEN214;
wire  _GEN2014 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2015 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2016 = io_x[11] ? _GEN2015 : _GEN2014;
wire  _GEN2017 = io_x[3] ? _GEN2016 : _GEN2013;
wire  _GEN2018 = io_x[7] ? _GEN2017 : _GEN203;
wire  _GEN2019 = io_x[2] ? _GEN2018 : _GEN2011;
wire  _GEN2020 = io_x[17] ? _GEN2019 : _GEN2004;
wire  _GEN2021 = io_x[15] ? _GEN2020 : _GEN1993;
wire  _GEN2022 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2023 = io_x[11] ? _GEN214 : _GEN2022;
wire  _GEN2024 = io_x[3] ? _GEN2023 : _GEN209;
wire  _GEN2025 = io_x[7] ? _GEN2024 : _GEN203;
wire  _GEN2026 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2027 = io_x[11] ? _GEN214 : _GEN2026;
wire  _GEN2028 = io_x[3] ? _GEN216 : _GEN2027;
wire  _GEN2029 = io_x[7] ? _GEN241 : _GEN2028;
wire  _GEN2030 = io_x[2] ? _GEN2029 : _GEN2025;
wire  _GEN2031 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2032 = io_x[3] ? _GEN2031 : _GEN216;
wire  _GEN2033 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2034 = io_x[11] ? _GEN2033 : _GEN207;
wire  _GEN2035 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2036 = io_x[11] ? _GEN214 : _GEN2035;
wire  _GEN2037 = io_x[3] ? _GEN2036 : _GEN2034;
wire  _GEN2038 = io_x[7] ? _GEN2037 : _GEN2032;
wire  _GEN2039 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2040 = io_x[11] ? _GEN214 : _GEN2039;
wire  _GEN2041 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2042 = io_x[11] ? _GEN214 : _GEN2041;
wire  _GEN2043 = io_x[3] ? _GEN2042 : _GEN2040;
wire  _GEN2044 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2045 = io_x[11] ? _GEN2044 : _GEN207;
wire  _GEN2046 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2047 = io_x[11] ? _GEN214 : _GEN2046;
wire  _GEN2048 = io_x[3] ? _GEN2047 : _GEN2045;
wire  _GEN2049 = io_x[7] ? _GEN2048 : _GEN2043;
wire  _GEN2050 = io_x[2] ? _GEN2049 : _GEN2038;
wire  _GEN2051 = io_x[17] ? _GEN2050 : _GEN2030;
wire  _GEN2052 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2053 = io_x[11] ? _GEN2052 : _GEN214;
wire  _GEN2054 = io_x[3] ? _GEN2053 : _GEN209;
wire  _GEN2055 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2056 = io_x[7] ? _GEN2055 : _GEN2054;
wire  _GEN2057 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2058 = io_x[11] ? _GEN2057 : _GEN214;
wire  _GEN2059 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2060 = io_x[11] ? _GEN2059 : _GEN214;
wire  _GEN2061 = io_x[3] ? _GEN2060 : _GEN2058;
wire  _GEN2062 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2063 = io_x[11] ? _GEN2062 : _GEN214;
wire  _GEN2064 = io_x[3] ? _GEN2063 : _GEN216;
wire  _GEN2065 = io_x[7] ? _GEN2064 : _GEN2061;
wire  _GEN2066 = io_x[2] ? _GEN2065 : _GEN2056;
wire  _GEN2067 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2068 = io_x[11] ? _GEN2067 : _GEN214;
wire  _GEN2069 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2070 = io_x[11] ? _GEN207 : _GEN2069;
wire  _GEN2071 = io_x[3] ? _GEN2070 : _GEN2068;
wire  _GEN2072 = io_x[7] ? _GEN2071 : _GEN241;
wire  _GEN2073 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2074 = io_x[11] ? _GEN2073 : _GEN214;
wire  _GEN2075 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2076 = io_x[11] ? _GEN2075 : _GEN207;
wire  _GEN2077 = io_x[3] ? _GEN2076 : _GEN2074;
wire  _GEN2078 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2079 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2080 = io_x[11] ? _GEN2079 : _GEN2078;
wire  _GEN2081 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2082 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2083 = io_x[11] ? _GEN2082 : _GEN2081;
wire  _GEN2084 = io_x[3] ? _GEN2083 : _GEN2080;
wire  _GEN2085 = io_x[7] ? _GEN2084 : _GEN2077;
wire  _GEN2086 = io_x[2] ? _GEN2085 : _GEN2072;
wire  _GEN2087 = io_x[17] ? _GEN2086 : _GEN2066;
wire  _GEN2088 = io_x[15] ? _GEN2087 : _GEN2051;
wire  _GEN2089 = io_x[12] ? _GEN2088 : _GEN2021;
wire  _GEN2090 = io_x[10] ? _GEN2089 : _GEN1967;
wire  _GEN2091 = io_x[4] ? _GEN2090 : _GEN1870;
wire  _GEN2092 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN2093 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2094 = io_x[11] ? _GEN2093 : _GEN214;
wire  _GEN2095 = io_x[3] ? _GEN2094 : _GEN216;
wire  _GEN2096 = io_x[7] ? _GEN2095 : _GEN241;
wire  _GEN2097 = io_x[2] ? _GEN2096 : _GEN2092;
wire  _GEN2098 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2099 = io_x[11] ? _GEN2098 : _GEN214;
wire  _GEN2100 = io_x[3] ? _GEN2099 : _GEN216;
wire  _GEN2101 = io_x[7] ? _GEN2100 : _GEN203;
wire  _GEN2102 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2103 = io_x[3] ? _GEN2102 : _GEN209;
wire  _GEN2104 = io_x[7] ? _GEN203 : _GEN2103;
wire  _GEN2105 = io_x[2] ? _GEN2104 : _GEN2101;
wire  _GEN2106 = io_x[17] ? _GEN2105 : _GEN2097;
wire  _GEN2107 = io_x[7] ? _GEN203 : _GEN241;
wire  _GEN2108 = io_x[7] ? _GEN203 : _GEN241;
wire  _GEN2109 = io_x[2] ? _GEN2108 : _GEN2107;
wire  _GEN2110 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2111 = io_x[11] ? _GEN2110 : _GEN214;
wire  _GEN2112 = io_x[3] ? _GEN2111 : _GEN209;
wire  _GEN2113 = io_x[7] ? _GEN2112 : _GEN241;
wire  _GEN2114 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2115 = io_x[11] ? _GEN2114 : _GEN214;
wire  _GEN2116 = io_x[3] ? _GEN216 : _GEN2115;
wire  _GEN2117 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2118 = io_x[11] ? _GEN2117 : _GEN214;
wire  _GEN2119 = io_x[3] ? _GEN2118 : _GEN209;
wire  _GEN2120 = io_x[7] ? _GEN2119 : _GEN2116;
wire  _GEN2121 = io_x[2] ? _GEN2120 : _GEN2113;
wire  _GEN2122 = io_x[17] ? _GEN2121 : _GEN2109;
wire  _GEN2123 = io_x[15] ? _GEN2122 : _GEN2106;
wire  _GEN2124 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2125 = io_x[3] ? _GEN216 : _GEN2124;
wire  _GEN2126 = io_x[7] ? _GEN241 : _GEN2125;
wire  _GEN2127 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2128 = io_x[3] ? _GEN2127 : _GEN216;
wire  _GEN2129 = io_x[7] ? _GEN2128 : _GEN203;
wire  _GEN2130 = io_x[2] ? _GEN2129 : _GEN2126;
wire  _GEN2131 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2132 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2133 = io_x[11] ? _GEN2132 : _GEN214;
wire  _GEN2134 = io_x[3] ? _GEN2133 : _GEN2131;
wire  _GEN2135 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2136 = io_x[11] ? _GEN2135 : _GEN214;
wire  _GEN2137 = io_x[3] ? _GEN2136 : _GEN216;
wire  _GEN2138 = io_x[7] ? _GEN2137 : _GEN2134;
wire  _GEN2139 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2140 = io_x[11] ? _GEN2139 : _GEN214;
wire  _GEN2141 = io_x[3] ? _GEN2140 : _GEN209;
wire  _GEN2142 = io_x[7] ? _GEN2141 : _GEN203;
wire  _GEN2143 = io_x[2] ? _GEN2142 : _GEN2138;
wire  _GEN2144 = io_x[17] ? _GEN2143 : _GEN2130;
wire  _GEN2145 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN2146 = io_x[2] ? _GEN2145 : _GEN202;
wire  _GEN2147 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2148 = io_x[11] ? _GEN214 : _GEN2147;
wire  _GEN2149 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2150 = io_x[11] ? _GEN2149 : _GEN214;
wire  _GEN2151 = io_x[3] ? _GEN2150 : _GEN2148;
wire  _GEN2152 = io_x[7] ? _GEN2151 : _GEN203;
wire  _GEN2153 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2154 = io_x[11] ? _GEN207 : _GEN2153;
wire  _GEN2155 = io_x[3] ? _GEN216 : _GEN2154;
wire  _GEN2156 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2157 = io_x[11] ? _GEN207 : _GEN2156;
wire  _GEN2158 = io_x[3] ? _GEN2157 : _GEN209;
wire  _GEN2159 = io_x[7] ? _GEN2158 : _GEN2155;
wire  _GEN2160 = io_x[2] ? _GEN2159 : _GEN2152;
wire  _GEN2161 = io_x[17] ? _GEN2160 : _GEN2146;
wire  _GEN2162 = io_x[15] ? _GEN2161 : _GEN2144;
wire  _GEN2163 = io_x[12] ? _GEN2162 : _GEN2123;
wire  _GEN2164 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2165 = io_x[3] ? _GEN216 : _GEN2164;
wire  _GEN2166 = io_x[7] ? _GEN203 : _GEN2165;
wire  _GEN2167 = io_x[2] ? _GEN2166 : _GEN233;
wire  _GEN2168 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2169 = io_x[11] ? _GEN2168 : _GEN214;
wire  _GEN2170 = io_x[3] ? _GEN2169 : _GEN216;
wire  _GEN2171 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2172 = io_x[11] ? _GEN214 : _GEN2171;
wire  _GEN2173 = io_x[3] ? _GEN2172 : _GEN216;
wire  _GEN2174 = io_x[7] ? _GEN2173 : _GEN2170;
wire  _GEN2175 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2176 = io_x[11] ? _GEN214 : _GEN2175;
wire  _GEN2177 = io_x[3] ? _GEN2176 : _GEN209;
wire  _GEN2178 = io_x[7] ? _GEN203 : _GEN2177;
wire  _GEN2179 = io_x[2] ? _GEN2178 : _GEN2174;
wire  _GEN2180 = io_x[17] ? _GEN2179 : _GEN2167;
wire  _GEN2181 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2182 = io_x[11] ? _GEN2181 : _GEN214;
wire  _GEN2183 = io_x[3] ? _GEN2182 : _GEN209;
wire  _GEN2184 = io_x[7] ? _GEN241 : _GEN2183;
wire  _GEN2185 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2186 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2187 = io_x[11] ? _GEN2186 : _GEN2185;
wire  _GEN2188 = io_x[3] ? _GEN2187 : _GEN216;
wire  _GEN2189 = io_x[7] ? _GEN2188 : _GEN203;
wire  _GEN2190 = io_x[2] ? _GEN2189 : _GEN2184;
wire  _GEN2191 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2192 = io_x[11] ? _GEN2191 : _GEN214;
wire  _GEN2193 = io_x[3] ? _GEN2192 : _GEN216;
wire  _GEN2194 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2195 = io_x[11] ? _GEN207 : _GEN2194;
wire  _GEN2196 = io_x[3] ? _GEN2195 : _GEN209;
wire  _GEN2197 = io_x[7] ? _GEN2196 : _GEN2193;
wire  _GEN2198 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2199 = io_x[11] ? _GEN207 : _GEN2198;
wire  _GEN2200 = io_x[3] ? _GEN209 : _GEN2199;
wire  _GEN2201 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2202 = io_x[11] ? _GEN2201 : _GEN207;
wire  _GEN2203 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2204 = io_x[11] ? _GEN2203 : _GEN214;
wire  _GEN2205 = io_x[3] ? _GEN2204 : _GEN2202;
wire  _GEN2206 = io_x[7] ? _GEN2205 : _GEN2200;
wire  _GEN2207 = io_x[2] ? _GEN2206 : _GEN2197;
wire  _GEN2208 = io_x[17] ? _GEN2207 : _GEN2190;
wire  _GEN2209 = io_x[15] ? _GEN2208 : _GEN2180;
wire  _GEN2210 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2211 = io_x[11] ? _GEN2210 : _GEN214;
wire  _GEN2212 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2213 = io_x[11] ? _GEN214 : _GEN2212;
wire  _GEN2214 = io_x[3] ? _GEN2213 : _GEN2211;
wire  _GEN2215 = io_x[7] ? _GEN2214 : _GEN241;
wire  _GEN2216 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2217 = io_x[3] ? _GEN2216 : _GEN216;
wire  _GEN2218 = io_x[7] ? _GEN203 : _GEN2217;
wire  _GEN2219 = io_x[2] ? _GEN2218 : _GEN2215;
wire  _GEN2220 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2221 = io_x[11] ? _GEN214 : _GEN2220;
wire  _GEN2222 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2223 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2224 = io_x[11] ? _GEN2223 : _GEN2222;
wire  _GEN2225 = io_x[3] ? _GEN2224 : _GEN2221;
wire  _GEN2226 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2227 = io_x[11] ? _GEN2226 : _GEN214;
wire  _GEN2228 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2229 = io_x[11] ? _GEN214 : _GEN2228;
wire  _GEN2230 = io_x[3] ? _GEN2229 : _GEN2227;
wire  _GEN2231 = io_x[7] ? _GEN2230 : _GEN2225;
wire  _GEN2232 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2233 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2234 = io_x[3] ? _GEN2233 : _GEN2232;
wire  _GEN2235 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2236 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2237 = io_x[11] ? _GEN2236 : _GEN207;
wire  _GEN2238 = io_x[3] ? _GEN2237 : _GEN2235;
wire  _GEN2239 = io_x[7] ? _GEN2238 : _GEN2234;
wire  _GEN2240 = io_x[2] ? _GEN2239 : _GEN2231;
wire  _GEN2241 = io_x[17] ? _GEN2240 : _GEN2219;
wire  _GEN2242 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2243 = io_x[7] ? _GEN2242 : _GEN203;
wire  _GEN2244 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2245 = io_x[11] ? _GEN2244 : _GEN207;
wire  _GEN2246 = io_x[3] ? _GEN2245 : _GEN216;
wire  _GEN2247 = io_x[7] ? _GEN2246 : _GEN203;
wire  _GEN2248 = io_x[2] ? _GEN2247 : _GEN2243;
wire  _GEN2249 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2250 = io_x[11] ? _GEN214 : _GEN2249;
wire  _GEN2251 = io_x[3] ? _GEN2250 : _GEN209;
wire  _GEN2252 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2253 = io_x[11] ? _GEN2252 : _GEN214;
wire  _GEN2254 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2255 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2256 = io_x[11] ? _GEN2255 : _GEN2254;
wire  _GEN2257 = io_x[3] ? _GEN2256 : _GEN2253;
wire  _GEN2258 = io_x[7] ? _GEN2257 : _GEN2251;
wire  _GEN2259 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2260 = io_x[11] ? _GEN207 : _GEN2259;
wire  _GEN2261 = io_x[3] ? _GEN216 : _GEN2260;
wire  _GEN2262 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2263 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2264 = io_x[11] ? _GEN2263 : _GEN2262;
wire  _GEN2265 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2266 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2267 = io_x[11] ? _GEN2266 : _GEN2265;
wire  _GEN2268 = io_x[3] ? _GEN2267 : _GEN2264;
wire  _GEN2269 = io_x[7] ? _GEN2268 : _GEN2261;
wire  _GEN2270 = io_x[2] ? _GEN2269 : _GEN2258;
wire  _GEN2271 = io_x[17] ? _GEN2270 : _GEN2248;
wire  _GEN2272 = io_x[15] ? _GEN2271 : _GEN2241;
wire  _GEN2273 = io_x[12] ? _GEN2272 : _GEN2209;
wire  _GEN2274 = io_x[10] ? _GEN2273 : _GEN2163;
wire  _GEN2275 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2276 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2277 = io_x[11] ? _GEN2276 : _GEN214;
wire  _GEN2278 = io_x[3] ? _GEN2277 : _GEN2275;
wire  _GEN2279 = io_x[7] ? _GEN203 : _GEN2278;
wire  _GEN2280 = io_x[2] ? _GEN2279 : _GEN202;
wire  _GEN2281 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2282 = io_x[11] ? _GEN2281 : _GEN207;
wire  _GEN2283 = io_x[3] ? _GEN2282 : _GEN209;
wire  _GEN2284 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2285 = io_x[11] ? _GEN2284 : _GEN207;
wire  _GEN2286 = io_x[3] ? _GEN2285 : _GEN209;
wire  _GEN2287 = io_x[7] ? _GEN2286 : _GEN2283;
wire  _GEN2288 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2289 = io_x[11] ? _GEN2288 : _GEN214;
wire  _GEN2290 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2291 = io_x[11] ? _GEN2290 : _GEN207;
wire  _GEN2292 = io_x[3] ? _GEN2291 : _GEN2289;
wire  _GEN2293 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2294 = io_x[11] ? _GEN2293 : _GEN214;
wire  _GEN2295 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2296 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2297 = io_x[11] ? _GEN2296 : _GEN2295;
wire  _GEN2298 = io_x[3] ? _GEN2297 : _GEN2294;
wire  _GEN2299 = io_x[7] ? _GEN2298 : _GEN2292;
wire  _GEN2300 = io_x[2] ? _GEN2299 : _GEN2287;
wire  _GEN2301 = io_x[17] ? _GEN2300 : _GEN2280;
wire  _GEN2302 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2303 = io_x[3] ? _GEN216 : _GEN2302;
wire  _GEN2304 = io_x[7] ? _GEN2303 : _GEN203;
wire  _GEN2305 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2306 = io_x[3] ? _GEN209 : _GEN2305;
wire  _GEN2307 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2308 = io_x[11] ? _GEN2307 : _GEN214;
wire  _GEN2309 = io_x[3] ? _GEN2308 : _GEN209;
wire  _GEN2310 = io_x[7] ? _GEN2309 : _GEN2306;
wire  _GEN2311 = io_x[2] ? _GEN2310 : _GEN2304;
wire  _GEN2312 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2313 = io_x[11] ? _GEN2312 : _GEN214;
wire  _GEN2314 = io_x[3] ? _GEN2313 : _GEN216;
wire  _GEN2315 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2316 = io_x[11] ? _GEN2315 : _GEN207;
wire  _GEN2317 = io_x[3] ? _GEN2316 : _GEN216;
wire  _GEN2318 = io_x[7] ? _GEN2317 : _GEN2314;
wire  _GEN2319 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2320 = io_x[11] ? _GEN2319 : _GEN214;
wire  _GEN2321 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2322 = io_x[11] ? _GEN2321 : _GEN214;
wire  _GEN2323 = io_x[3] ? _GEN2322 : _GEN2320;
wire  _GEN2324 = io_x[7] ? _GEN241 : _GEN2323;
wire  _GEN2325 = io_x[2] ? _GEN2324 : _GEN2318;
wire  _GEN2326 = io_x[17] ? _GEN2325 : _GEN2311;
wire  _GEN2327 = io_x[15] ? _GEN2326 : _GEN2301;
wire  _GEN2328 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2329 = io_x[3] ? _GEN2328 : _GEN209;
wire  _GEN2330 = io_x[7] ? _GEN2329 : _GEN203;
wire  _GEN2331 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2332 = io_x[11] ? _GEN2331 : _GEN214;
wire  _GEN2333 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2334 = io_x[11] ? _GEN2333 : _GEN207;
wire  _GEN2335 = io_x[3] ? _GEN2334 : _GEN2332;
wire  _GEN2336 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2337 = io_x[11] ? _GEN2336 : _GEN214;
wire  _GEN2338 = io_x[3] ? _GEN2337 : _GEN216;
wire  _GEN2339 = io_x[7] ? _GEN2338 : _GEN2335;
wire  _GEN2340 = io_x[2] ? _GEN2339 : _GEN2330;
wire  _GEN2341 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2342 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2343 = io_x[11] ? _GEN2342 : _GEN2341;
wire  _GEN2344 = io_x[3] ? _GEN2343 : _GEN209;
wire  _GEN2345 = io_x[7] ? _GEN2344 : _GEN203;
wire  _GEN2346 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2347 = io_x[11] ? _GEN2346 : _GEN214;
wire  _GEN2348 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2349 = io_x[11] ? _GEN2348 : _GEN214;
wire  _GEN2350 = io_x[3] ? _GEN2349 : _GEN2347;
wire  _GEN2351 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2352 = io_x[11] ? _GEN214 : _GEN2351;
wire  _GEN2353 = io_x[3] ? _GEN2352 : _GEN209;
wire  _GEN2354 = io_x[7] ? _GEN2353 : _GEN2350;
wire  _GEN2355 = io_x[2] ? _GEN2354 : _GEN2345;
wire  _GEN2356 = io_x[17] ? _GEN2355 : _GEN2340;
wire  _GEN2357 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2358 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2359 = io_x[3] ? _GEN2358 : _GEN2357;
wire  _GEN2360 = io_x[7] ? _GEN2359 : _GEN203;
wire  _GEN2361 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2362 = io_x[11] ? _GEN207 : _GEN2361;
wire  _GEN2363 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2364 = io_x[11] ? _GEN2363 : _GEN214;
wire  _GEN2365 = io_x[3] ? _GEN2364 : _GEN2362;
wire  _GEN2366 = io_x[7] ? _GEN2365 : _GEN241;
wire  _GEN2367 = io_x[2] ? _GEN2366 : _GEN2360;
wire  _GEN2368 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2369 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2370 = io_x[11] ? _GEN2369 : _GEN2368;
wire  _GEN2371 = io_x[3] ? _GEN2370 : _GEN209;
wire  _GEN2372 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2373 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2374 = io_x[11] ? _GEN2373 : _GEN2372;
wire  _GEN2375 = io_x[3] ? _GEN2374 : _GEN216;
wire  _GEN2376 = io_x[7] ? _GEN2375 : _GEN2371;
wire  _GEN2377 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2378 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2379 = io_x[11] ? _GEN2378 : _GEN2377;
wire  _GEN2380 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2381 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2382 = io_x[11] ? _GEN2381 : _GEN2380;
wire  _GEN2383 = io_x[3] ? _GEN2382 : _GEN2379;
wire  _GEN2384 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2385 = io_x[11] ? _GEN2384 : _GEN214;
wire  _GEN2386 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2387 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2388 = io_x[11] ? _GEN2387 : _GEN2386;
wire  _GEN2389 = io_x[3] ? _GEN2388 : _GEN2385;
wire  _GEN2390 = io_x[7] ? _GEN2389 : _GEN2383;
wire  _GEN2391 = io_x[2] ? _GEN2390 : _GEN2376;
wire  _GEN2392 = io_x[17] ? _GEN2391 : _GEN2367;
wire  _GEN2393 = io_x[15] ? _GEN2392 : _GEN2356;
wire  _GEN2394 = io_x[12] ? _GEN2393 : _GEN2327;
wire  _GEN2395 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2396 = io_x[3] ? _GEN2395 : _GEN216;
wire  _GEN2397 = io_x[7] ? _GEN2396 : _GEN241;
wire  _GEN2398 = io_x[2] ? _GEN2397 : _GEN233;
wire  _GEN2399 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2400 = io_x[3] ? _GEN2399 : _GEN216;
wire  _GEN2401 = io_x[7] ? _GEN2400 : _GEN203;
wire  _GEN2402 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2403 = io_x[11] ? _GEN2402 : _GEN207;
wire  _GEN2404 = io_x[3] ? _GEN2403 : _GEN216;
wire  _GEN2405 = io_x[7] ? _GEN2404 : _GEN241;
wire  _GEN2406 = io_x[2] ? _GEN2405 : _GEN2401;
wire  _GEN2407 = io_x[17] ? _GEN2406 : _GEN2398;
wire  _GEN2408 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2409 = io_x[11] ? _GEN2408 : _GEN214;
wire  _GEN2410 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2411 = io_x[3] ? _GEN2410 : _GEN2409;
wire  _GEN2412 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2413 = io_x[11] ? _GEN2412 : _GEN214;
wire  _GEN2414 = io_x[3] ? _GEN2413 : _GEN216;
wire  _GEN2415 = io_x[7] ? _GEN2414 : _GEN2411;
wire  _GEN2416 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2417 = io_x[11] ? _GEN2416 : _GEN214;
wire  _GEN2418 = io_x[3] ? _GEN2417 : _GEN216;
wire  _GEN2419 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2420 = io_x[11] ? _GEN2419 : _GEN214;
wire  _GEN2421 = io_x[3] ? _GEN2420 : _GEN209;
wire  _GEN2422 = io_x[7] ? _GEN2421 : _GEN2418;
wire  _GEN2423 = io_x[2] ? _GEN2422 : _GEN2415;
wire  _GEN2424 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2425 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2426 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2427 = io_x[11] ? _GEN2426 : _GEN2425;
wire  _GEN2428 = io_x[3] ? _GEN2427 : _GEN2424;
wire  _GEN2429 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2430 = io_x[11] ? _GEN214 : _GEN2429;
wire  _GEN2431 = io_x[3] ? _GEN209 : _GEN2430;
wire  _GEN2432 = io_x[7] ? _GEN2431 : _GEN2428;
wire  _GEN2433 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2434 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2435 = io_x[11] ? _GEN2434 : _GEN2433;
wire  _GEN2436 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2437 = io_x[11] ? _GEN2436 : _GEN214;
wire  _GEN2438 = io_x[3] ? _GEN2437 : _GEN2435;
wire  _GEN2439 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2440 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2441 = io_x[11] ? _GEN2440 : _GEN2439;
wire  _GEN2442 = io_x[3] ? _GEN2441 : _GEN216;
wire  _GEN2443 = io_x[7] ? _GEN2442 : _GEN2438;
wire  _GEN2444 = io_x[2] ? _GEN2443 : _GEN2432;
wire  _GEN2445 = io_x[17] ? _GEN2444 : _GEN2423;
wire  _GEN2446 = io_x[15] ? _GEN2445 : _GEN2407;
wire  _GEN2447 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2448 = io_x[3] ? _GEN2447 : _GEN209;
wire  _GEN2449 = io_x[7] ? _GEN203 : _GEN2448;
wire  _GEN2450 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2451 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2452 = io_x[11] ? _GEN2451 : _GEN2450;
wire  _GEN2453 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2454 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2455 = io_x[11] ? _GEN2454 : _GEN2453;
wire  _GEN2456 = io_x[3] ? _GEN2455 : _GEN2452;
wire  _GEN2457 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2458 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2459 = io_x[11] ? _GEN2458 : _GEN214;
wire  _GEN2460 = io_x[3] ? _GEN2459 : _GEN2457;
wire  _GEN2461 = io_x[7] ? _GEN2460 : _GEN2456;
wire  _GEN2462 = io_x[2] ? _GEN2461 : _GEN2449;
wire  _GEN2463 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2464 = io_x[11] ? _GEN214 : _GEN2463;
wire  _GEN2465 = io_x[3] ? _GEN2464 : _GEN209;
wire  _GEN2466 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2467 = io_x[11] ? _GEN207 : _GEN2466;
wire  _GEN2468 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2469 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2470 = io_x[11] ? _GEN2469 : _GEN2468;
wire  _GEN2471 = io_x[3] ? _GEN2470 : _GEN2467;
wire  _GEN2472 = io_x[7] ? _GEN2471 : _GEN2465;
wire  _GEN2473 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2474 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2475 = io_x[11] ? _GEN2474 : _GEN2473;
wire  _GEN2476 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2477 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2478 = io_x[11] ? _GEN2477 : _GEN2476;
wire  _GEN2479 = io_x[3] ? _GEN2478 : _GEN2475;
wire  _GEN2480 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2481 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2482 = io_x[11] ? _GEN2481 : _GEN2480;
wire  _GEN2483 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2484 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2485 = io_x[11] ? _GEN2484 : _GEN2483;
wire  _GEN2486 = io_x[3] ? _GEN2485 : _GEN2482;
wire  _GEN2487 = io_x[7] ? _GEN2486 : _GEN2479;
wire  _GEN2488 = io_x[2] ? _GEN2487 : _GEN2472;
wire  _GEN2489 = io_x[17] ? _GEN2488 : _GEN2462;
wire  _GEN2490 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2491 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2492 = io_x[11] ? _GEN2491 : _GEN214;
wire  _GEN2493 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2494 = io_x[11] ? _GEN2493 : _GEN207;
wire  _GEN2495 = io_x[3] ? _GEN2494 : _GEN2492;
wire  _GEN2496 = io_x[7] ? _GEN2495 : _GEN2490;
wire  _GEN2497 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2498 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2499 = io_x[11] ? _GEN2498 : _GEN214;
wire  _GEN2500 = io_x[3] ? _GEN2499 : _GEN2497;
wire  _GEN2501 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2502 = io_x[11] ? _GEN2501 : _GEN214;
wire  _GEN2503 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2504 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2505 = io_x[11] ? _GEN2504 : _GEN2503;
wire  _GEN2506 = io_x[3] ? _GEN2505 : _GEN2502;
wire  _GEN2507 = io_x[7] ? _GEN2506 : _GEN2500;
wire  _GEN2508 = io_x[2] ? _GEN2507 : _GEN2496;
wire  _GEN2509 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2510 = io_x[11] ? _GEN2509 : _GEN214;
wire  _GEN2511 = io_x[3] ? _GEN2510 : _GEN216;
wire  _GEN2512 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2513 = io_x[11] ? _GEN2512 : _GEN207;
wire  _GEN2514 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2515 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2516 = io_x[11] ? _GEN2515 : _GEN2514;
wire  _GEN2517 = io_x[3] ? _GEN2516 : _GEN2513;
wire  _GEN2518 = io_x[7] ? _GEN2517 : _GEN2511;
wire  _GEN2519 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2520 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2521 = io_x[11] ? _GEN2520 : _GEN2519;
wire  _GEN2522 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2523 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2524 = io_x[11] ? _GEN2523 : _GEN2522;
wire  _GEN2525 = io_x[3] ? _GEN2524 : _GEN2521;
wire  _GEN2526 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2527 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2528 = io_x[11] ? _GEN2527 : _GEN2526;
wire  _GEN2529 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2530 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2531 = io_x[11] ? _GEN2530 : _GEN2529;
wire  _GEN2532 = io_x[3] ? _GEN2531 : _GEN2528;
wire  _GEN2533 = io_x[7] ? _GEN2532 : _GEN2525;
wire  _GEN2534 = io_x[2] ? _GEN2533 : _GEN2518;
wire  _GEN2535 = io_x[17] ? _GEN2534 : _GEN2508;
wire  _GEN2536 = io_x[15] ? _GEN2535 : _GEN2489;
wire  _GEN2537 = io_x[12] ? _GEN2536 : _GEN2446;
wire  _GEN2538 = io_x[10] ? _GEN2537 : _GEN2394;
wire  _GEN2539 = io_x[4] ? _GEN2538 : _GEN2274;
wire  _GEN2540 = io_x[8] ? _GEN2539 : _GEN2091;
wire  _GEN2541 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN2542 = io_x[2] ? _GEN233 : _GEN2541;
wire  _GEN2543 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2544 = io_x[11] ? _GEN2543 : _GEN214;
wire  _GEN2545 = io_x[3] ? _GEN2544 : _GEN209;
wire  _GEN2546 = io_x[7] ? _GEN2545 : _GEN203;
wire  _GEN2547 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2548 = io_x[3] ? _GEN209 : _GEN2547;
wire  _GEN2549 = io_x[7] ? _GEN2548 : _GEN203;
wire  _GEN2550 = io_x[2] ? _GEN2549 : _GEN2546;
wire  _GEN2551 = io_x[17] ? _GEN2550 : _GEN2542;
wire  _GEN2552 = io_x[7] ? _GEN203 : _GEN241;
wire  _GEN2553 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2554 = io_x[11] ? _GEN2553 : _GEN214;
wire  _GEN2555 = io_x[3] ? _GEN2554 : _GEN216;
wire  _GEN2556 = io_x[7] ? _GEN2555 : _GEN203;
wire  _GEN2557 = io_x[2] ? _GEN2556 : _GEN2552;
wire  _GEN2558 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2559 = io_x[11] ? _GEN2558 : _GEN214;
wire  _GEN2560 = io_x[3] ? _GEN2559 : _GEN216;
wire  _GEN2561 = io_x[7] ? _GEN2560 : _GEN203;
wire  _GEN2562 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2563 = io_x[11] ? _GEN2562 : _GEN214;
wire  _GEN2564 = io_x[3] ? _GEN2563 : _GEN216;
wire  _GEN2565 = io_x[7] ? _GEN2564 : _GEN203;
wire  _GEN2566 = io_x[2] ? _GEN2565 : _GEN2561;
wire  _GEN2567 = io_x[17] ? _GEN2566 : _GEN2557;
wire  _GEN2568 = io_x[15] ? _GEN2567 : _GEN2551;
wire  _GEN2569 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2570 = io_x[11] ? _GEN214 : _GEN2569;
wire  _GEN2571 = io_x[3] ? _GEN2570 : _GEN216;
wire  _GEN2572 = io_x[7] ? _GEN203 : _GEN2571;
wire  _GEN2573 = io_x[2] ? _GEN233 : _GEN2572;
wire  _GEN2574 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN2575 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2576 = io_x[11] ? _GEN2575 : _GEN214;
wire  _GEN2577 = io_x[3] ? _GEN2576 : _GEN209;
wire  _GEN2578 = io_x[7] ? _GEN2577 : _GEN2574;
wire  _GEN2579 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2580 = io_x[11] ? _GEN2579 : _GEN214;
wire  _GEN2581 = io_x[3] ? _GEN2580 : _GEN209;
wire  _GEN2582 = io_x[7] ? _GEN2581 : _GEN203;
wire  _GEN2583 = io_x[2] ? _GEN2582 : _GEN2578;
wire  _GEN2584 = io_x[17] ? _GEN2583 : _GEN2573;
wire  _GEN2585 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN2586 = io_x[2] ? _GEN2585 : _GEN202;
wire  _GEN2587 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2588 = io_x[3] ? _GEN209 : _GEN2587;
wire  _GEN2589 = io_x[7] ? _GEN2588 : _GEN241;
wire  _GEN2590 = io_x[2] ? _GEN2589 : _GEN202;
wire  _GEN2591 = io_x[17] ? _GEN2590 : _GEN2586;
wire  _GEN2592 = io_x[15] ? _GEN2591 : _GEN2584;
wire  _GEN2593 = io_x[12] ? _GEN2592 : _GEN2568;
wire  _GEN2594 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2595 = io_x[11] ? _GEN2594 : _GEN214;
wire  _GEN2596 = io_x[3] ? _GEN2595 : _GEN216;
wire  _GEN2597 = io_x[7] ? _GEN203 : _GEN2596;
wire  _GEN2598 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2599 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN2600 = io_x[7] ? _GEN2599 : _GEN2598;
wire  _GEN2601 = io_x[2] ? _GEN2600 : _GEN2597;
wire  _GEN2602 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2603 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2604 = io_x[3] ? _GEN2603 : _GEN216;
wire  _GEN2605 = io_x[7] ? _GEN2604 : _GEN2602;
wire  _GEN2606 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2607 = io_x[3] ? _GEN209 : _GEN2606;
wire  _GEN2608 = io_x[7] ? _GEN241 : _GEN2607;
wire  _GEN2609 = io_x[2] ? _GEN2608 : _GEN2605;
wire  _GEN2610 = io_x[17] ? _GEN2609 : _GEN2601;
wire  _GEN2611 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN2612 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2613 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2614 = io_x[11] ? _GEN2613 : _GEN207;
wire  _GEN2615 = io_x[3] ? _GEN2614 : _GEN2612;
wire  _GEN2616 = io_x[7] ? _GEN2615 : _GEN2611;
wire  _GEN2617 = io_x[2] ? _GEN2616 : _GEN233;
wire  _GEN2618 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2619 = io_x[3] ? _GEN216 : _GEN2618;
wire  _GEN2620 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2621 = io_x[3] ? _GEN2620 : _GEN209;
wire  _GEN2622 = io_x[7] ? _GEN2621 : _GEN2619;
wire  _GEN2623 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2624 = io_x[3] ? _GEN2623 : _GEN216;
wire  _GEN2625 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2626 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2627 = io_x[3] ? _GEN2626 : _GEN2625;
wire  _GEN2628 = io_x[7] ? _GEN2627 : _GEN2624;
wire  _GEN2629 = io_x[2] ? _GEN2628 : _GEN2622;
wire  _GEN2630 = io_x[17] ? _GEN2629 : _GEN2617;
wire  _GEN2631 = io_x[15] ? _GEN2630 : _GEN2610;
wire  _GEN2632 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2633 = io_x[11] ? _GEN214 : _GEN2632;
wire  _GEN2634 = io_x[3] ? _GEN2633 : _GEN216;
wire  _GEN2635 = io_x[7] ? _GEN2634 : _GEN241;
wire  _GEN2636 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2637 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2638 = io_x[11] ? _GEN214 : _GEN2637;
wire  _GEN2639 = io_x[3] ? _GEN2638 : _GEN2636;
wire  _GEN2640 = io_x[7] ? _GEN2639 : _GEN241;
wire  _GEN2641 = io_x[2] ? _GEN2640 : _GEN2635;
wire  _GEN2642 = io_x[17] ? _GEN2641 : _GEN1283;
wire  _GEN2643 = io_x[7] ? _GEN203 : _GEN241;
wire  _GEN2644 = io_x[2] ? _GEN2643 : _GEN233;
wire  _GEN2645 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN2646 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2647 = io_x[3] ? _GEN2646 : _GEN216;
wire  _GEN2648 = io_x[7] ? _GEN2647 : _GEN2645;
wire  _GEN2649 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2650 = io_x[3] ? _GEN216 : _GEN2649;
wire  _GEN2651 = io_x[7] ? _GEN2650 : _GEN241;
wire  _GEN2652 = io_x[2] ? _GEN2651 : _GEN2648;
wire  _GEN2653 = io_x[17] ? _GEN2652 : _GEN2644;
wire  _GEN2654 = io_x[15] ? _GEN2653 : _GEN2642;
wire  _GEN2655 = io_x[12] ? _GEN2654 : _GEN2631;
wire  _GEN2656 = io_x[10] ? _GEN2655 : _GEN2593;
wire  _GEN2657 = 1'b1;
wire  _GEN2658 = io_x[7] ? _GEN203 : _GEN241;
wire  _GEN2659 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2660 = io_x[11] ? _GEN2659 : _GEN214;
wire  _GEN2661 = io_x[3] ? _GEN2660 : _GEN216;
wire  _GEN2662 = io_x[7] ? _GEN2661 : _GEN203;
wire  _GEN2663 = io_x[2] ? _GEN2662 : _GEN2658;
wire  _GEN2664 = io_x[17] ? _GEN2663 : _GEN2657;
wire  _GEN2665 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN2666 = io_x[7] ? _GEN2665 : _GEN241;
wire  _GEN2667 = io_x[2] ? _GEN2666 : _GEN202;
wire  _GEN2668 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2669 = io_x[11] ? _GEN2668 : _GEN214;
wire  _GEN2670 = io_x[3] ? _GEN2669 : _GEN216;
wire  _GEN2671 = io_x[7] ? _GEN2670 : _GEN203;
wire  _GEN2672 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2673 = io_x[11] ? _GEN2672 : _GEN214;
wire  _GEN2674 = io_x[3] ? _GEN2673 : _GEN209;
wire  _GEN2675 = io_x[7] ? _GEN2674 : _GEN203;
wire  _GEN2676 = io_x[2] ? _GEN2675 : _GEN2671;
wire  _GEN2677 = io_x[17] ? _GEN2676 : _GEN2667;
wire  _GEN2678 = io_x[15] ? _GEN2677 : _GEN2664;
wire  _GEN2679 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2680 = io_x[7] ? _GEN2679 : _GEN241;
wire  _GEN2681 = io_x[2] ? _GEN2680 : _GEN233;
wire  _GEN2682 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN2683 = io_x[7] ? _GEN203 : _GEN2682;
wire  _GEN2684 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2685 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2686 = io_x[3] ? _GEN2685 : _GEN2684;
wire  _GEN2687 = io_x[7] ? _GEN2686 : _GEN241;
wire  _GEN2688 = io_x[2] ? _GEN2687 : _GEN2683;
wire  _GEN2689 = io_x[17] ? _GEN2688 : _GEN2681;
wire  _GEN2690 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2691 = io_x[7] ? _GEN2690 : _GEN203;
wire  _GEN2692 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2693 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2694 = io_x[11] ? _GEN2693 : _GEN2692;
wire  _GEN2695 = io_x[3] ? _GEN2694 : _GEN209;
wire  _GEN2696 = io_x[7] ? _GEN2695 : _GEN203;
wire  _GEN2697 = io_x[2] ? _GEN2696 : _GEN2691;
wire  _GEN2698 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2699 = io_x[11] ? _GEN2698 : _GEN207;
wire  _GEN2700 = io_x[3] ? _GEN2699 : _GEN209;
wire  _GEN2701 = io_x[7] ? _GEN2700 : _GEN241;
wire  _GEN2702 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2703 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2704 = io_x[11] ? _GEN2703 : _GEN2702;
wire  _GEN2705 = io_x[3] ? _GEN2704 : _GEN209;
wire  _GEN2706 = io_x[7] ? _GEN2705 : _GEN203;
wire  _GEN2707 = io_x[2] ? _GEN2706 : _GEN2701;
wire  _GEN2708 = io_x[17] ? _GEN2707 : _GEN2697;
wire  _GEN2709 = io_x[15] ? _GEN2708 : _GEN2689;
wire  _GEN2710 = io_x[12] ? _GEN2709 : _GEN2678;
wire  _GEN2711 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2712 = io_x[3] ? _GEN216 : _GEN2711;
wire  _GEN2713 = io_x[7] ? _GEN2712 : _GEN203;
wire  _GEN2714 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2715 = io_x[3] ? _GEN209 : _GEN2714;
wire  _GEN2716 = io_x[7] ? _GEN2715 : _GEN203;
wire  _GEN2717 = io_x[2] ? _GEN2716 : _GEN2713;
wire  _GEN2718 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2719 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2720 = io_x[11] ? _GEN214 : _GEN2719;
wire  _GEN2721 = io_x[3] ? _GEN216 : _GEN2720;
wire  _GEN2722 = io_x[7] ? _GEN2721 : _GEN2718;
wire  _GEN2723 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2724 = io_x[3] ? _GEN2723 : _GEN216;
wire  _GEN2725 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2726 = io_x[11] ? _GEN207 : _GEN2725;
wire  _GEN2727 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2728 = io_x[3] ? _GEN2727 : _GEN2726;
wire  _GEN2729 = io_x[7] ? _GEN2728 : _GEN2724;
wire  _GEN2730 = io_x[2] ? _GEN2729 : _GEN2722;
wire  _GEN2731 = io_x[17] ? _GEN2730 : _GEN2717;
wire  _GEN2732 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2733 = io_x[7] ? _GEN2732 : _GEN203;
wire  _GEN2734 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2735 = io_x[3] ? _GEN216 : _GEN2734;
wire  _GEN2736 = io_x[7] ? _GEN2735 : _GEN241;
wire  _GEN2737 = io_x[2] ? _GEN2736 : _GEN2733;
wire  _GEN2738 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2739 = io_x[11] ? _GEN214 : _GEN2738;
wire  _GEN2740 = io_x[3] ? _GEN209 : _GEN2739;
wire  _GEN2741 = io_x[7] ? _GEN2740 : _GEN203;
wire  _GEN2742 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2743 = io_x[3] ? _GEN2742 : _GEN209;
wire  _GEN2744 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2745 = io_x[11] ? _GEN2744 : _GEN207;
wire  _GEN2746 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2747 = io_x[11] ? _GEN2746 : _GEN214;
wire  _GEN2748 = io_x[3] ? _GEN2747 : _GEN2745;
wire  _GEN2749 = io_x[7] ? _GEN2748 : _GEN2743;
wire  _GEN2750 = io_x[2] ? _GEN2749 : _GEN2741;
wire  _GEN2751 = io_x[17] ? _GEN2750 : _GEN2737;
wire  _GEN2752 = io_x[15] ? _GEN2751 : _GEN2731;
wire  _GEN2753 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2754 = io_x[11] ? _GEN214 : _GEN2753;
wire  _GEN2755 = io_x[3] ? _GEN216 : _GEN2754;
wire  _GEN2756 = io_x[7] ? _GEN241 : _GEN2755;
wire  _GEN2757 = io_x[2] ? _GEN2756 : _GEN202;
wire  _GEN2758 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2759 = io_x[3] ? _GEN2758 : _GEN216;
wire  _GEN2760 = io_x[7] ? _GEN241 : _GEN2759;
wire  _GEN2761 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2762 = io_x[3] ? _GEN2761 : _GEN216;
wire  _GEN2763 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2764 = io_x[11] ? _GEN2763 : _GEN207;
wire  _GEN2765 = io_x[3] ? _GEN2764 : _GEN209;
wire  _GEN2766 = io_x[7] ? _GEN2765 : _GEN2762;
wire  _GEN2767 = io_x[2] ? _GEN2766 : _GEN2760;
wire  _GEN2768 = io_x[17] ? _GEN2767 : _GEN2757;
wire  _GEN2769 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN2770 = io_x[7] ? _GEN2769 : _GEN203;
wire  _GEN2771 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2772 = io_x[3] ? _GEN2771 : _GEN216;
wire  _GEN2773 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2774 = io_x[7] ? _GEN2773 : _GEN2772;
wire  _GEN2775 = io_x[2] ? _GEN2774 : _GEN2770;
wire  _GEN2776 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2777 = io_x[11] ? _GEN2776 : _GEN214;
wire  _GEN2778 = io_x[3] ? _GEN216 : _GEN2777;
wire  _GEN2779 = io_x[7] ? _GEN2778 : _GEN203;
wire  _GEN2780 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2781 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2782 = io_x[11] ? _GEN2781 : _GEN2780;
wire  _GEN2783 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2784 = io_x[11] ? _GEN2783 : _GEN207;
wire  _GEN2785 = io_x[3] ? _GEN2784 : _GEN2782;
wire  _GEN2786 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2787 = io_x[11] ? _GEN2786 : _GEN214;
wire  _GEN2788 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2789 = io_x[11] ? _GEN2788 : _GEN207;
wire  _GEN2790 = io_x[3] ? _GEN2789 : _GEN2787;
wire  _GEN2791 = io_x[7] ? _GEN2790 : _GEN2785;
wire  _GEN2792 = io_x[2] ? _GEN2791 : _GEN2779;
wire  _GEN2793 = io_x[17] ? _GEN2792 : _GEN2775;
wire  _GEN2794 = io_x[15] ? _GEN2793 : _GEN2768;
wire  _GEN2795 = io_x[12] ? _GEN2794 : _GEN2752;
wire  _GEN2796 = io_x[10] ? _GEN2795 : _GEN2710;
wire  _GEN2797 = io_x[4] ? _GEN2796 : _GEN2656;
wire  _GEN2798 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2799 = io_x[11] ? _GEN2798 : _GEN214;
wire  _GEN2800 = io_x[3] ? _GEN209 : _GEN2799;
wire  _GEN2801 = io_x[7] ? _GEN241 : _GEN2800;
wire  _GEN2802 = io_x[2] ? _GEN2801 : _GEN233;
wire  _GEN2803 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2804 = io_x[3] ? _GEN2803 : _GEN209;
wire  _GEN2805 = io_x[7] ? _GEN2804 : _GEN241;
wire  _GEN2806 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2807 = io_x[11] ? _GEN2806 : _GEN214;
wire  _GEN2808 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2809 = io_x[11] ? _GEN2808 : _GEN214;
wire  _GEN2810 = io_x[3] ? _GEN2809 : _GEN2807;
wire  _GEN2811 = io_x[7] ? _GEN203 : _GEN2810;
wire  _GEN2812 = io_x[2] ? _GEN2811 : _GEN2805;
wire  _GEN2813 = io_x[17] ? _GEN2812 : _GEN2802;
wire  _GEN2814 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN2815 = io_x[7] ? _GEN203 : _GEN2814;
wire  _GEN2816 = io_x[2] ? _GEN2815 : _GEN202;
wire  _GEN2817 = io_x[7] ? _GEN241 : _GEN203;
wire  _GEN2818 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2819 = io_x[11] ? _GEN2818 : _GEN207;
wire  _GEN2820 = io_x[3] ? _GEN2819 : _GEN209;
wire  _GEN2821 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2822 = io_x[11] ? _GEN2821 : _GEN214;
wire  _GEN2823 = io_x[3] ? _GEN2822 : _GEN216;
wire  _GEN2824 = io_x[7] ? _GEN2823 : _GEN2820;
wire  _GEN2825 = io_x[2] ? _GEN2824 : _GEN2817;
wire  _GEN2826 = io_x[17] ? _GEN2825 : _GEN2816;
wire  _GEN2827 = io_x[15] ? _GEN2826 : _GEN2813;
wire  _GEN2828 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2829 = io_x[7] ? _GEN203 : _GEN2828;
wire  _GEN2830 = io_x[2] ? _GEN2829 : _GEN233;
wire  _GEN2831 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2832 = io_x[3] ? _GEN2831 : _GEN216;
wire  _GEN2833 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2834 = io_x[3] ? _GEN2833 : _GEN216;
wire  _GEN2835 = io_x[7] ? _GEN2834 : _GEN2832;
wire  _GEN2836 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2837 = io_x[3] ? _GEN2836 : _GEN209;
wire  _GEN2838 = io_x[7] ? _GEN2837 : _GEN203;
wire  _GEN2839 = io_x[2] ? _GEN2838 : _GEN2835;
wire  _GEN2840 = io_x[17] ? _GEN2839 : _GEN2830;
wire  _GEN2841 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN2842 = io_x[7] ? _GEN203 : _GEN2841;
wire  _GEN2843 = io_x[2] ? _GEN2842 : _GEN202;
wire  _GEN2844 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN2845 = io_x[7] ? _GEN2844 : _GEN203;
wire  _GEN2846 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2847 = io_x[3] ? _GEN216 : _GEN2846;
wire  _GEN2848 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2849 = io_x[3] ? _GEN2848 : _GEN216;
wire  _GEN2850 = io_x[7] ? _GEN2849 : _GEN2847;
wire  _GEN2851 = io_x[2] ? _GEN2850 : _GEN2845;
wire  _GEN2852 = io_x[17] ? _GEN2851 : _GEN2843;
wire  _GEN2853 = io_x[15] ? _GEN2852 : _GEN2840;
wire  _GEN2854 = io_x[12] ? _GEN2853 : _GEN2827;
wire  _GEN2855 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2856 = io_x[3] ? _GEN209 : _GEN2855;
wire  _GEN2857 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2858 = io_x[7] ? _GEN2857 : _GEN2856;
wire  _GEN2859 = io_x[2] ? _GEN2858 : _GEN233;
wire  _GEN2860 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2861 = io_x[3] ? _GEN2860 : _GEN216;
wire  _GEN2862 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2863 = io_x[3] ? _GEN2862 : _GEN216;
wire  _GEN2864 = io_x[7] ? _GEN2863 : _GEN2861;
wire  _GEN2865 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2866 = io_x[11] ? _GEN214 : _GEN2865;
wire  _GEN2867 = io_x[3] ? _GEN209 : _GEN2866;
wire  _GEN2868 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2869 = io_x[7] ? _GEN2868 : _GEN2867;
wire  _GEN2870 = io_x[2] ? _GEN2869 : _GEN2864;
wire  _GEN2871 = io_x[17] ? _GEN2870 : _GEN2859;
wire  _GEN2872 = io_x[2] ? _GEN233 : _GEN202;
wire  _GEN2873 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2874 = io_x[3] ? _GEN2873 : _GEN216;
wire  _GEN2875 = io_x[7] ? _GEN2874 : _GEN203;
wire  _GEN2876 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2877 = io_x[11] ? _GEN214 : _GEN2876;
wire  _GEN2878 = io_x[3] ? _GEN2877 : _GEN209;
wire  _GEN2879 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2880 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2881 = io_x[3] ? _GEN2880 : _GEN2879;
wire  _GEN2882 = io_x[7] ? _GEN2881 : _GEN2878;
wire  _GEN2883 = io_x[2] ? _GEN2882 : _GEN2875;
wire  _GEN2884 = io_x[17] ? _GEN2883 : _GEN2872;
wire  _GEN2885 = io_x[15] ? _GEN2884 : _GEN2871;
wire  _GEN2886 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2887 = io_x[11] ? _GEN214 : _GEN2886;
wire  _GEN2888 = io_x[3] ? _GEN2887 : _GEN216;
wire  _GEN2889 = io_x[7] ? _GEN2888 : _GEN203;
wire  _GEN2890 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2891 = io_x[11] ? _GEN2890 : _GEN214;
wire  _GEN2892 = io_x[3] ? _GEN2891 : _GEN209;
wire  _GEN2893 = io_x[7] ? _GEN2892 : _GEN203;
wire  _GEN2894 = io_x[2] ? _GEN2893 : _GEN2889;
wire  _GEN2895 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2896 = io_x[11] ? _GEN214 : _GEN2895;
wire  _GEN2897 = io_x[3] ? _GEN2896 : _GEN216;
wire  _GEN2898 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2899 = io_x[3] ? _GEN2898 : _GEN216;
wire  _GEN2900 = io_x[7] ? _GEN2899 : _GEN2897;
wire  _GEN2901 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2902 = io_x[11] ? _GEN214 : _GEN2901;
wire  _GEN2903 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2904 = io_x[11] ? _GEN214 : _GEN2903;
wire  _GEN2905 = io_x[3] ? _GEN2904 : _GEN2902;
wire  _GEN2906 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2907 = io_x[3] ? _GEN216 : _GEN2906;
wire  _GEN2908 = io_x[7] ? _GEN2907 : _GEN2905;
wire  _GEN2909 = io_x[2] ? _GEN2908 : _GEN2900;
wire  _GEN2910 = io_x[17] ? _GEN2909 : _GEN2894;
wire  _GEN2911 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2912 = io_x[11] ? _GEN2911 : _GEN214;
wire  _GEN2913 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2914 = io_x[3] ? _GEN2913 : _GEN2912;
wire  _GEN2915 = io_x[7] ? _GEN2914 : _GEN203;
wire  _GEN2916 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2917 = io_x[3] ? _GEN2916 : _GEN216;
wire  _GEN2918 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2919 = io_x[11] ? _GEN2918 : _GEN214;
wire  _GEN2920 = io_x[3] ? _GEN2919 : _GEN216;
wire  _GEN2921 = io_x[7] ? _GEN2920 : _GEN2917;
wire  _GEN2922 = io_x[2] ? _GEN2921 : _GEN2915;
wire  _GEN2923 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2924 = io_x[11] ? _GEN2923 : _GEN214;
wire  _GEN2925 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2926 = io_x[11] ? _GEN2925 : _GEN214;
wire  _GEN2927 = io_x[3] ? _GEN2926 : _GEN2924;
wire  _GEN2928 = io_x[7] ? _GEN2927 : _GEN241;
wire  _GEN2929 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2930 = io_x[11] ? _GEN207 : _GEN2929;
wire  _GEN2931 = io_x[3] ? _GEN209 : _GEN2930;
wire  _GEN2932 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2933 = io_x[11] ? _GEN2932 : _GEN214;
wire  _GEN2934 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2935 = io_x[11] ? _GEN2934 : _GEN214;
wire  _GEN2936 = io_x[3] ? _GEN2935 : _GEN2933;
wire  _GEN2937 = io_x[7] ? _GEN2936 : _GEN2931;
wire  _GEN2938 = io_x[2] ? _GEN2937 : _GEN2928;
wire  _GEN2939 = io_x[17] ? _GEN2938 : _GEN2922;
wire  _GEN2940 = io_x[15] ? _GEN2939 : _GEN2910;
wire  _GEN2941 = io_x[12] ? _GEN2940 : _GEN2885;
wire  _GEN2942 = io_x[10] ? _GEN2941 : _GEN2854;
wire  _GEN2943 = io_x[7] ? _GEN203 : _GEN241;
wire  _GEN2944 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2945 = io_x[11] ? _GEN2944 : _GEN214;
wire  _GEN2946 = io_x[3] ? _GEN216 : _GEN2945;
wire  _GEN2947 = io_x[7] ? _GEN241 : _GEN2946;
wire  _GEN2948 = io_x[2] ? _GEN2947 : _GEN2943;
wire  _GEN2949 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2950 = io_x[3] ? _GEN209 : _GEN2949;
wire  _GEN2951 = io_x[7] ? _GEN203 : _GEN2950;
wire  _GEN2952 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2953 = io_x[11] ? _GEN2952 : _GEN214;
wire  _GEN2954 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2955 = io_x[3] ? _GEN2954 : _GEN2953;
wire  _GEN2956 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2957 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2958 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2959 = io_x[11] ? _GEN2958 : _GEN2957;
wire  _GEN2960 = io_x[3] ? _GEN2959 : _GEN2956;
wire  _GEN2961 = io_x[7] ? _GEN2960 : _GEN2955;
wire  _GEN2962 = io_x[2] ? _GEN2961 : _GEN2951;
wire  _GEN2963 = io_x[17] ? _GEN2962 : _GEN2948;
wire  _GEN2964 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN2965 = io_x[11] ? _GEN2964 : _GEN214;
wire  _GEN2966 = io_x[3] ? _GEN216 : _GEN2965;
wire  _GEN2967 = io_x[7] ? _GEN203 : _GEN2966;
wire  _GEN2968 = io_x[2] ? _GEN2967 : _GEN233;
wire  _GEN2969 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2970 = io_x[11] ? _GEN2969 : _GEN214;
wire  _GEN2971 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2972 = io_x[3] ? _GEN2971 : _GEN2970;
wire  _GEN2973 = io_x[7] ? _GEN2972 : _GEN203;
wire  _GEN2974 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2975 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2976 = io_x[3] ? _GEN2975 : _GEN2974;
wire  _GEN2977 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2978 = io_x[3] ? _GEN2977 : _GEN216;
wire  _GEN2979 = io_x[7] ? _GEN2978 : _GEN2976;
wire  _GEN2980 = io_x[2] ? _GEN2979 : _GEN2973;
wire  _GEN2981 = io_x[17] ? _GEN2980 : _GEN2968;
wire  _GEN2982 = io_x[15] ? _GEN2981 : _GEN2963;
wire  _GEN2983 = io_x[3] ? _GEN209 : _GEN216;
wire  _GEN2984 = io_x[7] ? _GEN203 : _GEN2983;
wire  _GEN2985 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN2986 = io_x[11] ? _GEN2985 : _GEN214;
wire  _GEN2987 = io_x[3] ? _GEN209 : _GEN2986;
wire  _GEN2988 = io_x[7] ? _GEN241 : _GEN2987;
wire  _GEN2989 = io_x[2] ? _GEN2988 : _GEN2984;
wire  _GEN2990 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2991 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2992 = io_x[3] ? _GEN2991 : _GEN2990;
wire  _GEN2993 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN2994 = io_x[3] ? _GEN2993 : _GEN209;
wire  _GEN2995 = io_x[7] ? _GEN2994 : _GEN2992;
wire  _GEN2996 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2997 = io_x[3] ? _GEN2996 : _GEN216;
wire  _GEN2998 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN2999 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3000 = io_x[11] ? _GEN214 : _GEN2999;
wire  _GEN3001 = io_x[3] ? _GEN3000 : _GEN2998;
wire  _GEN3002 = io_x[7] ? _GEN3001 : _GEN2997;
wire  _GEN3003 = io_x[2] ? _GEN3002 : _GEN2995;
wire  _GEN3004 = io_x[17] ? _GEN3003 : _GEN2989;
wire  _GEN3005 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN3006 = io_x[7] ? _GEN3005 : _GEN203;
wire  _GEN3007 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3008 = io_x[11] ? _GEN3007 : _GEN207;
wire  _GEN3009 = io_x[3] ? _GEN216 : _GEN3008;
wire  _GEN3010 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN3011 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3012 = io_x[11] ? _GEN3011 : _GEN214;
wire  _GEN3013 = io_x[3] ? _GEN3012 : _GEN3010;
wire  _GEN3014 = io_x[7] ? _GEN3013 : _GEN3009;
wire  _GEN3015 = io_x[2] ? _GEN3014 : _GEN3006;
wire  _GEN3016 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN3017 = io_x[3] ? _GEN3016 : _GEN216;
wire  _GEN3018 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3019 = io_x[11] ? _GEN3018 : _GEN214;
wire  _GEN3020 = io_x[3] ? _GEN209 : _GEN3019;
wire  _GEN3021 = io_x[7] ? _GEN3020 : _GEN3017;
wire  _GEN3022 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3023 = io_x[11] ? _GEN214 : _GEN3022;
wire  _GEN3024 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3025 = io_x[11] ? _GEN214 : _GEN3024;
wire  _GEN3026 = io_x[3] ? _GEN3025 : _GEN3023;
wire  _GEN3027 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3028 = io_x[11] ? _GEN3027 : _GEN207;
wire  _GEN3029 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3030 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3031 = io_x[11] ? _GEN3030 : _GEN3029;
wire  _GEN3032 = io_x[3] ? _GEN3031 : _GEN3028;
wire  _GEN3033 = io_x[7] ? _GEN3032 : _GEN3026;
wire  _GEN3034 = io_x[2] ? _GEN3033 : _GEN3021;
wire  _GEN3035 = io_x[17] ? _GEN3034 : _GEN3015;
wire  _GEN3036 = io_x[15] ? _GEN3035 : _GEN3004;
wire  _GEN3037 = io_x[12] ? _GEN3036 : _GEN2982;
wire  _GEN3038 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN3039 = io_x[3] ? _GEN216 : _GEN3038;
wire  _GEN3040 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN3041 = io_x[3] ? _GEN216 : _GEN3040;
wire  _GEN3042 = io_x[7] ? _GEN3041 : _GEN3039;
wire  _GEN3043 = io_x[2] ? _GEN3042 : _GEN202;
wire  _GEN3044 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN3045 = io_x[3] ? _GEN3044 : _GEN209;
wire  _GEN3046 = io_x[7] ? _GEN3045 : _GEN241;
wire  _GEN3047 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN3048 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN3049 = io_x[3] ? _GEN3048 : _GEN3047;
wire  _GEN3050 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3051 = io_x[11] ? _GEN3050 : _GEN214;
wire  _GEN3052 = io_x[3] ? _GEN3051 : _GEN216;
wire  _GEN3053 = io_x[7] ? _GEN3052 : _GEN3049;
wire  _GEN3054 = io_x[2] ? _GEN3053 : _GEN3046;
wire  _GEN3055 = io_x[17] ? _GEN3054 : _GEN3043;
wire  _GEN3056 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN3057 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN3058 = io_x[3] ? _GEN3057 : _GEN209;
wire  _GEN3059 = io_x[7] ? _GEN3058 : _GEN3056;
wire  _GEN3060 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3061 = io_x[11] ? _GEN3060 : _GEN214;
wire  _GEN3062 = io_x[3] ? _GEN216 : _GEN3061;
wire  _GEN3063 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3064 = io_x[11] ? _GEN3063 : _GEN214;
wire  _GEN3065 = io_x[3] ? _GEN3064 : _GEN216;
wire  _GEN3066 = io_x[7] ? _GEN3065 : _GEN3062;
wire  _GEN3067 = io_x[2] ? _GEN3066 : _GEN3059;
wire  _GEN3068 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3069 = io_x[11] ? _GEN3068 : _GEN214;
wire  _GEN3070 = io_x[3] ? _GEN3069 : _GEN209;
wire  _GEN3071 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN3072 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3073 = io_x[11] ? _GEN3072 : _GEN214;
wire  _GEN3074 = io_x[3] ? _GEN3073 : _GEN3071;
wire  _GEN3075 = io_x[7] ? _GEN3074 : _GEN3070;
wire  _GEN3076 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3077 = io_x[11] ? _GEN3076 : _GEN214;
wire  _GEN3078 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3079 = io_x[11] ? _GEN3078 : _GEN207;
wire  _GEN3080 = io_x[3] ? _GEN3079 : _GEN3077;
wire  _GEN3081 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3082 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3083 = io_x[11] ? _GEN3082 : _GEN3081;
wire  _GEN3084 = io_x[3] ? _GEN3083 : _GEN209;
wire  _GEN3085 = io_x[7] ? _GEN3084 : _GEN3080;
wire  _GEN3086 = io_x[2] ? _GEN3085 : _GEN3075;
wire  _GEN3087 = io_x[17] ? _GEN3086 : _GEN3067;
wire  _GEN3088 = io_x[15] ? _GEN3087 : _GEN3055;
wire  _GEN3089 = io_x[3] ? _GEN216 : _GEN209;
wire  _GEN3090 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3091 = io_x[11] ? _GEN3090 : _GEN214;
wire  _GEN3092 = io_x[3] ? _GEN3091 : _GEN216;
wire  _GEN3093 = io_x[7] ? _GEN3092 : _GEN3089;
wire  _GEN3094 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3095 = io_x[11] ? _GEN214 : _GEN3094;
wire  _GEN3096 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3097 = io_x[11] ? _GEN207 : _GEN3096;
wire  _GEN3098 = io_x[3] ? _GEN3097 : _GEN3095;
wire  _GEN3099 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN3100 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3101 = io_x[11] ? _GEN3100 : _GEN214;
wire  _GEN3102 = io_x[3] ? _GEN3101 : _GEN3099;
wire  _GEN3103 = io_x[7] ? _GEN3102 : _GEN3098;
wire  _GEN3104 = io_x[2] ? _GEN3103 : _GEN3093;
wire  _GEN3105 = io_x[11] ? _GEN214 : _GEN207;
wire  _GEN3106 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3107 = io_x[11] ? _GEN214 : _GEN3106;
wire  _GEN3108 = io_x[3] ? _GEN3107 : _GEN3105;
wire  _GEN3109 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3110 = io_x[11] ? _GEN207 : _GEN3109;
wire  _GEN3111 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3112 = io_x[11] ? _GEN3111 : _GEN207;
wire  _GEN3113 = io_x[3] ? _GEN3112 : _GEN3110;
wire  _GEN3114 = io_x[7] ? _GEN3113 : _GEN3108;
wire  _GEN3115 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3116 = io_x[11] ? _GEN214 : _GEN3115;
wire  _GEN3117 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3118 = io_x[11] ? _GEN207 : _GEN3117;
wire  _GEN3119 = io_x[3] ? _GEN3118 : _GEN3116;
wire  _GEN3120 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3121 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3122 = io_x[11] ? _GEN3121 : _GEN3120;
wire  _GEN3123 = io_x[3] ? _GEN3122 : _GEN216;
wire  _GEN3124 = io_x[7] ? _GEN3123 : _GEN3119;
wire  _GEN3125 = io_x[2] ? _GEN3124 : _GEN3114;
wire  _GEN3126 = io_x[17] ? _GEN3125 : _GEN3104;
wire  _GEN3127 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3128 = io_x[11] ? _GEN3127 : _GEN207;
wire  _GEN3129 = io_x[3] ? _GEN3128 : _GEN209;
wire  _GEN3130 = io_x[7] ? _GEN3129 : _GEN241;
wire  _GEN3131 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3132 = io_x[11] ? _GEN207 : _GEN3131;
wire  _GEN3133 = io_x[3] ? _GEN216 : _GEN3132;
wire  _GEN3134 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3135 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3136 = io_x[11] ? _GEN3135 : _GEN3134;
wire  _GEN3137 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3138 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3139 = io_x[11] ? _GEN3138 : _GEN3137;
wire  _GEN3140 = io_x[3] ? _GEN3139 : _GEN3136;
wire  _GEN3141 = io_x[7] ? _GEN3140 : _GEN3133;
wire  _GEN3142 = io_x[2] ? _GEN3141 : _GEN3130;
wire  _GEN3143 = io_x[11] ? _GEN207 : _GEN214;
wire  _GEN3144 = io_x[3] ? _GEN209 : _GEN3143;
wire  _GEN3145 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3146 = io_x[11] ? _GEN3145 : _GEN207;
wire  _GEN3147 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3148 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3149 = io_x[11] ? _GEN3148 : _GEN3147;
wire  _GEN3150 = io_x[3] ? _GEN3149 : _GEN3146;
wire  _GEN3151 = io_x[7] ? _GEN3150 : _GEN3144;
wire  _GEN3152 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3153 = io_x[11] ? _GEN207 : _GEN3152;
wire  _GEN3154 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3155 = io_x[11] ? _GEN3154 : _GEN207;
wire  _GEN3156 = io_x[3] ? _GEN3155 : _GEN3153;
wire  _GEN3157 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3158 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3159 = io_x[11] ? _GEN3158 : _GEN3157;
wire  _GEN3160 = io_x[28] ? _GEN205 : _GEN204;
wire  _GEN3161 = io_x[28] ? _GEN204 : _GEN205;
wire  _GEN3162 = io_x[11] ? _GEN3161 : _GEN3160;
wire  _GEN3163 = io_x[3] ? _GEN3162 : _GEN3159;
wire  _GEN3164 = io_x[7] ? _GEN3163 : _GEN3156;
wire  _GEN3165 = io_x[2] ? _GEN3164 : _GEN3151;
wire  _GEN3166 = io_x[17] ? _GEN3165 : _GEN3142;
wire  _GEN3167 = io_x[15] ? _GEN3166 : _GEN3126;
wire  _GEN3168 = io_x[12] ? _GEN3167 : _GEN3088;
wire  _GEN3169 = io_x[10] ? _GEN3168 : _GEN3037;
wire  _GEN3170 = io_x[4] ? _GEN3169 : _GEN2942;
wire  _GEN3171 = io_x[8] ? _GEN3170 : _GEN2797;
wire  _GEN3172 = io_x[29] ? _GEN3171 : _GEN2540;
wire  _GEN3173 = io_x[23] ? _GEN3172 : _GEN1732;
assign io_y[8] = _GEN3173;
wire  _GEN3174 = 1'b1;
wire  _GEN3175 = 1'b0;
wire  _GEN3176 = 1'b1;
wire  _GEN3177 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3178 = 1'b1;
wire  _GEN3179 = io_x[10] ? _GEN3178 : _GEN3177;
wire  _GEN3180 = 1'b1;
wire  _GEN3181 = io_x[24] ? _GEN3180 : _GEN3179;
wire  _GEN3182 = io_x[17] ? _GEN3181 : _GEN3174;
wire  _GEN3183 = 1'b0;
wire  _GEN3184 = 1'b0;
wire  _GEN3185 = 1'b1;
wire  _GEN3186 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3187 = io_x[14] ? _GEN3186 : _GEN3176;
wire  _GEN3188 = io_x[10] ? _GEN3187 : _GEN3183;
wire  _GEN3189 = io_x[24] ? _GEN3180 : _GEN3188;
wire  _GEN3190 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3191 = io_x[14] ? _GEN3190 : _GEN3176;
wire  _GEN3192 = io_x[10] ? _GEN3191 : _GEN3183;
wire  _GEN3193 = io_x[24] ? _GEN3180 : _GEN3192;
wire  _GEN3194 = io_x[17] ? _GEN3193 : _GEN3189;
wire  _GEN3195 = io_x[12] ? _GEN3194 : _GEN3182;
wire  _GEN3196 = 1'b0;
wire  _GEN3197 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3198 = io_x[24] ? _GEN3197 : _GEN3196;
wire  _GEN3199 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3200 = io_x[14] ? _GEN3199 : _GEN3176;
wire  _GEN3201 = io_x[10] ? _GEN3200 : _GEN3183;
wire  _GEN3202 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3203 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3204 = io_x[14] ? _GEN3203 : _GEN3202;
wire  _GEN3205 = io_x[10] ? _GEN3183 : _GEN3204;
wire  _GEN3206 = io_x[24] ? _GEN3205 : _GEN3201;
wire  _GEN3207 = io_x[17] ? _GEN3206 : _GEN3198;
wire  _GEN3208 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3209 = io_x[10] ? _GEN3208 : _GEN3178;
wire  _GEN3210 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3211 = io_x[24] ? _GEN3210 : _GEN3209;
wire  _GEN3212 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3213 = io_x[14] ? _GEN3212 : _GEN3176;
wire  _GEN3214 = io_x[10] ? _GEN3213 : _GEN3178;
wire  _GEN3215 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3216 = io_x[14] ? _GEN3215 : _GEN3176;
wire  _GEN3217 = io_x[10] ? _GEN3183 : _GEN3216;
wire  _GEN3218 = io_x[24] ? _GEN3217 : _GEN3214;
wire  _GEN3219 = io_x[17] ? _GEN3218 : _GEN3211;
wire  _GEN3220 = io_x[12] ? _GEN3219 : _GEN3207;
wire  _GEN3221 = io_x[2] ? _GEN3220 : _GEN3195;
wire  _GEN3222 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3223 = io_x[10] ? _GEN3222 : _GEN3178;
wire  _GEN3224 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3225 = io_x[10] ? _GEN3224 : _GEN3178;
wire  _GEN3226 = io_x[24] ? _GEN3225 : _GEN3223;
wire  _GEN3227 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3228 = io_x[14] ? _GEN3227 : _GEN3175;
wire  _GEN3229 = io_x[10] ? _GEN3228 : _GEN3178;
wire  _GEN3230 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3231 = io_x[10] ? _GEN3230 : _GEN3178;
wire  _GEN3232 = io_x[24] ? _GEN3231 : _GEN3229;
wire  _GEN3233 = io_x[17] ? _GEN3232 : _GEN3226;
wire  _GEN3234 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3235 = io_x[14] ? _GEN3234 : _GEN3176;
wire  _GEN3236 = io_x[10] ? _GEN3235 : _GEN3183;
wire  _GEN3237 = io_x[24] ? _GEN3180 : _GEN3236;
wire  _GEN3238 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3239 = io_x[10] ? _GEN3238 : _GEN3183;
wire  _GEN3240 = io_x[24] ? _GEN3196 : _GEN3239;
wire  _GEN3241 = io_x[17] ? _GEN3240 : _GEN3237;
wire  _GEN3242 = io_x[12] ? _GEN3241 : _GEN3233;
wire  _GEN3243 = 1'b0;
wire  _GEN3244 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3245 = io_x[14] ? _GEN3244 : _GEN3176;
wire  _GEN3246 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3247 = io_x[14] ? _GEN3246 : _GEN3176;
wire  _GEN3248 = io_x[10] ? _GEN3247 : _GEN3245;
wire  _GEN3249 = io_x[24] ? _GEN3196 : _GEN3248;
wire  _GEN3250 = io_x[17] ? _GEN3249 : _GEN3243;
wire  _GEN3251 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3252 = io_x[14] ? _GEN3251 : _GEN3176;
wire  _GEN3253 = io_x[10] ? _GEN3252 : _GEN3178;
wire  _GEN3254 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3255 = io_x[24] ? _GEN3254 : _GEN3253;
wire  _GEN3256 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3257 = io_x[14] ? _GEN3256 : _GEN3175;
wire  _GEN3258 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3259 = io_x[10] ? _GEN3258 : _GEN3257;
wire  _GEN3260 = io_x[24] ? _GEN3259 : _GEN3196;
wire  _GEN3261 = io_x[17] ? _GEN3260 : _GEN3255;
wire  _GEN3262 = io_x[12] ? _GEN3261 : _GEN3250;
wire  _GEN3263 = io_x[2] ? _GEN3262 : _GEN3242;
wire  _GEN3264 = io_x[9] ? _GEN3263 : _GEN3221;
wire  _GEN3265 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3266 = io_x[24] ? _GEN3196 : _GEN3265;
wire  _GEN3267 = io_x[17] ? _GEN3266 : _GEN3243;
wire  _GEN3268 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3269 = io_x[14] ? _GEN3176 : _GEN3268;
wire  _GEN3270 = io_x[10] ? _GEN3183 : _GEN3269;
wire  _GEN3271 = io_x[24] ? _GEN3180 : _GEN3270;
wire  _GEN3272 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3273 = io_x[14] ? _GEN3176 : _GEN3272;
wire  _GEN3274 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3275 = io_x[10] ? _GEN3274 : _GEN3273;
wire  _GEN3276 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3277 = io_x[14] ? _GEN3276 : _GEN3176;
wire  _GEN3278 = io_x[10] ? _GEN3277 : _GEN3178;
wire  _GEN3279 = io_x[24] ? _GEN3278 : _GEN3275;
wire  _GEN3280 = io_x[17] ? _GEN3279 : _GEN3271;
wire  _GEN3281 = io_x[12] ? _GEN3280 : _GEN3267;
wire  _GEN3282 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3283 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN3284 = io_x[24] ? _GEN3283 : _GEN3282;
wire  _GEN3285 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3286 = io_x[10] ? _GEN3285 : _GEN3183;
wire  _GEN3287 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3288 = io_x[10] ? _GEN3287 : _GEN3178;
wire  _GEN3289 = io_x[24] ? _GEN3288 : _GEN3286;
wire  _GEN3290 = io_x[17] ? _GEN3289 : _GEN3284;
wire  _GEN3291 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3292 = io_x[10] ? _GEN3291 : _GEN3183;
wire  _GEN3293 = io_x[24] ? _GEN3292 : _GEN3196;
wire  _GEN3294 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3295 = io_x[14] ? _GEN3294 : _GEN3175;
wire  _GEN3296 = io_x[10] ? _GEN3295 : _GEN3178;
wire  _GEN3297 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3298 = io_x[10] ? _GEN3297 : _GEN3178;
wire  _GEN3299 = io_x[24] ? _GEN3298 : _GEN3296;
wire  _GEN3300 = io_x[17] ? _GEN3299 : _GEN3293;
wire  _GEN3301 = io_x[12] ? _GEN3300 : _GEN3290;
wire  _GEN3302 = io_x[2] ? _GEN3301 : _GEN3281;
wire  _GEN3303 = io_x[24] ? _GEN3196 : _GEN3180;
wire  _GEN3304 = io_x[17] ? _GEN3303 : _GEN3174;
wire  _GEN3305 = io_x[24] ? _GEN3180 : _GEN3196;
wire  _GEN3306 = io_x[17] ? _GEN3305 : _GEN3174;
wire  _GEN3307 = io_x[12] ? _GEN3306 : _GEN3304;
wire  _GEN3308 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3309 = io_x[10] ? _GEN3308 : _GEN3178;
wire  _GEN3310 = io_x[24] ? _GEN3196 : _GEN3309;
wire  _GEN3311 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3312 = io_x[14] ? _GEN3311 : _GEN3176;
wire  _GEN3313 = io_x[10] ? _GEN3183 : _GEN3312;
wire  _GEN3314 = io_x[24] ? _GEN3180 : _GEN3313;
wire  _GEN3315 = io_x[17] ? _GEN3314 : _GEN3310;
wire  _GEN3316 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3317 = io_x[14] ? _GEN3316 : _GEN3176;
wire  _GEN3318 = io_x[10] ? _GEN3317 : _GEN3178;
wire  _GEN3319 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3320 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3321 = io_x[10] ? _GEN3320 : _GEN3319;
wire  _GEN3322 = io_x[24] ? _GEN3321 : _GEN3318;
wire  _GEN3323 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3324 = io_x[14] ? _GEN3323 : _GEN3176;
wire  _GEN3325 = io_x[10] ? _GEN3324 : _GEN3178;
wire  _GEN3326 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3327 = io_x[14] ? _GEN3175 : _GEN3326;
wire  _GEN3328 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3329 = io_x[10] ? _GEN3328 : _GEN3327;
wire  _GEN3330 = io_x[24] ? _GEN3329 : _GEN3325;
wire  _GEN3331 = io_x[17] ? _GEN3330 : _GEN3322;
wire  _GEN3332 = io_x[12] ? _GEN3331 : _GEN3315;
wire  _GEN3333 = io_x[2] ? _GEN3332 : _GEN3307;
wire  _GEN3334 = io_x[9] ? _GEN3333 : _GEN3302;
wire  _GEN3335 = io_x[13] ? _GEN3334 : _GEN3264;
wire  _GEN3336 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3337 = io_x[24] ? _GEN3180 : _GEN3336;
wire  _GEN3338 = io_x[17] ? _GEN3337 : _GEN3174;
wire  _GEN3339 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3340 = io_x[24] ? _GEN3180 : _GEN3339;
wire  _GEN3341 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3342 = io_x[14] ? _GEN3341 : _GEN3176;
wire  _GEN3343 = io_x[10] ? _GEN3183 : _GEN3342;
wire  _GEN3344 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3345 = io_x[24] ? _GEN3344 : _GEN3343;
wire  _GEN3346 = io_x[17] ? _GEN3345 : _GEN3340;
wire  _GEN3347 = io_x[12] ? _GEN3346 : _GEN3338;
wire  _GEN3348 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3349 = io_x[14] ? _GEN3348 : _GEN3176;
wire  _GEN3350 = io_x[10] ? _GEN3349 : _GEN3183;
wire  _GEN3351 = io_x[24] ? _GEN3180 : _GEN3350;
wire  _GEN3352 = io_x[17] ? _GEN3243 : _GEN3351;
wire  _GEN3353 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3354 = io_x[10] ? _GEN3353 : _GEN3178;
wire  _GEN3355 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3356 = io_x[14] ? _GEN3175 : _GEN3355;
wire  _GEN3357 = io_x[10] ? _GEN3356 : _GEN3178;
wire  _GEN3358 = io_x[24] ? _GEN3357 : _GEN3354;
wire  _GEN3359 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3360 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3361 = io_x[14] ? _GEN3360 : _GEN3359;
wire  _GEN3362 = io_x[10] ? _GEN3361 : _GEN3178;
wire  _GEN3363 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3364 = io_x[14] ? _GEN3175 : _GEN3363;
wire  _GEN3365 = io_x[10] ? _GEN3364 : _GEN3183;
wire  _GEN3366 = io_x[24] ? _GEN3365 : _GEN3362;
wire  _GEN3367 = io_x[17] ? _GEN3366 : _GEN3358;
wire  _GEN3368 = io_x[12] ? _GEN3367 : _GEN3352;
wire  _GEN3369 = io_x[2] ? _GEN3368 : _GEN3347;
wire  _GEN3370 = 1'b1;
wire  _GEN3371 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN3372 = io_x[24] ? _GEN3371 : _GEN3180;
wire  _GEN3373 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3374 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3375 = io_x[14] ? _GEN3374 : _GEN3373;
wire  _GEN3376 = io_x[10] ? _GEN3375 : _GEN3178;
wire  _GEN3377 = io_x[24] ? _GEN3180 : _GEN3376;
wire  _GEN3378 = io_x[17] ? _GEN3377 : _GEN3372;
wire  _GEN3379 = io_x[12] ? _GEN3378 : _GEN3370;
wire  _GEN3380 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3381 = io_x[24] ? _GEN3180 : _GEN3380;
wire  _GEN3382 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3383 = io_x[24] ? _GEN3382 : _GEN3196;
wire  _GEN3384 = io_x[17] ? _GEN3383 : _GEN3381;
wire  _GEN3385 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3386 = io_x[14] ? _GEN3385 : _GEN3176;
wire  _GEN3387 = io_x[10] ? _GEN3183 : _GEN3386;
wire  _GEN3388 = io_x[24] ? _GEN3196 : _GEN3387;
wire  _GEN3389 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3390 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3391 = io_x[14] ? _GEN3175 : _GEN3390;
wire  _GEN3392 = io_x[10] ? _GEN3391 : _GEN3389;
wire  _GEN3393 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3394 = io_x[10] ? _GEN3183 : _GEN3393;
wire  _GEN3395 = io_x[24] ? _GEN3394 : _GEN3392;
wire  _GEN3396 = io_x[17] ? _GEN3395 : _GEN3388;
wire  _GEN3397 = io_x[12] ? _GEN3396 : _GEN3384;
wire  _GEN3398 = io_x[2] ? _GEN3397 : _GEN3379;
wire  _GEN3399 = io_x[9] ? _GEN3398 : _GEN3369;
wire  _GEN3400 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3401 = io_x[14] ? _GEN3175 : _GEN3400;
wire  _GEN3402 = io_x[10] ? _GEN3401 : _GEN3178;
wire  _GEN3403 = io_x[24] ? _GEN3180 : _GEN3402;
wire  _GEN3404 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3405 = io_x[10] ? _GEN3404 : _GEN3178;
wire  _GEN3406 = io_x[24] ? _GEN3180 : _GEN3405;
wire  _GEN3407 = io_x[17] ? _GEN3406 : _GEN3403;
wire  _GEN3408 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3409 = io_x[14] ? _GEN3175 : _GEN3408;
wire  _GEN3410 = io_x[10] ? _GEN3409 : _GEN3178;
wire  _GEN3411 = io_x[24] ? _GEN3196 : _GEN3410;
wire  _GEN3412 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3413 = io_x[14] ? _GEN3176 : _GEN3412;
wire  _GEN3414 = io_x[10] ? _GEN3413 : _GEN3178;
wire  _GEN3415 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3416 = io_x[14] ? _GEN3415 : _GEN3175;
wire  _GEN3417 = io_x[10] ? _GEN3416 : _GEN3183;
wire  _GEN3418 = io_x[24] ? _GEN3417 : _GEN3414;
wire  _GEN3419 = io_x[17] ? _GEN3418 : _GEN3411;
wire  _GEN3420 = io_x[12] ? _GEN3419 : _GEN3407;
wire  _GEN3421 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3422 = io_x[10] ? _GEN3421 : _GEN3183;
wire  _GEN3423 = io_x[24] ? _GEN3422 : _GEN3196;
wire  _GEN3424 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3425 = io_x[14] ? _GEN3424 : _GEN3175;
wire  _GEN3426 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3427 = io_x[10] ? _GEN3426 : _GEN3425;
wire  _GEN3428 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN3429 = io_x[24] ? _GEN3428 : _GEN3427;
wire  _GEN3430 = io_x[17] ? _GEN3429 : _GEN3423;
wire  _GEN3431 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3432 = io_x[14] ? _GEN3431 : _GEN3176;
wire  _GEN3433 = io_x[10] ? _GEN3432 : _GEN3178;
wire  _GEN3434 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3435 = io_x[14] ? _GEN3434 : _GEN3176;
wire  _GEN3436 = io_x[10] ? _GEN3435 : _GEN3178;
wire  _GEN3437 = io_x[24] ? _GEN3436 : _GEN3433;
wire  _GEN3438 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3439 = io_x[14] ? _GEN3438 : _GEN3176;
wire  _GEN3440 = io_x[10] ? _GEN3439 : _GEN3178;
wire  _GEN3441 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3442 = io_x[10] ? _GEN3178 : _GEN3441;
wire  _GEN3443 = io_x[24] ? _GEN3442 : _GEN3440;
wire  _GEN3444 = io_x[17] ? _GEN3443 : _GEN3437;
wire  _GEN3445 = io_x[12] ? _GEN3444 : _GEN3430;
wire  _GEN3446 = io_x[2] ? _GEN3445 : _GEN3420;
wire  _GEN3447 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3448 = io_x[14] ? _GEN3175 : _GEN3447;
wire  _GEN3449 = io_x[10] ? _GEN3183 : _GEN3448;
wire  _GEN3450 = io_x[24] ? _GEN3180 : _GEN3449;
wire  _GEN3451 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3452 = io_x[14] ? _GEN3175 : _GEN3451;
wire  _GEN3453 = io_x[10] ? _GEN3178 : _GEN3452;
wire  _GEN3454 = io_x[24] ? _GEN3180 : _GEN3453;
wire  _GEN3455 = io_x[17] ? _GEN3454 : _GEN3450;
wire  _GEN3456 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3457 = io_x[10] ? _GEN3456 : _GEN3183;
wire  _GEN3458 = io_x[24] ? _GEN3180 : _GEN3457;
wire  _GEN3459 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3460 = io_x[14] ? _GEN3459 : _GEN3175;
wire  _GEN3461 = io_x[10] ? _GEN3460 : _GEN3178;
wire  _GEN3462 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3463 = io_x[10] ? _GEN3183 : _GEN3462;
wire  _GEN3464 = io_x[24] ? _GEN3463 : _GEN3461;
wire  _GEN3465 = io_x[17] ? _GEN3464 : _GEN3458;
wire  _GEN3466 = io_x[12] ? _GEN3465 : _GEN3455;
wire  _GEN3467 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3468 = io_x[14] ? _GEN3467 : _GEN3176;
wire  _GEN3469 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3470 = io_x[14] ? _GEN3175 : _GEN3469;
wire  _GEN3471 = io_x[10] ? _GEN3470 : _GEN3468;
wire  _GEN3472 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3473 = io_x[10] ? _GEN3183 : _GEN3472;
wire  _GEN3474 = io_x[24] ? _GEN3473 : _GEN3471;
wire  _GEN3475 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3476 = io_x[10] ? _GEN3183 : _GEN3475;
wire  _GEN3477 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3478 = io_x[14] ? _GEN3176 : _GEN3477;
wire  _GEN3479 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3480 = io_x[10] ? _GEN3479 : _GEN3478;
wire  _GEN3481 = io_x[24] ? _GEN3480 : _GEN3476;
wire  _GEN3482 = io_x[17] ? _GEN3481 : _GEN3474;
wire  _GEN3483 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3484 = io_x[10] ? _GEN3483 : _GEN3178;
wire  _GEN3485 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3486 = io_x[14] ? _GEN3485 : _GEN3176;
wire  _GEN3487 = io_x[10] ? _GEN3486 : _GEN3183;
wire  _GEN3488 = io_x[24] ? _GEN3487 : _GEN3484;
wire  _GEN3489 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3490 = io_x[14] ? _GEN3489 : _GEN3176;
wire  _GEN3491 = io_x[10] ? _GEN3490 : _GEN3178;
wire  _GEN3492 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3493 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3494 = io_x[10] ? _GEN3493 : _GEN3492;
wire  _GEN3495 = io_x[24] ? _GEN3494 : _GEN3491;
wire  _GEN3496 = io_x[17] ? _GEN3495 : _GEN3488;
wire  _GEN3497 = io_x[12] ? _GEN3496 : _GEN3482;
wire  _GEN3498 = io_x[2] ? _GEN3497 : _GEN3466;
wire  _GEN3499 = io_x[9] ? _GEN3498 : _GEN3446;
wire  _GEN3500 = io_x[13] ? _GEN3499 : _GEN3399;
wire  _GEN3501 = io_x[7] ? _GEN3500 : _GEN3335;
wire  _GEN3502 = io_x[24] ? _GEN3180 : _GEN3196;
wire  _GEN3503 = io_x[17] ? _GEN3243 : _GEN3502;
wire  _GEN3504 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3505 = io_x[10] ? _GEN3178 : _GEN3504;
wire  _GEN3506 = io_x[24] ? _GEN3180 : _GEN3505;
wire  _GEN3507 = io_x[17] ? _GEN3243 : _GEN3506;
wire  _GEN3508 = io_x[12] ? _GEN3507 : _GEN3503;
wire  _GEN3509 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3510 = io_x[10] ? _GEN3509 : _GEN3178;
wire  _GEN3511 = io_x[24] ? _GEN3196 : _GEN3510;
wire  _GEN3512 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3513 = io_x[10] ? _GEN3183 : _GEN3512;
wire  _GEN3514 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3515 = io_x[14] ? _GEN3514 : _GEN3176;
wire  _GEN3516 = io_x[10] ? _GEN3515 : _GEN3183;
wire  _GEN3517 = io_x[24] ? _GEN3516 : _GEN3513;
wire  _GEN3518 = io_x[17] ? _GEN3517 : _GEN3511;
wire  _GEN3519 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3520 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3521 = io_x[14] ? _GEN3520 : _GEN3176;
wire  _GEN3522 = io_x[10] ? _GEN3521 : _GEN3519;
wire  _GEN3523 = io_x[24] ? _GEN3196 : _GEN3522;
wire  _GEN3524 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3525 = io_x[14] ? _GEN3176 : _GEN3524;
wire  _GEN3526 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3527 = io_x[14] ? _GEN3526 : _GEN3176;
wire  _GEN3528 = io_x[10] ? _GEN3527 : _GEN3525;
wire  _GEN3529 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3530 = io_x[10] ? _GEN3529 : _GEN3178;
wire  _GEN3531 = io_x[24] ? _GEN3530 : _GEN3528;
wire  _GEN3532 = io_x[17] ? _GEN3531 : _GEN3523;
wire  _GEN3533 = io_x[12] ? _GEN3532 : _GEN3518;
wire  _GEN3534 = io_x[2] ? _GEN3533 : _GEN3508;
wire  _GEN3535 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3536 = io_x[14] ? _GEN3535 : _GEN3176;
wire  _GEN3537 = io_x[10] ? _GEN3536 : _GEN3178;
wire  _GEN3538 = io_x[24] ? _GEN3196 : _GEN3537;
wire  _GEN3539 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3540 = io_x[14] ? _GEN3176 : _GEN3539;
wire  _GEN3541 = io_x[10] ? _GEN3540 : _GEN3178;
wire  _GEN3542 = io_x[24] ? _GEN3180 : _GEN3541;
wire  _GEN3543 = io_x[17] ? _GEN3542 : _GEN3538;
wire  _GEN3544 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3545 = io_x[14] ? _GEN3176 : _GEN3544;
wire  _GEN3546 = io_x[10] ? _GEN3183 : _GEN3545;
wire  _GEN3547 = io_x[24] ? _GEN3180 : _GEN3546;
wire  _GEN3548 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3549 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3550 = io_x[10] ? _GEN3549 : _GEN3548;
wire  _GEN3551 = io_x[24] ? _GEN3180 : _GEN3550;
wire  _GEN3552 = io_x[17] ? _GEN3551 : _GEN3547;
wire  _GEN3553 = io_x[12] ? _GEN3552 : _GEN3543;
wire  _GEN3554 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3555 = io_x[14] ? _GEN3554 : _GEN3176;
wire  _GEN3556 = io_x[10] ? _GEN3555 : _GEN3178;
wire  _GEN3557 = io_x[24] ? _GEN3556 : _GEN3180;
wire  _GEN3558 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3559 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3560 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3561 = io_x[14] ? _GEN3560 : _GEN3559;
wire  _GEN3562 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3563 = io_x[10] ? _GEN3562 : _GEN3561;
wire  _GEN3564 = io_x[24] ? _GEN3563 : _GEN3558;
wire  _GEN3565 = io_x[17] ? _GEN3564 : _GEN3557;
wire  _GEN3566 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3567 = io_x[10] ? _GEN3566 : _GEN3178;
wire  _GEN3568 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3569 = io_x[14] ? _GEN3568 : _GEN3176;
wire  _GEN3570 = io_x[10] ? _GEN3569 : _GEN3183;
wire  _GEN3571 = io_x[24] ? _GEN3570 : _GEN3567;
wire  _GEN3572 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3573 = io_x[14] ? _GEN3572 : _GEN3176;
wire  _GEN3574 = io_x[10] ? _GEN3573 : _GEN3178;
wire  _GEN3575 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3576 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3577 = io_x[14] ? _GEN3576 : _GEN3176;
wire  _GEN3578 = io_x[10] ? _GEN3577 : _GEN3575;
wire  _GEN3579 = io_x[24] ? _GEN3578 : _GEN3574;
wire  _GEN3580 = io_x[17] ? _GEN3579 : _GEN3571;
wire  _GEN3581 = io_x[12] ? _GEN3580 : _GEN3565;
wire  _GEN3582 = io_x[2] ? _GEN3581 : _GEN3553;
wire  _GEN3583 = io_x[9] ? _GEN3582 : _GEN3534;
wire  _GEN3584 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3585 = io_x[10] ? _GEN3178 : _GEN3584;
wire  _GEN3586 = io_x[24] ? _GEN3585 : _GEN3196;
wire  _GEN3587 = io_x[17] ? _GEN3586 : _GEN3174;
wire  _GEN3588 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3589 = io_x[14] ? _GEN3588 : _GEN3176;
wire  _GEN3590 = io_x[10] ? _GEN3589 : _GEN3178;
wire  _GEN3591 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3592 = io_x[24] ? _GEN3591 : _GEN3590;
wire  _GEN3593 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3594 = io_x[10] ? _GEN3593 : _GEN3178;
wire  _GEN3595 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3596 = io_x[14] ? _GEN3595 : _GEN3175;
wire  _GEN3597 = io_x[10] ? _GEN3596 : _GEN3178;
wire  _GEN3598 = io_x[24] ? _GEN3597 : _GEN3594;
wire  _GEN3599 = io_x[17] ? _GEN3598 : _GEN3592;
wire  _GEN3600 = io_x[12] ? _GEN3599 : _GEN3587;
wire  _GEN3601 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3602 = io_x[10] ? _GEN3601 : _GEN3178;
wire  _GEN3603 = io_x[24] ? _GEN3180 : _GEN3602;
wire  _GEN3604 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3605 = io_x[14] ? _GEN3604 : _GEN3176;
wire  _GEN3606 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3607 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3608 = io_x[14] ? _GEN3607 : _GEN3606;
wire  _GEN3609 = io_x[10] ? _GEN3608 : _GEN3605;
wire  _GEN3610 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3611 = io_x[10] ? _GEN3610 : _GEN3183;
wire  _GEN3612 = io_x[24] ? _GEN3611 : _GEN3609;
wire  _GEN3613 = io_x[17] ? _GEN3612 : _GEN3603;
wire  _GEN3614 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3615 = io_x[14] ? _GEN3176 : _GEN3614;
wire  _GEN3616 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3617 = io_x[14] ? _GEN3616 : _GEN3176;
wire  _GEN3618 = io_x[10] ? _GEN3617 : _GEN3615;
wire  _GEN3619 = io_x[24] ? _GEN3196 : _GEN3618;
wire  _GEN3620 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3621 = io_x[14] ? _GEN3620 : _GEN3175;
wire  _GEN3622 = io_x[10] ? _GEN3183 : _GEN3621;
wire  _GEN3623 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3624 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3625 = io_x[14] ? _GEN3624 : _GEN3176;
wire  _GEN3626 = io_x[10] ? _GEN3625 : _GEN3623;
wire  _GEN3627 = io_x[24] ? _GEN3626 : _GEN3622;
wire  _GEN3628 = io_x[17] ? _GEN3627 : _GEN3619;
wire  _GEN3629 = io_x[12] ? _GEN3628 : _GEN3613;
wire  _GEN3630 = io_x[2] ? _GEN3629 : _GEN3600;
wire  _GEN3631 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3632 = io_x[14] ? _GEN3631 : _GEN3176;
wire  _GEN3633 = io_x[10] ? _GEN3632 : _GEN3178;
wire  _GEN3634 = io_x[24] ? _GEN3196 : _GEN3633;
wire  _GEN3635 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3636 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3637 = io_x[14] ? _GEN3636 : _GEN3635;
wire  _GEN3638 = io_x[10] ? _GEN3637 : _GEN3183;
wire  _GEN3639 = io_x[24] ? _GEN3196 : _GEN3638;
wire  _GEN3640 = io_x[17] ? _GEN3639 : _GEN3634;
wire  _GEN3641 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3642 = io_x[24] ? _GEN3180 : _GEN3641;
wire  _GEN3643 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3644 = io_x[14] ? _GEN3643 : _GEN3176;
wire  _GEN3645 = io_x[10] ? _GEN3644 : _GEN3178;
wire  _GEN3646 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3647 = io_x[14] ? _GEN3646 : _GEN3175;
wire  _GEN3648 = io_x[10] ? _GEN3647 : _GEN3178;
wire  _GEN3649 = io_x[24] ? _GEN3648 : _GEN3645;
wire  _GEN3650 = io_x[17] ? _GEN3649 : _GEN3642;
wire  _GEN3651 = io_x[12] ? _GEN3650 : _GEN3640;
wire  _GEN3652 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN3653 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3654 = io_x[14] ? _GEN3176 : _GEN3653;
wire  _GEN3655 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3656 = io_x[14] ? _GEN3176 : _GEN3655;
wire  _GEN3657 = io_x[10] ? _GEN3656 : _GEN3654;
wire  _GEN3658 = io_x[24] ? _GEN3657 : _GEN3652;
wire  _GEN3659 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3660 = io_x[14] ? _GEN3176 : _GEN3659;
wire  _GEN3661 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3662 = io_x[14] ? _GEN3661 : _GEN3176;
wire  _GEN3663 = io_x[10] ? _GEN3662 : _GEN3660;
wire  _GEN3664 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3665 = io_x[14] ? _GEN3664 : _GEN3175;
wire  _GEN3666 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3667 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3668 = io_x[14] ? _GEN3667 : _GEN3666;
wire  _GEN3669 = io_x[10] ? _GEN3668 : _GEN3665;
wire  _GEN3670 = io_x[24] ? _GEN3669 : _GEN3663;
wire  _GEN3671 = io_x[17] ? _GEN3670 : _GEN3658;
wire  _GEN3672 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3673 = io_x[14] ? _GEN3672 : _GEN3176;
wire  _GEN3674 = io_x[10] ? _GEN3673 : _GEN3178;
wire  _GEN3675 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3676 = io_x[10] ? _GEN3675 : _GEN3178;
wire  _GEN3677 = io_x[24] ? _GEN3676 : _GEN3674;
wire  _GEN3678 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3679 = io_x[14] ? _GEN3678 : _GEN3175;
wire  _GEN3680 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3681 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3682 = io_x[14] ? _GEN3681 : _GEN3680;
wire  _GEN3683 = io_x[10] ? _GEN3682 : _GEN3679;
wire  _GEN3684 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3685 = io_x[14] ? _GEN3684 : _GEN3176;
wire  _GEN3686 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3687 = io_x[14] ? _GEN3686 : _GEN3176;
wire  _GEN3688 = io_x[10] ? _GEN3687 : _GEN3685;
wire  _GEN3689 = io_x[24] ? _GEN3688 : _GEN3683;
wire  _GEN3690 = io_x[17] ? _GEN3689 : _GEN3677;
wire  _GEN3691 = io_x[12] ? _GEN3690 : _GEN3671;
wire  _GEN3692 = io_x[2] ? _GEN3691 : _GEN3651;
wire  _GEN3693 = io_x[9] ? _GEN3692 : _GEN3630;
wire  _GEN3694 = io_x[13] ? _GEN3693 : _GEN3583;
wire  _GEN3695 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3696 = io_x[14] ? _GEN3695 : _GEN3176;
wire  _GEN3697 = io_x[10] ? _GEN3696 : _GEN3178;
wire  _GEN3698 = io_x[24] ? _GEN3180 : _GEN3697;
wire  _GEN3699 = io_x[17] ? _GEN3698 : _GEN3174;
wire  _GEN3700 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3701 = io_x[24] ? _GEN3700 : _GEN3180;
wire  _GEN3702 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3703 = io_x[14] ? _GEN3702 : _GEN3175;
wire  _GEN3704 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3705 = io_x[14] ? _GEN3176 : _GEN3704;
wire  _GEN3706 = io_x[10] ? _GEN3705 : _GEN3703;
wire  _GEN3707 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3708 = io_x[24] ? _GEN3707 : _GEN3706;
wire  _GEN3709 = io_x[17] ? _GEN3708 : _GEN3701;
wire  _GEN3710 = io_x[12] ? _GEN3709 : _GEN3699;
wire  _GEN3711 = io_x[24] ? _GEN3196 : _GEN3180;
wire  _GEN3712 = io_x[17] ? _GEN3711 : _GEN3174;
wire  _GEN3713 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3714 = io_x[14] ? _GEN3713 : _GEN3175;
wire  _GEN3715 = io_x[10] ? _GEN3714 : _GEN3178;
wire  _GEN3716 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3717 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3718 = io_x[14] ? _GEN3717 : _GEN3716;
wire  _GEN3719 = io_x[10] ? _GEN3718 : _GEN3183;
wire  _GEN3720 = io_x[24] ? _GEN3719 : _GEN3715;
wire  _GEN3721 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3722 = io_x[14] ? _GEN3721 : _GEN3175;
wire  _GEN3723 = io_x[10] ? _GEN3722 : _GEN3178;
wire  _GEN3724 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3725 = io_x[14] ? _GEN3176 : _GEN3724;
wire  _GEN3726 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3727 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3728 = io_x[14] ? _GEN3727 : _GEN3726;
wire  _GEN3729 = io_x[10] ? _GEN3728 : _GEN3725;
wire  _GEN3730 = io_x[24] ? _GEN3729 : _GEN3723;
wire  _GEN3731 = io_x[17] ? _GEN3730 : _GEN3720;
wire  _GEN3732 = io_x[12] ? _GEN3731 : _GEN3712;
wire  _GEN3733 = io_x[2] ? _GEN3732 : _GEN3710;
wire  _GEN3734 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3735 = io_x[24] ? _GEN3180 : _GEN3734;
wire  _GEN3736 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3737 = io_x[10] ? _GEN3736 : _GEN3183;
wire  _GEN3738 = io_x[24] ? _GEN3180 : _GEN3737;
wire  _GEN3739 = io_x[17] ? _GEN3738 : _GEN3735;
wire  _GEN3740 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN3741 = io_x[24] ? _GEN3180 : _GEN3740;
wire  _GEN3742 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3743 = io_x[14] ? _GEN3742 : _GEN3176;
wire  _GEN3744 = io_x[10] ? _GEN3743 : _GEN3178;
wire  _GEN3745 = io_x[24] ? _GEN3180 : _GEN3744;
wire  _GEN3746 = io_x[17] ? _GEN3745 : _GEN3741;
wire  _GEN3747 = io_x[12] ? _GEN3746 : _GEN3739;
wire  _GEN3748 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3749 = io_x[14] ? _GEN3175 : _GEN3748;
wire  _GEN3750 = io_x[10] ? _GEN3183 : _GEN3749;
wire  _GEN3751 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3752 = io_x[14] ? _GEN3751 : _GEN3176;
wire  _GEN3753 = io_x[10] ? _GEN3752 : _GEN3183;
wire  _GEN3754 = io_x[24] ? _GEN3753 : _GEN3750;
wire  _GEN3755 = io_x[17] ? _GEN3754 : _GEN3243;
wire  _GEN3756 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3757 = io_x[14] ? _GEN3756 : _GEN3176;
wire  _GEN3758 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3759 = io_x[14] ? _GEN3758 : _GEN3176;
wire  _GEN3760 = io_x[10] ? _GEN3759 : _GEN3757;
wire  _GEN3761 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3762 = io_x[14] ? _GEN3761 : _GEN3176;
wire  _GEN3763 = io_x[10] ? _GEN3762 : _GEN3178;
wire  _GEN3764 = io_x[24] ? _GEN3763 : _GEN3760;
wire  _GEN3765 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3766 = io_x[14] ? _GEN3765 : _GEN3176;
wire  _GEN3767 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3768 = io_x[14] ? _GEN3767 : _GEN3176;
wire  _GEN3769 = io_x[10] ? _GEN3768 : _GEN3766;
wire  _GEN3770 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3771 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3772 = io_x[14] ? _GEN3771 : _GEN3770;
wire  _GEN3773 = io_x[10] ? _GEN3772 : _GEN3178;
wire  _GEN3774 = io_x[24] ? _GEN3773 : _GEN3769;
wire  _GEN3775 = io_x[17] ? _GEN3774 : _GEN3764;
wire  _GEN3776 = io_x[12] ? _GEN3775 : _GEN3755;
wire  _GEN3777 = io_x[2] ? _GEN3776 : _GEN3747;
wire  _GEN3778 = io_x[9] ? _GEN3777 : _GEN3733;
wire  _GEN3779 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3780 = io_x[14] ? _GEN3779 : _GEN3176;
wire  _GEN3781 = io_x[10] ? _GEN3183 : _GEN3780;
wire  _GEN3782 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3783 = io_x[10] ? _GEN3178 : _GEN3782;
wire  _GEN3784 = io_x[24] ? _GEN3783 : _GEN3781;
wire  _GEN3785 = io_x[17] ? _GEN3784 : _GEN3174;
wire  _GEN3786 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3787 = io_x[24] ? _GEN3180 : _GEN3786;
wire  _GEN3788 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3789 = io_x[14] ? _GEN3788 : _GEN3176;
wire  _GEN3790 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3791 = io_x[14] ? _GEN3790 : _GEN3175;
wire  _GEN3792 = io_x[10] ? _GEN3791 : _GEN3789;
wire  _GEN3793 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN3794 = io_x[24] ? _GEN3793 : _GEN3792;
wire  _GEN3795 = io_x[17] ? _GEN3794 : _GEN3787;
wire  _GEN3796 = io_x[12] ? _GEN3795 : _GEN3785;
wire  _GEN3797 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3798 = io_x[14] ? _GEN3176 : _GEN3797;
wire  _GEN3799 = io_x[10] ? _GEN3798 : _GEN3178;
wire  _GEN3800 = io_x[24] ? _GEN3180 : _GEN3799;
wire  _GEN3801 = io_x[24] ? _GEN3180 : _GEN3196;
wire  _GEN3802 = io_x[17] ? _GEN3801 : _GEN3800;
wire  _GEN3803 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3804 = io_x[14] ? _GEN3175 : _GEN3803;
wire  _GEN3805 = io_x[10] ? _GEN3804 : _GEN3178;
wire  _GEN3806 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3807 = io_x[10] ? _GEN3806 : _GEN3178;
wire  _GEN3808 = io_x[24] ? _GEN3807 : _GEN3805;
wire  _GEN3809 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3810 = io_x[10] ? _GEN3809 : _GEN3178;
wire  _GEN3811 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3812 = io_x[10] ? _GEN3811 : _GEN3178;
wire  _GEN3813 = io_x[24] ? _GEN3812 : _GEN3810;
wire  _GEN3814 = io_x[17] ? _GEN3813 : _GEN3808;
wire  _GEN3815 = io_x[12] ? _GEN3814 : _GEN3802;
wire  _GEN3816 = io_x[2] ? _GEN3815 : _GEN3796;
wire  _GEN3817 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3818 = io_x[14] ? _GEN3176 : _GEN3817;
wire  _GEN3819 = io_x[10] ? _GEN3178 : _GEN3818;
wire  _GEN3820 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN3821 = io_x[24] ? _GEN3820 : _GEN3819;
wire  _GEN3822 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3823 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3824 = io_x[14] ? _GEN3823 : _GEN3822;
wire  _GEN3825 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3826 = io_x[14] ? _GEN3825 : _GEN3175;
wire  _GEN3827 = io_x[10] ? _GEN3826 : _GEN3824;
wire  _GEN3828 = io_x[24] ? _GEN3180 : _GEN3827;
wire  _GEN3829 = io_x[17] ? _GEN3828 : _GEN3821;
wire  _GEN3830 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3831 = io_x[14] ? _GEN3830 : _GEN3175;
wire  _GEN3832 = io_x[10] ? _GEN3831 : _GEN3178;
wire  _GEN3833 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3834 = io_x[10] ? _GEN3833 : _GEN3183;
wire  _GEN3835 = io_x[24] ? _GEN3834 : _GEN3832;
wire  _GEN3836 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3837 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3838 = io_x[14] ? _GEN3837 : _GEN3836;
wire  _GEN3839 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3840 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3841 = io_x[14] ? _GEN3840 : _GEN3839;
wire  _GEN3842 = io_x[10] ? _GEN3841 : _GEN3838;
wire  _GEN3843 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3844 = io_x[14] ? _GEN3843 : _GEN3176;
wire  _GEN3845 = io_x[10] ? _GEN3844 : _GEN3183;
wire  _GEN3846 = io_x[24] ? _GEN3845 : _GEN3842;
wire  _GEN3847 = io_x[17] ? _GEN3846 : _GEN3835;
wire  _GEN3848 = io_x[12] ? _GEN3847 : _GEN3829;
wire  _GEN3849 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3850 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3851 = io_x[14] ? _GEN3850 : _GEN3849;
wire  _GEN3852 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3853 = io_x[10] ? _GEN3852 : _GEN3851;
wire  _GEN3854 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3855 = io_x[14] ? _GEN3176 : _GEN3854;
wire  _GEN3856 = io_x[10] ? _GEN3178 : _GEN3855;
wire  _GEN3857 = io_x[24] ? _GEN3856 : _GEN3853;
wire  _GEN3858 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3859 = io_x[14] ? _GEN3858 : _GEN3176;
wire  _GEN3860 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3861 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3862 = io_x[14] ? _GEN3861 : _GEN3860;
wire  _GEN3863 = io_x[10] ? _GEN3862 : _GEN3859;
wire  _GEN3864 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3865 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3866 = io_x[14] ? _GEN3865 : _GEN3864;
wire  _GEN3867 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3868 = io_x[14] ? _GEN3175 : _GEN3867;
wire  _GEN3869 = io_x[10] ? _GEN3868 : _GEN3866;
wire  _GEN3870 = io_x[24] ? _GEN3869 : _GEN3863;
wire  _GEN3871 = io_x[17] ? _GEN3870 : _GEN3857;
wire  _GEN3872 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3873 = io_x[14] ? _GEN3176 : _GEN3872;
wire  _GEN3874 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3875 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3876 = io_x[14] ? _GEN3875 : _GEN3874;
wire  _GEN3877 = io_x[10] ? _GEN3876 : _GEN3873;
wire  _GEN3878 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3879 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3880 = io_x[14] ? _GEN3879 : _GEN3878;
wire  _GEN3881 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3882 = io_x[14] ? _GEN3881 : _GEN3176;
wire  _GEN3883 = io_x[10] ? _GEN3882 : _GEN3880;
wire  _GEN3884 = io_x[24] ? _GEN3883 : _GEN3877;
wire  _GEN3885 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3886 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3887 = io_x[14] ? _GEN3886 : _GEN3885;
wire  _GEN3888 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3889 = io_x[14] ? _GEN3888 : _GEN3176;
wire  _GEN3890 = io_x[10] ? _GEN3889 : _GEN3887;
wire  _GEN3891 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3892 = io_x[14] ? _GEN3176 : _GEN3891;
wire  _GEN3893 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3894 = io_x[14] ? _GEN3893 : _GEN3176;
wire  _GEN3895 = io_x[10] ? _GEN3894 : _GEN3892;
wire  _GEN3896 = io_x[24] ? _GEN3895 : _GEN3890;
wire  _GEN3897 = io_x[17] ? _GEN3896 : _GEN3884;
wire  _GEN3898 = io_x[12] ? _GEN3897 : _GEN3871;
wire  _GEN3899 = io_x[2] ? _GEN3898 : _GEN3848;
wire  _GEN3900 = io_x[9] ? _GEN3899 : _GEN3816;
wire  _GEN3901 = io_x[13] ? _GEN3900 : _GEN3778;
wire  _GEN3902 = io_x[7] ? _GEN3901 : _GEN3694;
wire  _GEN3903 = io_x[15] ? _GEN3902 : _GEN3501;
wire  _GEN3904 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3905 = io_x[14] ? _GEN3904 : _GEN3176;
wire  _GEN3906 = io_x[10] ? _GEN3905 : _GEN3178;
wire  _GEN3907 = io_x[24] ? _GEN3180 : _GEN3906;
wire  _GEN3908 = io_x[17] ? _GEN3907 : _GEN3174;
wire  _GEN3909 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN3910 = io_x[24] ? _GEN3909 : _GEN3180;
wire  _GEN3911 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3912 = io_x[10] ? _GEN3911 : _GEN3178;
wire  _GEN3913 = io_x[24] ? _GEN3196 : _GEN3912;
wire  _GEN3914 = io_x[17] ? _GEN3913 : _GEN3910;
wire  _GEN3915 = io_x[12] ? _GEN3914 : _GEN3908;
wire  _GEN3916 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3917 = io_x[14] ? _GEN3916 : _GEN3176;
wire  _GEN3918 = io_x[10] ? _GEN3917 : _GEN3178;
wire  _GEN3919 = io_x[24] ? _GEN3918 : _GEN3180;
wire  _GEN3920 = io_x[17] ? _GEN3919 : _GEN3243;
wire  _GEN3921 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3922 = io_x[14] ? _GEN3921 : _GEN3176;
wire  _GEN3923 = io_x[10] ? _GEN3922 : _GEN3178;
wire  _GEN3924 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN3925 = io_x[24] ? _GEN3924 : _GEN3923;
wire  _GEN3926 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3927 = io_x[14] ? _GEN3926 : _GEN3176;
wire  _GEN3928 = io_x[10] ? _GEN3183 : _GEN3927;
wire  _GEN3929 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3930 = io_x[14] ? _GEN3929 : _GEN3176;
wire  _GEN3931 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3932 = io_x[14] ? _GEN3931 : _GEN3175;
wire  _GEN3933 = io_x[10] ? _GEN3932 : _GEN3930;
wire  _GEN3934 = io_x[24] ? _GEN3933 : _GEN3928;
wire  _GEN3935 = io_x[17] ? _GEN3934 : _GEN3925;
wire  _GEN3936 = io_x[12] ? _GEN3935 : _GEN3920;
wire  _GEN3937 = io_x[2] ? _GEN3936 : _GEN3915;
wire  _GEN3938 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN3939 = io_x[24] ? _GEN3938 : _GEN3180;
wire  _GEN3940 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3941 = io_x[10] ? _GEN3940 : _GEN3178;
wire  _GEN3942 = io_x[24] ? _GEN3180 : _GEN3941;
wire  _GEN3943 = io_x[17] ? _GEN3942 : _GEN3939;
wire  _GEN3944 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3945 = io_x[10] ? _GEN3944 : _GEN3178;
wire  _GEN3946 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3947 = io_x[14] ? _GEN3946 : _GEN3176;
wire  _GEN3948 = io_x[10] ? _GEN3178 : _GEN3947;
wire  _GEN3949 = io_x[24] ? _GEN3948 : _GEN3945;
wire  _GEN3950 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3951 = io_x[14] ? _GEN3950 : _GEN3176;
wire  _GEN3952 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3953 = io_x[14] ? _GEN3952 : _GEN3175;
wire  _GEN3954 = io_x[10] ? _GEN3953 : _GEN3951;
wire  _GEN3955 = io_x[24] ? _GEN3180 : _GEN3954;
wire  _GEN3956 = io_x[17] ? _GEN3955 : _GEN3949;
wire  _GEN3957 = io_x[12] ? _GEN3956 : _GEN3943;
wire  _GEN3958 = 1'b0;
wire  _GEN3959 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3960 = io_x[14] ? _GEN3959 : _GEN3176;
wire  _GEN3961 = io_x[10] ? _GEN3960 : _GEN3183;
wire  _GEN3962 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3963 = io_x[10] ? _GEN3962 : _GEN3178;
wire  _GEN3964 = io_x[24] ? _GEN3963 : _GEN3961;
wire  _GEN3965 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3966 = io_x[14] ? _GEN3965 : _GEN3176;
wire  _GEN3967 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3968 = io_x[14] ? _GEN3967 : _GEN3176;
wire  _GEN3969 = io_x[10] ? _GEN3968 : _GEN3966;
wire  _GEN3970 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3971 = io_x[10] ? _GEN3178 : _GEN3970;
wire  _GEN3972 = io_x[24] ? _GEN3971 : _GEN3969;
wire  _GEN3973 = io_x[17] ? _GEN3972 : _GEN3964;
wire  _GEN3974 = io_x[12] ? _GEN3973 : _GEN3958;
wire  _GEN3975 = io_x[2] ? _GEN3974 : _GEN3957;
wire  _GEN3976 = io_x[9] ? _GEN3975 : _GEN3937;
wire  _GEN3977 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3978 = io_x[14] ? _GEN3176 : _GEN3977;
wire  _GEN3979 = io_x[10] ? _GEN3978 : _GEN3178;
wire  _GEN3980 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN3981 = io_x[24] ? _GEN3980 : _GEN3979;
wire  _GEN3982 = io_x[17] ? _GEN3981 : _GEN3174;
wire  _GEN3983 = io_x[24] ? _GEN3180 : _GEN3196;
wire  _GEN3984 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3985 = io_x[14] ? _GEN3984 : _GEN3176;
wire  _GEN3986 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN3987 = io_x[10] ? _GEN3986 : _GEN3985;
wire  _GEN3988 = io_x[24] ? _GEN3196 : _GEN3987;
wire  _GEN3989 = io_x[17] ? _GEN3988 : _GEN3983;
wire  _GEN3990 = io_x[12] ? _GEN3989 : _GEN3982;
wire  _GEN3991 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN3992 = io_x[10] ? _GEN3991 : _GEN3178;
wire  _GEN3993 = io_x[24] ? _GEN3992 : _GEN3196;
wire  _GEN3994 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN3995 = io_x[14] ? _GEN3994 : _GEN3176;
wire  _GEN3996 = io_x[10] ? _GEN3995 : _GEN3183;
wire  _GEN3997 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN3998 = io_x[14] ? _GEN3175 : _GEN3997;
wire  _GEN3999 = io_x[10] ? _GEN3998 : _GEN3178;
wire  _GEN4000 = io_x[24] ? _GEN3999 : _GEN3996;
wire  _GEN4001 = io_x[17] ? _GEN4000 : _GEN3993;
wire  _GEN4002 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4003 = io_x[10] ? _GEN4002 : _GEN3178;
wire  _GEN4004 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4005 = io_x[10] ? _GEN4004 : _GEN3178;
wire  _GEN4006 = io_x[24] ? _GEN4005 : _GEN4003;
wire  _GEN4007 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4008 = io_x[10] ? _GEN3183 : _GEN4007;
wire  _GEN4009 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4010 = io_x[10] ? _GEN4009 : _GEN3178;
wire  _GEN4011 = io_x[24] ? _GEN4010 : _GEN4008;
wire  _GEN4012 = io_x[17] ? _GEN4011 : _GEN4006;
wire  _GEN4013 = io_x[12] ? _GEN4012 : _GEN4001;
wire  _GEN4014 = io_x[2] ? _GEN4013 : _GEN3990;
wire  _GEN4015 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4016 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4017 = io_x[10] ? _GEN4016 : _GEN4015;
wire  _GEN4018 = io_x[24] ? _GEN4017 : _GEN3196;
wire  _GEN4019 = io_x[17] ? _GEN4018 : _GEN3243;
wire  _GEN4020 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4021 = io_x[10] ? _GEN4020 : _GEN3178;
wire  _GEN4022 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4023 = io_x[14] ? _GEN3175 : _GEN4022;
wire  _GEN4024 = io_x[10] ? _GEN4023 : _GEN3183;
wire  _GEN4025 = io_x[24] ? _GEN4024 : _GEN4021;
wire  _GEN4026 = io_x[17] ? _GEN4025 : _GEN3174;
wire  _GEN4027 = io_x[12] ? _GEN4026 : _GEN4019;
wire  _GEN4028 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4029 = io_x[10] ? _GEN3178 : _GEN4028;
wire  _GEN4030 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4031 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4032 = io_x[10] ? _GEN4031 : _GEN4030;
wire  _GEN4033 = io_x[24] ? _GEN4032 : _GEN4029;
wire  _GEN4034 = io_x[17] ? _GEN4033 : _GEN3174;
wire  _GEN4035 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4036 = io_x[14] ? _GEN4035 : _GEN3176;
wire  _GEN4037 = io_x[10] ? _GEN4036 : _GEN3178;
wire  _GEN4038 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4039 = io_x[14] ? _GEN3176 : _GEN4038;
wire  _GEN4040 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4041 = io_x[14] ? _GEN4040 : _GEN3176;
wire  _GEN4042 = io_x[10] ? _GEN4041 : _GEN4039;
wire  _GEN4043 = io_x[24] ? _GEN4042 : _GEN4037;
wire  _GEN4044 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4045 = io_x[14] ? _GEN4044 : _GEN3176;
wire  _GEN4046 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4047 = io_x[14] ? _GEN4046 : _GEN3175;
wire  _GEN4048 = io_x[10] ? _GEN4047 : _GEN4045;
wire  _GEN4049 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4050 = io_x[14] ? _GEN4049 : _GEN3176;
wire  _GEN4051 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4052 = io_x[14] ? _GEN4051 : _GEN3176;
wire  _GEN4053 = io_x[10] ? _GEN4052 : _GEN4050;
wire  _GEN4054 = io_x[24] ? _GEN4053 : _GEN4048;
wire  _GEN4055 = io_x[17] ? _GEN4054 : _GEN4043;
wire  _GEN4056 = io_x[12] ? _GEN4055 : _GEN4034;
wire  _GEN4057 = io_x[2] ? _GEN4056 : _GEN4027;
wire  _GEN4058 = io_x[9] ? _GEN4057 : _GEN4014;
wire  _GEN4059 = io_x[13] ? _GEN4058 : _GEN3976;
wire  _GEN4060 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN4061 = io_x[24] ? _GEN4060 : _GEN3180;
wire  _GEN4062 = io_x[17] ? _GEN4061 : _GEN3174;
wire  _GEN4063 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN4064 = io_x[24] ? _GEN3196 : _GEN4063;
wire  _GEN4065 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4066 = io_x[14] ? _GEN4065 : _GEN3176;
wire  _GEN4067 = io_x[10] ? _GEN4066 : _GEN3178;
wire  _GEN4068 = io_x[24] ? _GEN3180 : _GEN4067;
wire  _GEN4069 = io_x[17] ? _GEN4068 : _GEN4064;
wire  _GEN4070 = io_x[12] ? _GEN4069 : _GEN4062;
wire  _GEN4071 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4072 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4073 = io_x[14] ? _GEN4072 : _GEN3176;
wire  _GEN4074 = io_x[10] ? _GEN3183 : _GEN4073;
wire  _GEN4075 = io_x[24] ? _GEN4074 : _GEN4071;
wire  _GEN4076 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4077 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4078 = io_x[14] ? _GEN4077 : _GEN3176;
wire  _GEN4079 = io_x[10] ? _GEN4078 : _GEN4076;
wire  _GEN4080 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4081 = io_x[14] ? _GEN4080 : _GEN3176;
wire  _GEN4082 = io_x[10] ? _GEN4081 : _GEN3178;
wire  _GEN4083 = io_x[24] ? _GEN4082 : _GEN4079;
wire  _GEN4084 = io_x[17] ? _GEN4083 : _GEN4075;
wire  _GEN4085 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4086 = io_x[10] ? _GEN4085 : _GEN3183;
wire  _GEN4087 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4088 = io_x[14] ? _GEN4087 : _GEN3176;
wire  _GEN4089 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4090 = io_x[14] ? _GEN4089 : _GEN3176;
wire  _GEN4091 = io_x[10] ? _GEN4090 : _GEN4088;
wire  _GEN4092 = io_x[24] ? _GEN4091 : _GEN4086;
wire  _GEN4093 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4094 = io_x[14] ? _GEN3176 : _GEN4093;
wire  _GEN4095 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4096 = io_x[14] ? _GEN4095 : _GEN3176;
wire  _GEN4097 = io_x[10] ? _GEN4096 : _GEN4094;
wire  _GEN4098 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4099 = io_x[14] ? _GEN3175 : _GEN4098;
wire  _GEN4100 = io_x[10] ? _GEN4099 : _GEN3178;
wire  _GEN4101 = io_x[24] ? _GEN4100 : _GEN4097;
wire  _GEN4102 = io_x[17] ? _GEN4101 : _GEN4092;
wire  _GEN4103 = io_x[12] ? _GEN4102 : _GEN4084;
wire  _GEN4104 = io_x[2] ? _GEN4103 : _GEN4070;
wire  _GEN4105 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4106 = io_x[14] ? _GEN3176 : _GEN4105;
wire  _GEN4107 = io_x[10] ? _GEN3178 : _GEN4106;
wire  _GEN4108 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4109 = io_x[14] ? _GEN4108 : _GEN3176;
wire  _GEN4110 = io_x[10] ? _GEN3178 : _GEN4109;
wire  _GEN4111 = io_x[24] ? _GEN4110 : _GEN4107;
wire  _GEN4112 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4113 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4114 = io_x[14] ? _GEN4113 : _GEN3176;
wire  _GEN4115 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4116 = io_x[14] ? _GEN4115 : _GEN3176;
wire  _GEN4117 = io_x[10] ? _GEN4116 : _GEN4114;
wire  _GEN4118 = io_x[24] ? _GEN4117 : _GEN4112;
wire  _GEN4119 = io_x[17] ? _GEN4118 : _GEN4111;
wire  _GEN4120 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4121 = io_x[14] ? _GEN4120 : _GEN3175;
wire  _GEN4122 = io_x[10] ? _GEN4121 : _GEN3183;
wire  _GEN4123 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4124 = io_x[10] ? _GEN4123 : _GEN3183;
wire  _GEN4125 = io_x[24] ? _GEN4124 : _GEN4122;
wire  _GEN4126 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4127 = io_x[14] ? _GEN4126 : _GEN3175;
wire  _GEN4128 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4129 = io_x[14] ? _GEN4128 : _GEN3175;
wire  _GEN4130 = io_x[10] ? _GEN4129 : _GEN4127;
wire  _GEN4131 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4132 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4133 = io_x[10] ? _GEN4132 : _GEN4131;
wire  _GEN4134 = io_x[24] ? _GEN4133 : _GEN4130;
wire  _GEN4135 = io_x[17] ? _GEN4134 : _GEN4125;
wire  _GEN4136 = io_x[12] ? _GEN4135 : _GEN4119;
wire  _GEN4137 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4138 = io_x[14] ? _GEN4137 : _GEN3176;
wire  _GEN4139 = io_x[10] ? _GEN4138 : _GEN3178;
wire  _GEN4140 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4141 = io_x[14] ? _GEN4140 : _GEN3176;
wire  _GEN4142 = io_x[10] ? _GEN4141 : _GEN3178;
wire  _GEN4143 = io_x[24] ? _GEN4142 : _GEN4139;
wire  _GEN4144 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4145 = io_x[10] ? _GEN4144 : _GEN3178;
wire  _GEN4146 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4147 = io_x[14] ? _GEN4146 : _GEN3175;
wire  _GEN4148 = io_x[10] ? _GEN3183 : _GEN4147;
wire  _GEN4149 = io_x[24] ? _GEN4148 : _GEN4145;
wire  _GEN4150 = io_x[17] ? _GEN4149 : _GEN4143;
wire  _GEN4151 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4152 = io_x[14] ? _GEN4151 : _GEN3176;
wire  _GEN4153 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4154 = io_x[10] ? _GEN4153 : _GEN4152;
wire  _GEN4155 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4156 = io_x[14] ? _GEN3175 : _GEN4155;
wire  _GEN4157 = io_x[10] ? _GEN4156 : _GEN3178;
wire  _GEN4158 = io_x[24] ? _GEN4157 : _GEN4154;
wire  _GEN4159 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4160 = io_x[14] ? _GEN4159 : _GEN3175;
wire  _GEN4161 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4162 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4163 = io_x[14] ? _GEN4162 : _GEN4161;
wire  _GEN4164 = io_x[10] ? _GEN4163 : _GEN4160;
wire  _GEN4165 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4166 = io_x[14] ? _GEN3175 : _GEN4165;
wire  _GEN4167 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4168 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4169 = io_x[14] ? _GEN4168 : _GEN4167;
wire  _GEN4170 = io_x[10] ? _GEN4169 : _GEN4166;
wire  _GEN4171 = io_x[24] ? _GEN4170 : _GEN4164;
wire  _GEN4172 = io_x[17] ? _GEN4171 : _GEN4158;
wire  _GEN4173 = io_x[12] ? _GEN4172 : _GEN4150;
wire  _GEN4174 = io_x[2] ? _GEN4173 : _GEN4136;
wire  _GEN4175 = io_x[9] ? _GEN4174 : _GEN4104;
wire  _GEN4176 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4177 = io_x[14] ? _GEN3175 : _GEN4176;
wire  _GEN4178 = io_x[10] ? _GEN4177 : _GEN3178;
wire  _GEN4179 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4180 = io_x[10] ? _GEN3178 : _GEN4179;
wire  _GEN4181 = io_x[24] ? _GEN4180 : _GEN4178;
wire  _GEN4182 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4183 = io_x[14] ? _GEN4182 : _GEN3176;
wire  _GEN4184 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4185 = io_x[14] ? _GEN3176 : _GEN4184;
wire  _GEN4186 = io_x[10] ? _GEN4185 : _GEN4183;
wire  _GEN4187 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4188 = io_x[10] ? _GEN4187 : _GEN3183;
wire  _GEN4189 = io_x[24] ? _GEN4188 : _GEN4186;
wire  _GEN4190 = io_x[17] ? _GEN4189 : _GEN4181;
wire  _GEN4191 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4192 = io_x[10] ? _GEN4191 : _GEN3178;
wire  _GEN4193 = io_x[24] ? _GEN3180 : _GEN4192;
wire  _GEN4194 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4195 = io_x[14] ? _GEN4194 : _GEN3175;
wire  _GEN4196 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4197 = io_x[14] ? _GEN4196 : _GEN3176;
wire  _GEN4198 = io_x[10] ? _GEN4197 : _GEN4195;
wire  _GEN4199 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4200 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4201 = io_x[10] ? _GEN4200 : _GEN4199;
wire  _GEN4202 = io_x[24] ? _GEN4201 : _GEN4198;
wire  _GEN4203 = io_x[17] ? _GEN4202 : _GEN4193;
wire  _GEN4204 = io_x[12] ? _GEN4203 : _GEN4190;
wire  _GEN4205 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4206 = io_x[10] ? _GEN3178 : _GEN4205;
wire  _GEN4207 = io_x[24] ? _GEN4206 : _GEN3196;
wire  _GEN4208 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4209 = io_x[14] ? _GEN4208 : _GEN3176;
wire  _GEN4210 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4211 = io_x[10] ? _GEN4210 : _GEN4209;
wire  _GEN4212 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4213 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4214 = io_x[10] ? _GEN4213 : _GEN4212;
wire  _GEN4215 = io_x[24] ? _GEN4214 : _GEN4211;
wire  _GEN4216 = io_x[17] ? _GEN4215 : _GEN4207;
wire  _GEN4217 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4218 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4219 = io_x[14] ? _GEN4218 : _GEN4217;
wire  _GEN4220 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4221 = io_x[10] ? _GEN4220 : _GEN4219;
wire  _GEN4222 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4223 = io_x[24] ? _GEN4222 : _GEN4221;
wire  _GEN4224 = io_x[17] ? _GEN4223 : _GEN3243;
wire  _GEN4225 = io_x[12] ? _GEN4224 : _GEN4216;
wire  _GEN4226 = io_x[2] ? _GEN4225 : _GEN4204;
wire  _GEN4227 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4228 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4229 = io_x[14] ? _GEN4228 : _GEN4227;
wire  _GEN4230 = io_x[10] ? _GEN3178 : _GEN4229;
wire  _GEN4231 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4232 = io_x[14] ? _GEN4231 : _GEN3176;
wire  _GEN4233 = io_x[10] ? _GEN4232 : _GEN3183;
wire  _GEN4234 = io_x[24] ? _GEN4233 : _GEN4230;
wire  _GEN4235 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4236 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4237 = io_x[14] ? _GEN4236 : _GEN4235;
wire  _GEN4238 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4239 = io_x[14] ? _GEN4238 : _GEN3176;
wire  _GEN4240 = io_x[10] ? _GEN4239 : _GEN4237;
wire  _GEN4241 = io_x[24] ? _GEN3196 : _GEN4240;
wire  _GEN4242 = io_x[17] ? _GEN4241 : _GEN4234;
wire  _GEN4243 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4244 = io_x[14] ? _GEN4243 : _GEN3176;
wire  _GEN4245 = io_x[10] ? _GEN4244 : _GEN3183;
wire  _GEN4246 = io_x[24] ? _GEN3180 : _GEN4245;
wire  _GEN4247 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4248 = io_x[14] ? _GEN4247 : _GEN3175;
wire  _GEN4249 = io_x[10] ? _GEN4248 : _GEN3183;
wire  _GEN4250 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4251 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4252 = io_x[14] ? _GEN4251 : _GEN4250;
wire  _GEN4253 = io_x[10] ? _GEN4252 : _GEN3178;
wire  _GEN4254 = io_x[24] ? _GEN4253 : _GEN4249;
wire  _GEN4255 = io_x[17] ? _GEN4254 : _GEN4246;
wire  _GEN4256 = io_x[12] ? _GEN4255 : _GEN4242;
wire  _GEN4257 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4258 = io_x[10] ? _GEN4257 : _GEN3178;
wire  _GEN4259 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4260 = io_x[14] ? _GEN3176 : _GEN4259;
wire  _GEN4261 = io_x[10] ? _GEN3178 : _GEN4260;
wire  _GEN4262 = io_x[24] ? _GEN4261 : _GEN4258;
wire  _GEN4263 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4264 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4265 = io_x[10] ? _GEN4264 : _GEN4263;
wire  _GEN4266 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4267 = io_x[10] ? _GEN4266 : _GEN3178;
wire  _GEN4268 = io_x[24] ? _GEN4267 : _GEN4265;
wire  _GEN4269 = io_x[17] ? _GEN4268 : _GEN4262;
wire  _GEN4270 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4271 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4272 = io_x[14] ? _GEN4271 : _GEN3176;
wire  _GEN4273 = io_x[10] ? _GEN4272 : _GEN4270;
wire  _GEN4274 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4275 = io_x[14] ? _GEN4274 : _GEN3175;
wire  _GEN4276 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4277 = io_x[14] ? _GEN4276 : _GEN3176;
wire  _GEN4278 = io_x[10] ? _GEN4277 : _GEN4275;
wire  _GEN4279 = io_x[24] ? _GEN4278 : _GEN4273;
wire  _GEN4280 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4281 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4282 = io_x[14] ? _GEN4281 : _GEN4280;
wire  _GEN4283 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4284 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4285 = io_x[14] ? _GEN4284 : _GEN4283;
wire  _GEN4286 = io_x[10] ? _GEN4285 : _GEN4282;
wire  _GEN4287 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4288 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4289 = io_x[14] ? _GEN4288 : _GEN4287;
wire  _GEN4290 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4291 = io_x[14] ? _GEN4290 : _GEN3176;
wire  _GEN4292 = io_x[10] ? _GEN4291 : _GEN4289;
wire  _GEN4293 = io_x[24] ? _GEN4292 : _GEN4286;
wire  _GEN4294 = io_x[17] ? _GEN4293 : _GEN4279;
wire  _GEN4295 = io_x[12] ? _GEN4294 : _GEN4269;
wire  _GEN4296 = io_x[2] ? _GEN4295 : _GEN4256;
wire  _GEN4297 = io_x[9] ? _GEN4296 : _GEN4226;
wire  _GEN4298 = io_x[13] ? _GEN4297 : _GEN4175;
wire  _GEN4299 = io_x[7] ? _GEN4298 : _GEN4059;
wire  _GEN4300 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4301 = io_x[10] ? _GEN4300 : _GEN3178;
wire  _GEN4302 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4303 = io_x[10] ? _GEN3178 : _GEN4302;
wire  _GEN4304 = io_x[24] ? _GEN4303 : _GEN4301;
wire  _GEN4305 = io_x[17] ? _GEN4304 : _GEN3174;
wire  _GEN4306 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4307 = io_x[10] ? _GEN4306 : _GEN3178;
wire  _GEN4308 = io_x[24] ? _GEN3180 : _GEN4307;
wire  _GEN4309 = io_x[17] ? _GEN4308 : _GEN3174;
wire  _GEN4310 = io_x[12] ? _GEN4309 : _GEN4305;
wire  _GEN4311 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4312 = io_x[10] ? _GEN4311 : _GEN3178;
wire  _GEN4313 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4314 = io_x[14] ? _GEN4313 : _GEN3176;
wire  _GEN4315 = io_x[10] ? _GEN3178 : _GEN4314;
wire  _GEN4316 = io_x[24] ? _GEN4315 : _GEN4312;
wire  _GEN4317 = io_x[17] ? _GEN4316 : _GEN3243;
wire  _GEN4318 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4319 = io_x[14] ? _GEN4318 : _GEN3176;
wire  _GEN4320 = io_x[10] ? _GEN4319 : _GEN3183;
wire  _GEN4321 = io_x[24] ? _GEN4320 : _GEN3196;
wire  _GEN4322 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4323 = io_x[14] ? _GEN3176 : _GEN4322;
wire  _GEN4324 = io_x[10] ? _GEN3183 : _GEN4323;
wire  _GEN4325 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4326 = io_x[14] ? _GEN4325 : _GEN3175;
wire  _GEN4327 = io_x[10] ? _GEN4326 : _GEN3178;
wire  _GEN4328 = io_x[24] ? _GEN4327 : _GEN4324;
wire  _GEN4329 = io_x[17] ? _GEN4328 : _GEN4321;
wire  _GEN4330 = io_x[12] ? _GEN4329 : _GEN4317;
wire  _GEN4331 = io_x[2] ? _GEN4330 : _GEN4310;
wire  _GEN4332 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4333 = io_x[10] ? _GEN3178 : _GEN4332;
wire  _GEN4334 = io_x[24] ? _GEN3180 : _GEN4333;
wire  _GEN4335 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4336 = io_x[14] ? _GEN4335 : _GEN3176;
wire  _GEN4337 = io_x[10] ? _GEN3178 : _GEN4336;
wire  _GEN4338 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4339 = io_x[10] ? _GEN3183 : _GEN4338;
wire  _GEN4340 = io_x[24] ? _GEN4339 : _GEN4337;
wire  _GEN4341 = io_x[17] ? _GEN4340 : _GEN4334;
wire  _GEN4342 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4343 = io_x[10] ? _GEN3178 : _GEN4342;
wire  _GEN4344 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4345 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4346 = io_x[14] ? _GEN4345 : _GEN3176;
wire  _GEN4347 = io_x[10] ? _GEN4346 : _GEN4344;
wire  _GEN4348 = io_x[24] ? _GEN4347 : _GEN4343;
wire  _GEN4349 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4350 = io_x[14] ? _GEN4349 : _GEN3176;
wire  _GEN4351 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4352 = io_x[14] ? _GEN4351 : _GEN3175;
wire  _GEN4353 = io_x[10] ? _GEN4352 : _GEN4350;
wire  _GEN4354 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4355 = io_x[14] ? _GEN3175 : _GEN4354;
wire  _GEN4356 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4357 = io_x[14] ? _GEN4356 : _GEN3176;
wire  _GEN4358 = io_x[10] ? _GEN4357 : _GEN4355;
wire  _GEN4359 = io_x[24] ? _GEN4358 : _GEN4353;
wire  _GEN4360 = io_x[17] ? _GEN4359 : _GEN4348;
wire  _GEN4361 = io_x[12] ? _GEN4360 : _GEN4341;
wire  _GEN4362 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN4363 = io_x[24] ? _GEN3180 : _GEN4362;
wire  _GEN4364 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4365 = io_x[10] ? _GEN3183 : _GEN4364;
wire  _GEN4366 = io_x[24] ? _GEN4365 : _GEN3180;
wire  _GEN4367 = io_x[17] ? _GEN4366 : _GEN4363;
wire  _GEN4368 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4369 = io_x[14] ? _GEN3176 : _GEN4368;
wire  _GEN4370 = io_x[10] ? _GEN3183 : _GEN4369;
wire  _GEN4371 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4372 = io_x[14] ? _GEN4371 : _GEN3176;
wire  _GEN4373 = io_x[10] ? _GEN4372 : _GEN3178;
wire  _GEN4374 = io_x[24] ? _GEN4373 : _GEN4370;
wire  _GEN4375 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4376 = io_x[10] ? _GEN4375 : _GEN3178;
wire  _GEN4377 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4378 = io_x[14] ? _GEN3176 : _GEN4377;
wire  _GEN4379 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4380 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4381 = io_x[14] ? _GEN4380 : _GEN4379;
wire  _GEN4382 = io_x[10] ? _GEN4381 : _GEN4378;
wire  _GEN4383 = io_x[24] ? _GEN4382 : _GEN4376;
wire  _GEN4384 = io_x[17] ? _GEN4383 : _GEN4374;
wire  _GEN4385 = io_x[12] ? _GEN4384 : _GEN4367;
wire  _GEN4386 = io_x[2] ? _GEN4385 : _GEN4361;
wire  _GEN4387 = io_x[9] ? _GEN4386 : _GEN4331;
wire  _GEN4388 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4389 = io_x[14] ? _GEN4388 : _GEN3175;
wire  _GEN4390 = io_x[10] ? _GEN4389 : _GEN3178;
wire  _GEN4391 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4392 = io_x[14] ? _GEN3176 : _GEN4391;
wire  _GEN4393 = io_x[10] ? _GEN4392 : _GEN3178;
wire  _GEN4394 = io_x[24] ? _GEN4393 : _GEN4390;
wire  _GEN4395 = io_x[17] ? _GEN4394 : _GEN3174;
wire  _GEN4396 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4397 = io_x[24] ? _GEN3180 : _GEN4396;
wire  _GEN4398 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4399 = io_x[14] ? _GEN4398 : _GEN3175;
wire  _GEN4400 = io_x[10] ? _GEN4399 : _GEN3183;
wire  _GEN4401 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4402 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4403 = io_x[14] ? _GEN4402 : _GEN4401;
wire  _GEN4404 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4405 = io_x[10] ? _GEN4404 : _GEN4403;
wire  _GEN4406 = io_x[24] ? _GEN4405 : _GEN4400;
wire  _GEN4407 = io_x[17] ? _GEN4406 : _GEN4397;
wire  _GEN4408 = io_x[12] ? _GEN4407 : _GEN4395;
wire  _GEN4409 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4410 = io_x[10] ? _GEN4409 : _GEN3178;
wire  _GEN4411 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4412 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4413 = io_x[14] ? _GEN3175 : _GEN4412;
wire  _GEN4414 = io_x[10] ? _GEN4413 : _GEN4411;
wire  _GEN4415 = io_x[24] ? _GEN4414 : _GEN4410;
wire  _GEN4416 = io_x[17] ? _GEN4415 : _GEN3174;
wire  _GEN4417 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4418 = io_x[14] ? _GEN4417 : _GEN3176;
wire  _GEN4419 = io_x[10] ? _GEN4418 : _GEN3183;
wire  _GEN4420 = io_x[24] ? _GEN4419 : _GEN3180;
wire  _GEN4421 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4422 = io_x[14] ? _GEN4421 : _GEN3176;
wire  _GEN4423 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4424 = io_x[14] ? _GEN4423 : _GEN3176;
wire  _GEN4425 = io_x[10] ? _GEN4424 : _GEN4422;
wire  _GEN4426 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4427 = io_x[14] ? _GEN4426 : _GEN3176;
wire  _GEN4428 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4429 = io_x[14] ? _GEN3175 : _GEN4428;
wire  _GEN4430 = io_x[10] ? _GEN4429 : _GEN4427;
wire  _GEN4431 = io_x[24] ? _GEN4430 : _GEN4425;
wire  _GEN4432 = io_x[17] ? _GEN4431 : _GEN4420;
wire  _GEN4433 = io_x[12] ? _GEN4432 : _GEN4416;
wire  _GEN4434 = io_x[2] ? _GEN4433 : _GEN4408;
wire  _GEN4435 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4436 = io_x[14] ? _GEN4435 : _GEN3176;
wire  _GEN4437 = io_x[10] ? _GEN4436 : _GEN3183;
wire  _GEN4438 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4439 = io_x[10] ? _GEN3178 : _GEN4438;
wire  _GEN4440 = io_x[24] ? _GEN4439 : _GEN4437;
wire  _GEN4441 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4442 = io_x[14] ? _GEN3176 : _GEN4441;
wire  _GEN4443 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4444 = io_x[14] ? _GEN4443 : _GEN3176;
wire  _GEN4445 = io_x[10] ? _GEN4444 : _GEN4442;
wire  _GEN4446 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4447 = io_x[14] ? _GEN3176 : _GEN4446;
wire  _GEN4448 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4449 = io_x[10] ? _GEN4448 : _GEN4447;
wire  _GEN4450 = io_x[24] ? _GEN4449 : _GEN4445;
wire  _GEN4451 = io_x[17] ? _GEN4450 : _GEN4440;
wire  _GEN4452 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4453 = io_x[14] ? _GEN4452 : _GEN3176;
wire  _GEN4454 = io_x[10] ? _GEN4453 : _GEN3178;
wire  _GEN4455 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4456 = io_x[14] ? _GEN3176 : _GEN4455;
wire  _GEN4457 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4458 = io_x[10] ? _GEN4457 : _GEN4456;
wire  _GEN4459 = io_x[24] ? _GEN4458 : _GEN4454;
wire  _GEN4460 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4461 = io_x[14] ? _GEN4460 : _GEN3176;
wire  _GEN4462 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4463 = io_x[14] ? _GEN4462 : _GEN3175;
wire  _GEN4464 = io_x[10] ? _GEN4463 : _GEN4461;
wire  _GEN4465 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4466 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4467 = io_x[14] ? _GEN4466 : _GEN4465;
wire  _GEN4468 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4469 = io_x[14] ? _GEN4468 : _GEN3175;
wire  _GEN4470 = io_x[10] ? _GEN4469 : _GEN4467;
wire  _GEN4471 = io_x[24] ? _GEN4470 : _GEN4464;
wire  _GEN4472 = io_x[17] ? _GEN4471 : _GEN4459;
wire  _GEN4473 = io_x[12] ? _GEN4472 : _GEN4451;
wire  _GEN4474 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4475 = io_x[14] ? _GEN3176 : _GEN4474;
wire  _GEN4476 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4477 = io_x[14] ? _GEN4476 : _GEN3176;
wire  _GEN4478 = io_x[10] ? _GEN4477 : _GEN4475;
wire  _GEN4479 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4480 = io_x[14] ? _GEN4479 : _GEN3175;
wire  _GEN4481 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4482 = io_x[14] ? _GEN4481 : _GEN3176;
wire  _GEN4483 = io_x[10] ? _GEN4482 : _GEN4480;
wire  _GEN4484 = io_x[24] ? _GEN4483 : _GEN4478;
wire  _GEN4485 = io_x[17] ? _GEN4484 : _GEN3243;
wire  _GEN4486 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4487 = io_x[14] ? _GEN4486 : _GEN3176;
wire  _GEN4488 = io_x[10] ? _GEN4487 : _GEN3183;
wire  _GEN4489 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4490 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4491 = io_x[14] ? _GEN4490 : _GEN3176;
wire  _GEN4492 = io_x[10] ? _GEN4491 : _GEN4489;
wire  _GEN4493 = io_x[24] ? _GEN4492 : _GEN4488;
wire  _GEN4494 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4495 = io_x[14] ? _GEN4494 : _GEN3175;
wire  _GEN4496 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4497 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4498 = io_x[14] ? _GEN4497 : _GEN4496;
wire  _GEN4499 = io_x[10] ? _GEN4498 : _GEN4495;
wire  _GEN4500 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4501 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4502 = io_x[14] ? _GEN4501 : _GEN4500;
wire  _GEN4503 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4504 = io_x[14] ? _GEN4503 : _GEN3176;
wire  _GEN4505 = io_x[10] ? _GEN4504 : _GEN4502;
wire  _GEN4506 = io_x[24] ? _GEN4505 : _GEN4499;
wire  _GEN4507 = io_x[17] ? _GEN4506 : _GEN4493;
wire  _GEN4508 = io_x[12] ? _GEN4507 : _GEN4485;
wire  _GEN4509 = io_x[2] ? _GEN4508 : _GEN4473;
wire  _GEN4510 = io_x[9] ? _GEN4509 : _GEN4434;
wire  _GEN4511 = io_x[13] ? _GEN4510 : _GEN4387;
wire  _GEN4512 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4513 = io_x[14] ? _GEN3176 : _GEN4512;
wire  _GEN4514 = io_x[10] ? _GEN3183 : _GEN4513;
wire  _GEN4515 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4516 = io_x[14] ? _GEN4515 : _GEN3176;
wire  _GEN4517 = io_x[10] ? _GEN4516 : _GEN3178;
wire  _GEN4518 = io_x[24] ? _GEN4517 : _GEN4514;
wire  _GEN4519 = io_x[17] ? _GEN4518 : _GEN3243;
wire  _GEN4520 = io_x[24] ? _GEN3180 : _GEN3196;
wire  _GEN4521 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4522 = io_x[14] ? _GEN4521 : _GEN3176;
wire  _GEN4523 = io_x[10] ? _GEN4522 : _GEN3183;
wire  _GEN4524 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4525 = io_x[14] ? _GEN3176 : _GEN4524;
wire  _GEN4526 = io_x[10] ? _GEN4525 : _GEN3183;
wire  _GEN4527 = io_x[24] ? _GEN4526 : _GEN4523;
wire  _GEN4528 = io_x[17] ? _GEN4527 : _GEN4520;
wire  _GEN4529 = io_x[12] ? _GEN4528 : _GEN4519;
wire  _GEN4530 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4531 = io_x[10] ? _GEN4530 : _GEN3183;
wire  _GEN4532 = io_x[24] ? _GEN4531 : _GEN3180;
wire  _GEN4533 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4534 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4535 = io_x[14] ? _GEN4534 : _GEN4533;
wire  _GEN4536 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4537 = io_x[10] ? _GEN4536 : _GEN4535;
wire  _GEN4538 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4539 = io_x[10] ? _GEN4538 : _GEN3183;
wire  _GEN4540 = io_x[24] ? _GEN4539 : _GEN4537;
wire  _GEN4541 = io_x[17] ? _GEN4540 : _GEN4532;
wire  _GEN4542 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4543 = io_x[14] ? _GEN4542 : _GEN3176;
wire  _GEN4544 = io_x[10] ? _GEN4543 : _GEN3183;
wire  _GEN4545 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4546 = io_x[10] ? _GEN4545 : _GEN3183;
wire  _GEN4547 = io_x[24] ? _GEN4546 : _GEN4544;
wire  _GEN4548 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4549 = io_x[14] ? _GEN4548 : _GEN3175;
wire  _GEN4550 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4551 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4552 = io_x[14] ? _GEN4551 : _GEN4550;
wire  _GEN4553 = io_x[10] ? _GEN4552 : _GEN4549;
wire  _GEN4554 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4555 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4556 = io_x[14] ? _GEN4555 : _GEN4554;
wire  _GEN4557 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4558 = io_x[10] ? _GEN4557 : _GEN4556;
wire  _GEN4559 = io_x[24] ? _GEN4558 : _GEN4553;
wire  _GEN4560 = io_x[17] ? _GEN4559 : _GEN4547;
wire  _GEN4561 = io_x[12] ? _GEN4560 : _GEN4541;
wire  _GEN4562 = io_x[2] ? _GEN4561 : _GEN4529;
wire  _GEN4563 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4564 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4565 = io_x[14] ? _GEN4564 : _GEN4563;
wire  _GEN4566 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4567 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4568 = io_x[14] ? _GEN4567 : _GEN4566;
wire  _GEN4569 = io_x[10] ? _GEN4568 : _GEN4565;
wire  _GEN4570 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4571 = io_x[14] ? _GEN4570 : _GEN3176;
wire  _GEN4572 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4573 = io_x[10] ? _GEN4572 : _GEN4571;
wire  _GEN4574 = io_x[24] ? _GEN4573 : _GEN4569;
wire  _GEN4575 = io_x[17] ? _GEN4574 : _GEN3243;
wire  _GEN4576 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4577 = io_x[14] ? _GEN3176 : _GEN4576;
wire  _GEN4578 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4579 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4580 = io_x[14] ? _GEN4579 : _GEN4578;
wire  _GEN4581 = io_x[10] ? _GEN4580 : _GEN4577;
wire  _GEN4582 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4583 = io_x[10] ? _GEN4582 : _GEN3178;
wire  _GEN4584 = io_x[24] ? _GEN4583 : _GEN4581;
wire  _GEN4585 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4586 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4587 = io_x[14] ? _GEN4586 : _GEN4585;
wire  _GEN4588 = io_x[10] ? _GEN4587 : _GEN3183;
wire  _GEN4589 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN4590 = io_x[24] ? _GEN4589 : _GEN4588;
wire  _GEN4591 = io_x[17] ? _GEN4590 : _GEN4584;
wire  _GEN4592 = io_x[12] ? _GEN4591 : _GEN4575;
wire  _GEN4593 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4594 = io_x[14] ? _GEN4593 : _GEN3176;
wire  _GEN4595 = io_x[10] ? _GEN4594 : _GEN3183;
wire  _GEN4596 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4597 = io_x[14] ? _GEN4596 : _GEN3176;
wire  _GEN4598 = io_x[10] ? _GEN4597 : _GEN3178;
wire  _GEN4599 = io_x[24] ? _GEN4598 : _GEN4595;
wire  _GEN4600 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4601 = io_x[14] ? _GEN4600 : _GEN3176;
wire  _GEN4602 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4603 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4604 = io_x[14] ? _GEN4603 : _GEN4602;
wire  _GEN4605 = io_x[10] ? _GEN4604 : _GEN4601;
wire  _GEN4606 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4607 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4608 = io_x[14] ? _GEN3175 : _GEN4607;
wire  _GEN4609 = io_x[10] ? _GEN4608 : _GEN4606;
wire  _GEN4610 = io_x[24] ? _GEN4609 : _GEN4605;
wire  _GEN4611 = io_x[17] ? _GEN4610 : _GEN4599;
wire  _GEN4612 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4613 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4614 = io_x[14] ? _GEN4613 : _GEN4612;
wire  _GEN4615 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4616 = io_x[14] ? _GEN4615 : _GEN3176;
wire  _GEN4617 = io_x[10] ? _GEN4616 : _GEN4614;
wire  _GEN4618 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4619 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4620 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4621 = io_x[14] ? _GEN4620 : _GEN4619;
wire  _GEN4622 = io_x[10] ? _GEN4621 : _GEN4618;
wire  _GEN4623 = io_x[24] ? _GEN4622 : _GEN4617;
wire  _GEN4624 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4625 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4626 = io_x[14] ? _GEN4625 : _GEN4624;
wire  _GEN4627 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4628 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4629 = io_x[14] ? _GEN4628 : _GEN4627;
wire  _GEN4630 = io_x[10] ? _GEN4629 : _GEN4626;
wire  _GEN4631 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4632 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4633 = io_x[14] ? _GEN4632 : _GEN4631;
wire  _GEN4634 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4635 = io_x[14] ? _GEN4634 : _GEN3176;
wire  _GEN4636 = io_x[10] ? _GEN4635 : _GEN4633;
wire  _GEN4637 = io_x[24] ? _GEN4636 : _GEN4630;
wire  _GEN4638 = io_x[17] ? _GEN4637 : _GEN4623;
wire  _GEN4639 = io_x[12] ? _GEN4638 : _GEN4611;
wire  _GEN4640 = io_x[2] ? _GEN4639 : _GEN4592;
wire  _GEN4641 = io_x[9] ? _GEN4640 : _GEN4562;
wire  _GEN4642 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4643 = io_x[14] ? _GEN3176 : _GEN4642;
wire  _GEN4644 = io_x[10] ? _GEN4643 : _GEN3178;
wire  _GEN4645 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4646 = io_x[24] ? _GEN4645 : _GEN4644;
wire  _GEN4647 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4648 = io_x[14] ? _GEN4647 : _GEN3175;
wire  _GEN4649 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4650 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4651 = io_x[14] ? _GEN4650 : _GEN4649;
wire  _GEN4652 = io_x[10] ? _GEN4651 : _GEN4648;
wire  _GEN4653 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4654 = io_x[14] ? _GEN4653 : _GEN3176;
wire  _GEN4655 = io_x[10] ? _GEN4654 : _GEN3183;
wire  _GEN4656 = io_x[24] ? _GEN4655 : _GEN4652;
wire  _GEN4657 = io_x[17] ? _GEN4656 : _GEN4646;
wire  _GEN4658 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4659 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4660 = io_x[14] ? _GEN4659 : _GEN4658;
wire  _GEN4661 = io_x[10] ? _GEN4660 : _GEN3178;
wire  _GEN4662 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4663 = io_x[14] ? _GEN4662 : _GEN3176;
wire  _GEN4664 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4665 = io_x[14] ? _GEN4664 : _GEN3175;
wire  _GEN4666 = io_x[10] ? _GEN4665 : _GEN4663;
wire  _GEN4667 = io_x[24] ? _GEN4666 : _GEN4661;
wire  _GEN4668 = io_x[17] ? _GEN4667 : _GEN3174;
wire  _GEN4669 = io_x[12] ? _GEN4668 : _GEN4657;
wire  _GEN4670 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4671 = io_x[14] ? _GEN3175 : _GEN4670;
wire  _GEN4672 = io_x[10] ? _GEN4671 : _GEN3178;
wire  _GEN4673 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4674 = io_x[14] ? _GEN3176 : _GEN4673;
wire  _GEN4675 = io_x[10] ? _GEN4674 : _GEN3183;
wire  _GEN4676 = io_x[24] ? _GEN4675 : _GEN4672;
wire  _GEN4677 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4678 = io_x[14] ? _GEN4677 : _GEN3175;
wire  _GEN4679 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4680 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4681 = io_x[14] ? _GEN4680 : _GEN4679;
wire  _GEN4682 = io_x[10] ? _GEN4681 : _GEN4678;
wire  _GEN4683 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4684 = io_x[10] ? _GEN3183 : _GEN4683;
wire  _GEN4685 = io_x[24] ? _GEN4684 : _GEN4682;
wire  _GEN4686 = io_x[17] ? _GEN4685 : _GEN4676;
wire  _GEN4687 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4688 = io_x[14] ? _GEN4687 : _GEN3175;
wire  _GEN4689 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4690 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4691 = io_x[14] ? _GEN4690 : _GEN4689;
wire  _GEN4692 = io_x[10] ? _GEN4691 : _GEN4688;
wire  _GEN4693 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4694 = io_x[14] ? _GEN4693 : _GEN3176;
wire  _GEN4695 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4696 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4697 = io_x[14] ? _GEN4696 : _GEN4695;
wire  _GEN4698 = io_x[10] ? _GEN4697 : _GEN4694;
wire  _GEN4699 = io_x[24] ? _GEN4698 : _GEN4692;
wire  _GEN4700 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4701 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4702 = io_x[14] ? _GEN4701 : _GEN4700;
wire  _GEN4703 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4704 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4705 = io_x[14] ? _GEN4704 : _GEN4703;
wire  _GEN4706 = io_x[10] ? _GEN4705 : _GEN4702;
wire  _GEN4707 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4708 = io_x[14] ? _GEN4707 : _GEN3176;
wire  _GEN4709 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4710 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4711 = io_x[14] ? _GEN4710 : _GEN4709;
wire  _GEN4712 = io_x[10] ? _GEN4711 : _GEN4708;
wire  _GEN4713 = io_x[24] ? _GEN4712 : _GEN4706;
wire  _GEN4714 = io_x[17] ? _GEN4713 : _GEN4699;
wire  _GEN4715 = io_x[12] ? _GEN4714 : _GEN4686;
wire  _GEN4716 = io_x[2] ? _GEN4715 : _GEN4669;
wire  _GEN4717 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4718 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4719 = io_x[14] ? _GEN3175 : _GEN4718;
wire  _GEN4720 = io_x[10] ? _GEN4719 : _GEN4717;
wire  _GEN4721 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4722 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4723 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4724 = io_x[14] ? _GEN4723 : _GEN4722;
wire  _GEN4725 = io_x[10] ? _GEN4724 : _GEN4721;
wire  _GEN4726 = io_x[24] ? _GEN4725 : _GEN4720;
wire  _GEN4727 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4728 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4729 = io_x[14] ? _GEN4728 : _GEN4727;
wire  _GEN4730 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4731 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4732 = io_x[14] ? _GEN4731 : _GEN4730;
wire  _GEN4733 = io_x[10] ? _GEN4732 : _GEN4729;
wire  _GEN4734 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4735 = io_x[14] ? _GEN3176 : _GEN4734;
wire  _GEN4736 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4737 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4738 = io_x[14] ? _GEN4737 : _GEN4736;
wire  _GEN4739 = io_x[10] ? _GEN4738 : _GEN4735;
wire  _GEN4740 = io_x[24] ? _GEN4739 : _GEN4733;
wire  _GEN4741 = io_x[17] ? _GEN4740 : _GEN4726;
wire  _GEN4742 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4743 = io_x[14] ? _GEN4742 : _GEN3175;
wire  _GEN4744 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4745 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4746 = io_x[14] ? _GEN4745 : _GEN4744;
wire  _GEN4747 = io_x[10] ? _GEN4746 : _GEN4743;
wire  _GEN4748 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4749 = io_x[14] ? _GEN3176 : _GEN4748;
wire  _GEN4750 = io_x[10] ? _GEN4749 : _GEN3183;
wire  _GEN4751 = io_x[24] ? _GEN4750 : _GEN4747;
wire  _GEN4752 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4753 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4754 = io_x[14] ? _GEN4753 : _GEN4752;
wire  _GEN4755 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4756 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4757 = io_x[14] ? _GEN4756 : _GEN4755;
wire  _GEN4758 = io_x[10] ? _GEN4757 : _GEN4754;
wire  _GEN4759 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4760 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4761 = io_x[14] ? _GEN4760 : _GEN4759;
wire  _GEN4762 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4763 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4764 = io_x[14] ? _GEN4763 : _GEN4762;
wire  _GEN4765 = io_x[10] ? _GEN4764 : _GEN4761;
wire  _GEN4766 = io_x[24] ? _GEN4765 : _GEN4758;
wire  _GEN4767 = io_x[17] ? _GEN4766 : _GEN4751;
wire  _GEN4768 = io_x[12] ? _GEN4767 : _GEN4741;
wire  _GEN4769 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4770 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4771 = io_x[14] ? _GEN4770 : _GEN4769;
wire  _GEN4772 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4773 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4774 = io_x[14] ? _GEN4773 : _GEN4772;
wire  _GEN4775 = io_x[10] ? _GEN4774 : _GEN4771;
wire  _GEN4776 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4777 = io_x[14] ? _GEN3175 : _GEN4776;
wire  _GEN4778 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4779 = io_x[14] ? _GEN4778 : _GEN3176;
wire  _GEN4780 = io_x[10] ? _GEN4779 : _GEN4777;
wire  _GEN4781 = io_x[24] ? _GEN4780 : _GEN4775;
wire  _GEN4782 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4783 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4784 = io_x[14] ? _GEN4783 : _GEN4782;
wire  _GEN4785 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4786 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4787 = io_x[14] ? _GEN4786 : _GEN4785;
wire  _GEN4788 = io_x[10] ? _GEN4787 : _GEN4784;
wire  _GEN4789 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4790 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4791 = io_x[14] ? _GEN4790 : _GEN4789;
wire  _GEN4792 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4793 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4794 = io_x[14] ? _GEN4793 : _GEN4792;
wire  _GEN4795 = io_x[10] ? _GEN4794 : _GEN4791;
wire  _GEN4796 = io_x[24] ? _GEN4795 : _GEN4788;
wire  _GEN4797 = io_x[17] ? _GEN4796 : _GEN4781;
wire  _GEN4798 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4799 = io_x[14] ? _GEN4798 : _GEN3176;
wire  _GEN4800 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4801 = io_x[14] ? _GEN4800 : _GEN3176;
wire  _GEN4802 = io_x[10] ? _GEN4801 : _GEN4799;
wire  _GEN4803 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4804 = io_x[14] ? _GEN4803 : _GEN3176;
wire  _GEN4805 = io_x[10] ? _GEN4804 : _GEN3178;
wire  _GEN4806 = io_x[24] ? _GEN4805 : _GEN4802;
wire  _GEN4807 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4808 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4809 = io_x[14] ? _GEN4808 : _GEN4807;
wire  _GEN4810 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4811 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4812 = io_x[14] ? _GEN4811 : _GEN4810;
wire  _GEN4813 = io_x[10] ? _GEN4812 : _GEN4809;
wire  _GEN4814 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4815 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4816 = io_x[14] ? _GEN4815 : _GEN4814;
wire  _GEN4817 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4818 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4819 = io_x[14] ? _GEN4818 : _GEN4817;
wire  _GEN4820 = io_x[10] ? _GEN4819 : _GEN4816;
wire  _GEN4821 = io_x[24] ? _GEN4820 : _GEN4813;
wire  _GEN4822 = io_x[17] ? _GEN4821 : _GEN4806;
wire  _GEN4823 = io_x[12] ? _GEN4822 : _GEN4797;
wire  _GEN4824 = io_x[2] ? _GEN4823 : _GEN4768;
wire  _GEN4825 = io_x[9] ? _GEN4824 : _GEN4716;
wire  _GEN4826 = io_x[13] ? _GEN4825 : _GEN4641;
wire  _GEN4827 = io_x[7] ? _GEN4826 : _GEN4511;
wire  _GEN4828 = io_x[15] ? _GEN4827 : _GEN4299;
wire  _GEN4829 = io_x[3] ? _GEN4828 : _GEN3903;
wire  _GEN4830 = io_x[24] ? _GEN3180 : _GEN3196;
wire  _GEN4831 = io_x[17] ? _GEN4830 : _GEN3174;
wire  _GEN4832 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4833 = io_x[10] ? _GEN3183 : _GEN4832;
wire  _GEN4834 = io_x[24] ? _GEN4833 : _GEN3196;
wire  _GEN4835 = io_x[24] ? _GEN3180 : _GEN3196;
wire  _GEN4836 = io_x[17] ? _GEN4835 : _GEN4834;
wire  _GEN4837 = io_x[12] ? _GEN4836 : _GEN4831;
wire  _GEN4838 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN4839 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4840 = io_x[14] ? _GEN4839 : _GEN3176;
wire  _GEN4841 = io_x[10] ? _GEN4840 : _GEN3178;
wire  _GEN4842 = io_x[24] ? _GEN4841 : _GEN4838;
wire  _GEN4843 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4844 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4845 = io_x[14] ? _GEN4844 : _GEN3176;
wire  _GEN4846 = io_x[10] ? _GEN4845 : _GEN4843;
wire  _GEN4847 = io_x[24] ? _GEN4846 : _GEN3180;
wire  _GEN4848 = io_x[17] ? _GEN4847 : _GEN4842;
wire  _GEN4849 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4850 = io_x[14] ? _GEN4849 : _GEN3176;
wire  _GEN4851 = io_x[10] ? _GEN4850 : _GEN3183;
wire  _GEN4852 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4853 = io_x[24] ? _GEN4852 : _GEN4851;
wire  _GEN4854 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4855 = io_x[14] ? _GEN4854 : _GEN3176;
wire  _GEN4856 = io_x[10] ? _GEN4855 : _GEN3183;
wire  _GEN4857 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4858 = io_x[24] ? _GEN4857 : _GEN4856;
wire  _GEN4859 = io_x[17] ? _GEN4858 : _GEN4853;
wire  _GEN4860 = io_x[12] ? _GEN4859 : _GEN4848;
wire  _GEN4861 = io_x[2] ? _GEN4860 : _GEN4837;
wire  _GEN4862 = io_x[24] ? _GEN3196 : _GEN3180;
wire  _GEN4863 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4864 = io_x[14] ? _GEN4863 : _GEN3176;
wire  _GEN4865 = io_x[10] ? _GEN4864 : _GEN3178;
wire  _GEN4866 = io_x[24] ? _GEN4865 : _GEN3180;
wire  _GEN4867 = io_x[17] ? _GEN4866 : _GEN4862;
wire  _GEN4868 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4869 = io_x[10] ? _GEN4868 : _GEN3183;
wire  _GEN4870 = io_x[24] ? _GEN4869 : _GEN3180;
wire  _GEN4871 = io_x[17] ? _GEN4870 : _GEN3243;
wire  _GEN4872 = io_x[12] ? _GEN4871 : _GEN4867;
wire  _GEN4873 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4874 = io_x[24] ? _GEN3196 : _GEN4873;
wire  _GEN4875 = io_x[17] ? _GEN4874 : _GEN3243;
wire  _GEN4876 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4877 = io_x[14] ? _GEN3176 : _GEN4876;
wire  _GEN4878 = io_x[10] ? _GEN4877 : _GEN3183;
wire  _GEN4879 = io_x[24] ? _GEN3180 : _GEN4878;
wire  _GEN4880 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4881 = io_x[14] ? _GEN4880 : _GEN3176;
wire  _GEN4882 = io_x[10] ? _GEN4881 : _GEN3178;
wire  _GEN4883 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4884 = io_x[14] ? _GEN4883 : _GEN3175;
wire  _GEN4885 = io_x[10] ? _GEN4884 : _GEN3183;
wire  _GEN4886 = io_x[24] ? _GEN4885 : _GEN4882;
wire  _GEN4887 = io_x[17] ? _GEN4886 : _GEN4879;
wire  _GEN4888 = io_x[12] ? _GEN4887 : _GEN4875;
wire  _GEN4889 = io_x[2] ? _GEN4888 : _GEN4872;
wire  _GEN4890 = io_x[9] ? _GEN4889 : _GEN4861;
wire  _GEN4891 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4892 = io_x[14] ? _GEN4891 : _GEN3176;
wire  _GEN4893 = io_x[10] ? _GEN3178 : _GEN4892;
wire  _GEN4894 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN4895 = io_x[24] ? _GEN4894 : _GEN4893;
wire  _GEN4896 = io_x[17] ? _GEN4895 : _GEN3174;
wire  _GEN4897 = io_x[12] ? _GEN3958 : _GEN4896;
wire  _GEN4898 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4899 = io_x[10] ? _GEN4898 : _GEN3178;
wire  _GEN4900 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4901 = io_x[10] ? _GEN4900 : _GEN3178;
wire  _GEN4902 = io_x[24] ? _GEN4901 : _GEN4899;
wire  _GEN4903 = io_x[17] ? _GEN4902 : _GEN3243;
wire  _GEN4904 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4905 = io_x[10] ? _GEN4904 : _GEN3178;
wire  _GEN4906 = io_x[24] ? _GEN3180 : _GEN4905;
wire  _GEN4907 = io_x[17] ? _GEN3174 : _GEN4906;
wire  _GEN4908 = io_x[12] ? _GEN4907 : _GEN4903;
wire  _GEN4909 = io_x[2] ? _GEN4908 : _GEN4897;
wire  _GEN4910 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4911 = io_x[10] ? _GEN4910 : _GEN3178;
wire  _GEN4912 = io_x[24] ? _GEN3196 : _GEN4911;
wire  _GEN4913 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN4914 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4915 = io_x[24] ? _GEN4914 : _GEN4913;
wire  _GEN4916 = io_x[17] ? _GEN4915 : _GEN4912;
wire  _GEN4917 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN4918 = io_x[24] ? _GEN3180 : _GEN4917;
wire  _GEN4919 = io_x[17] ? _GEN4918 : _GEN3174;
wire  _GEN4920 = io_x[12] ? _GEN4919 : _GEN4916;
wire  _GEN4921 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4922 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4923 = io_x[14] ? _GEN4922 : _GEN4921;
wire  _GEN4924 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4925 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4926 = io_x[14] ? _GEN4925 : _GEN4924;
wire  _GEN4927 = io_x[10] ? _GEN4926 : _GEN4923;
wire  _GEN4928 = io_x[24] ? _GEN3196 : _GEN4927;
wire  _GEN4929 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4930 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4931 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4932 = io_x[14] ? _GEN4931 : _GEN4930;
wire  _GEN4933 = io_x[10] ? _GEN4932 : _GEN4929;
wire  _GEN4934 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4935 = io_x[14] ? _GEN3176 : _GEN4934;
wire  _GEN4936 = io_x[10] ? _GEN4935 : _GEN3183;
wire  _GEN4937 = io_x[24] ? _GEN4936 : _GEN4933;
wire  _GEN4938 = io_x[17] ? _GEN4937 : _GEN4928;
wire  _GEN4939 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4940 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4941 = io_x[24] ? _GEN4940 : _GEN4939;
wire  _GEN4942 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4943 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4944 = io_x[14] ? _GEN3176 : _GEN4943;
wire  _GEN4945 = io_x[10] ? _GEN4944 : _GEN3183;
wire  _GEN4946 = io_x[24] ? _GEN4945 : _GEN4942;
wire  _GEN4947 = io_x[17] ? _GEN4946 : _GEN4941;
wire  _GEN4948 = io_x[12] ? _GEN4947 : _GEN4938;
wire  _GEN4949 = io_x[2] ? _GEN4948 : _GEN4920;
wire  _GEN4950 = io_x[9] ? _GEN4949 : _GEN4909;
wire  _GEN4951 = io_x[13] ? _GEN4950 : _GEN4890;
wire  _GEN4952 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4953 = io_x[14] ? _GEN4952 : _GEN3176;
wire  _GEN4954 = io_x[10] ? _GEN4953 : _GEN3178;
wire  _GEN4955 = io_x[24] ? _GEN3196 : _GEN4954;
wire  _GEN4956 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4957 = io_x[10] ? _GEN4956 : _GEN3183;
wire  _GEN4958 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN4959 = io_x[24] ? _GEN4958 : _GEN4957;
wire  _GEN4960 = io_x[17] ? _GEN4959 : _GEN4955;
wire  _GEN4961 = io_x[12] ? _GEN4960 : _GEN3370;
wire  _GEN4962 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4963 = io_x[14] ? _GEN4962 : _GEN3175;
wire  _GEN4964 = io_x[10] ? _GEN3183 : _GEN4963;
wire  _GEN4965 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN4966 = io_x[24] ? _GEN4965 : _GEN4964;
wire  _GEN4967 = io_x[17] ? _GEN4966 : _GEN3243;
wire  _GEN4968 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4969 = io_x[14] ? _GEN4968 : _GEN3176;
wire  _GEN4970 = io_x[10] ? _GEN4969 : _GEN3178;
wire  _GEN4971 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4972 = io_x[14] ? _GEN4971 : _GEN3176;
wire  _GEN4973 = io_x[10] ? _GEN4972 : _GEN3178;
wire  _GEN4974 = io_x[24] ? _GEN4973 : _GEN4970;
wire  _GEN4975 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4976 = io_x[14] ? _GEN4975 : _GEN3176;
wire  _GEN4977 = io_x[10] ? _GEN4976 : _GEN3183;
wire  _GEN4978 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4979 = io_x[14] ? _GEN4978 : _GEN3176;
wire  _GEN4980 = io_x[10] ? _GEN4979 : _GEN3178;
wire  _GEN4981 = io_x[24] ? _GEN4980 : _GEN4977;
wire  _GEN4982 = io_x[17] ? _GEN4981 : _GEN4974;
wire  _GEN4983 = io_x[12] ? _GEN4982 : _GEN4967;
wire  _GEN4984 = io_x[2] ? _GEN4983 : _GEN4961;
wire  _GEN4985 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN4986 = io_x[10] ? _GEN3183 : _GEN4985;
wire  _GEN4987 = io_x[24] ? _GEN4986 : _GEN3196;
wire  _GEN4988 = io_x[17] ? _GEN4987 : _GEN3243;
wire  _GEN4989 = io_x[12] ? _GEN4988 : _GEN3958;
wire  _GEN4990 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN4991 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN4992 = io_x[14] ? _GEN4991 : _GEN3176;
wire  _GEN4993 = io_x[10] ? _GEN4992 : _GEN4990;
wire  _GEN4994 = io_x[24] ? _GEN3180 : _GEN4993;
wire  _GEN4995 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN4996 = io_x[24] ? _GEN3180 : _GEN4995;
wire  _GEN4997 = io_x[17] ? _GEN4996 : _GEN4994;
wire  _GEN4998 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN4999 = io_x[14] ? _GEN4998 : _GEN3175;
wire  _GEN5000 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5001 = io_x[14] ? _GEN5000 : _GEN3176;
wire  _GEN5002 = io_x[10] ? _GEN5001 : _GEN4999;
wire  _GEN5003 = io_x[24] ? _GEN3180 : _GEN5002;
wire  _GEN5004 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5005 = io_x[14] ? _GEN5004 : _GEN3175;
wire  _GEN5006 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5007 = io_x[14] ? _GEN5006 : _GEN3176;
wire  _GEN5008 = io_x[10] ? _GEN5007 : _GEN5005;
wire  _GEN5009 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5010 = io_x[14] ? _GEN5009 : _GEN3175;
wire  _GEN5011 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5012 = io_x[14] ? _GEN5011 : _GEN3176;
wire  _GEN5013 = io_x[10] ? _GEN5012 : _GEN5010;
wire  _GEN5014 = io_x[24] ? _GEN5013 : _GEN5008;
wire  _GEN5015 = io_x[17] ? _GEN5014 : _GEN5003;
wire  _GEN5016 = io_x[12] ? _GEN5015 : _GEN4997;
wire  _GEN5017 = io_x[2] ? _GEN5016 : _GEN4989;
wire  _GEN5018 = io_x[9] ? _GEN5017 : _GEN4984;
wire  _GEN5019 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5020 = io_x[14] ? _GEN3176 : _GEN5019;
wire  _GEN5021 = io_x[10] ? _GEN5020 : _GEN3178;
wire  _GEN5022 = io_x[24] ? _GEN3196 : _GEN5021;
wire  _GEN5023 = io_x[17] ? _GEN5022 : _GEN3243;
wire  _GEN5024 = io_x[12] ? _GEN3370 : _GEN5023;
wire  _GEN5025 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5026 = io_x[14] ? _GEN3176 : _GEN5025;
wire  _GEN5027 = io_x[10] ? _GEN5026 : _GEN3178;
wire  _GEN5028 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5029 = io_x[10] ? _GEN5028 : _GEN3178;
wire  _GEN5030 = io_x[24] ? _GEN5029 : _GEN5027;
wire  _GEN5031 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5032 = io_x[14] ? _GEN3176 : _GEN5031;
wire  _GEN5033 = io_x[10] ? _GEN5032 : _GEN3178;
wire  _GEN5034 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5035 = io_x[14] ? _GEN3176 : _GEN5034;
wire  _GEN5036 = io_x[10] ? _GEN5035 : _GEN3178;
wire  _GEN5037 = io_x[24] ? _GEN5036 : _GEN5033;
wire  _GEN5038 = io_x[17] ? _GEN5037 : _GEN5030;
wire  _GEN5039 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5040 = io_x[14] ? _GEN5039 : _GEN3176;
wire  _GEN5041 = io_x[10] ? _GEN3183 : _GEN5040;
wire  _GEN5042 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5043 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5044 = io_x[14] ? _GEN5043 : _GEN3176;
wire  _GEN5045 = io_x[10] ? _GEN5044 : _GEN5042;
wire  _GEN5046 = io_x[24] ? _GEN5045 : _GEN5041;
wire  _GEN5047 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5048 = io_x[14] ? _GEN3176 : _GEN5047;
wire  _GEN5049 = io_x[10] ? _GEN3183 : _GEN5048;
wire  _GEN5050 = io_x[24] ? _GEN5049 : _GEN3180;
wire  _GEN5051 = io_x[17] ? _GEN5050 : _GEN5046;
wire  _GEN5052 = io_x[12] ? _GEN5051 : _GEN5038;
wire  _GEN5053 = io_x[2] ? _GEN5052 : _GEN5024;
wire  _GEN5054 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5055 = io_x[14] ? _GEN5054 : _GEN3176;
wire  _GEN5056 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5057 = io_x[14] ? _GEN5056 : _GEN3176;
wire  _GEN5058 = io_x[10] ? _GEN5057 : _GEN5055;
wire  _GEN5059 = io_x[24] ? _GEN3196 : _GEN5058;
wire  _GEN5060 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5061 = io_x[14] ? _GEN5060 : _GEN3176;
wire  _GEN5062 = io_x[10] ? _GEN3178 : _GEN5061;
wire  _GEN5063 = io_x[24] ? _GEN3196 : _GEN5062;
wire  _GEN5064 = io_x[17] ? _GEN5063 : _GEN5059;
wire  _GEN5065 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5066 = io_x[10] ? _GEN3178 : _GEN5065;
wire  _GEN5067 = io_x[24] ? _GEN3180 : _GEN5066;
wire  _GEN5068 = io_x[24] ? _GEN3196 : _GEN3180;
wire  _GEN5069 = io_x[17] ? _GEN5068 : _GEN5067;
wire  _GEN5070 = io_x[12] ? _GEN5069 : _GEN5064;
wire  _GEN5071 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5072 = io_x[10] ? _GEN3178 : _GEN5071;
wire  _GEN5073 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5074 = io_x[14] ? _GEN5073 : _GEN3176;
wire  _GEN5075 = io_x[10] ? _GEN3178 : _GEN5074;
wire  _GEN5076 = io_x[24] ? _GEN5075 : _GEN5072;
wire  _GEN5077 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5078 = io_x[14] ? _GEN5077 : _GEN3176;
wire  _GEN5079 = io_x[10] ? _GEN3178 : _GEN5078;
wire  _GEN5080 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5081 = io_x[14] ? _GEN5080 : _GEN3176;
wire  _GEN5082 = io_x[10] ? _GEN3178 : _GEN5081;
wire  _GEN5083 = io_x[24] ? _GEN5082 : _GEN5079;
wire  _GEN5084 = io_x[17] ? _GEN5083 : _GEN5076;
wire  _GEN5085 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5086 = io_x[14] ? _GEN5085 : _GEN3176;
wire  _GEN5087 = io_x[10] ? _GEN5086 : _GEN3183;
wire  _GEN5088 = io_x[24] ? _GEN3196 : _GEN5087;
wire  _GEN5089 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5090 = io_x[14] ? _GEN5089 : _GEN3175;
wire  _GEN5091 = io_x[10] ? _GEN5090 : _GEN3183;
wire  _GEN5092 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5093 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5094 = io_x[14] ? _GEN5093 : _GEN3176;
wire  _GEN5095 = io_x[10] ? _GEN5094 : _GEN5092;
wire  _GEN5096 = io_x[24] ? _GEN5095 : _GEN5091;
wire  _GEN5097 = io_x[17] ? _GEN5096 : _GEN5088;
wire  _GEN5098 = io_x[12] ? _GEN5097 : _GEN5084;
wire  _GEN5099 = io_x[2] ? _GEN5098 : _GEN5070;
wire  _GEN5100 = io_x[9] ? _GEN5099 : _GEN5053;
wire  _GEN5101 = io_x[13] ? _GEN5100 : _GEN5018;
wire  _GEN5102 = io_x[7] ? _GEN5101 : _GEN4951;
wire  _GEN5103 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5104 = io_x[14] ? _GEN3176 : _GEN5103;
wire  _GEN5105 = io_x[10] ? _GEN5104 : _GEN3178;
wire  _GEN5106 = io_x[24] ? _GEN5105 : _GEN3180;
wire  _GEN5107 = io_x[17] ? _GEN5106 : _GEN3174;
wire  _GEN5108 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5109 = io_x[10] ? _GEN5108 : _GEN3178;
wire  _GEN5110 = io_x[24] ? _GEN3180 : _GEN5109;
wire  _GEN5111 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5112 = io_x[10] ? _GEN5111 : _GEN3178;
wire  _GEN5113 = io_x[24] ? _GEN3180 : _GEN5112;
wire  _GEN5114 = io_x[17] ? _GEN5113 : _GEN5110;
wire  _GEN5115 = io_x[12] ? _GEN5114 : _GEN5107;
wire  _GEN5116 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5117 = io_x[10] ? _GEN5116 : _GEN3178;
wire  _GEN5118 = io_x[24] ? _GEN3180 : _GEN5117;
wire  _GEN5119 = io_x[17] ? _GEN5118 : _GEN3174;
wire  _GEN5120 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5121 = io_x[10] ? _GEN5120 : _GEN3178;
wire  _GEN5122 = io_x[24] ? _GEN5121 : _GEN3196;
wire  _GEN5123 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5124 = io_x[14] ? _GEN5123 : _GEN3175;
wire  _GEN5125 = io_x[10] ? _GEN5124 : _GEN3178;
wire  _GEN5126 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5127 = io_x[14] ? _GEN5126 : _GEN3175;
wire  _GEN5128 = io_x[10] ? _GEN5127 : _GEN3178;
wire  _GEN5129 = io_x[24] ? _GEN5128 : _GEN5125;
wire  _GEN5130 = io_x[17] ? _GEN5129 : _GEN5122;
wire  _GEN5131 = io_x[12] ? _GEN5130 : _GEN5119;
wire  _GEN5132 = io_x[2] ? _GEN5131 : _GEN5115;
wire  _GEN5133 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5134 = io_x[14] ? _GEN5133 : _GEN3176;
wire  _GEN5135 = io_x[10] ? _GEN5134 : _GEN3178;
wire  _GEN5136 = io_x[24] ? _GEN5135 : _GEN3180;
wire  _GEN5137 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5138 = io_x[14] ? _GEN5137 : _GEN3175;
wire  _GEN5139 = io_x[10] ? _GEN5138 : _GEN3178;
wire  _GEN5140 = io_x[24] ? _GEN5139 : _GEN3180;
wire  _GEN5141 = io_x[17] ? _GEN5140 : _GEN5136;
wire  _GEN5142 = io_x[12] ? _GEN3958 : _GEN5141;
wire  _GEN5143 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5144 = io_x[14] ? _GEN5143 : _GEN3175;
wire  _GEN5145 = io_x[10] ? _GEN3178 : _GEN5144;
wire  _GEN5146 = io_x[24] ? _GEN3196 : _GEN5145;
wire  _GEN5147 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN5148 = io_x[24] ? _GEN3180 : _GEN5147;
wire  _GEN5149 = io_x[17] ? _GEN5148 : _GEN5146;
wire  _GEN5150 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5151 = io_x[14] ? _GEN3176 : _GEN5150;
wire  _GEN5152 = io_x[10] ? _GEN3183 : _GEN5151;
wire  _GEN5153 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5154 = io_x[14] ? _GEN3175 : _GEN5153;
wire  _GEN5155 = io_x[10] ? _GEN3178 : _GEN5154;
wire  _GEN5156 = io_x[24] ? _GEN5155 : _GEN5152;
wire  _GEN5157 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5158 = io_x[14] ? _GEN3175 : _GEN5157;
wire  _GEN5159 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5160 = io_x[14] ? _GEN5159 : _GEN3175;
wire  _GEN5161 = io_x[10] ? _GEN5160 : _GEN5158;
wire  _GEN5162 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5163 = io_x[14] ? _GEN5162 : _GEN3176;
wire  _GEN5164 = io_x[10] ? _GEN5163 : _GEN3183;
wire  _GEN5165 = io_x[24] ? _GEN5164 : _GEN5161;
wire  _GEN5166 = io_x[17] ? _GEN5165 : _GEN5156;
wire  _GEN5167 = io_x[12] ? _GEN5166 : _GEN5149;
wire  _GEN5168 = io_x[2] ? _GEN5167 : _GEN5142;
wire  _GEN5169 = io_x[9] ? _GEN5168 : _GEN5132;
wire  _GEN5170 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5171 = io_x[10] ? _GEN5170 : _GEN3183;
wire  _GEN5172 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5173 = io_x[14] ? _GEN5172 : _GEN3176;
wire  _GEN5174 = io_x[10] ? _GEN5173 : _GEN3178;
wire  _GEN5175 = io_x[24] ? _GEN5174 : _GEN5171;
wire  _GEN5176 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5177 = io_x[10] ? _GEN5176 : _GEN3183;
wire  _GEN5178 = io_x[24] ? _GEN3180 : _GEN5177;
wire  _GEN5179 = io_x[17] ? _GEN5178 : _GEN5175;
wire  _GEN5180 = io_x[24] ? _GEN3196 : _GEN3180;
wire  _GEN5181 = io_x[17] ? _GEN3174 : _GEN5180;
wire  _GEN5182 = io_x[12] ? _GEN5181 : _GEN5179;
wire  _GEN5183 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5184 = io_x[10] ? _GEN5183 : _GEN3183;
wire  _GEN5185 = io_x[24] ? _GEN3180 : _GEN5184;
wire  _GEN5186 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5187 = io_x[14] ? _GEN5186 : _GEN3176;
wire  _GEN5188 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5189 = io_x[10] ? _GEN5188 : _GEN5187;
wire  _GEN5190 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5191 = io_x[14] ? _GEN5190 : _GEN3175;
wire  _GEN5192 = io_x[10] ? _GEN5191 : _GEN3178;
wire  _GEN5193 = io_x[24] ? _GEN5192 : _GEN5189;
wire  _GEN5194 = io_x[17] ? _GEN5193 : _GEN5185;
wire  _GEN5195 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5196 = io_x[14] ? _GEN3176 : _GEN5195;
wire  _GEN5197 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5198 = io_x[10] ? _GEN5197 : _GEN5196;
wire  _GEN5199 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN5200 = io_x[24] ? _GEN5199 : _GEN5198;
wire  _GEN5201 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5202 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5203 = io_x[14] ? _GEN5202 : _GEN5201;
wire  _GEN5204 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5205 = io_x[10] ? _GEN5204 : _GEN5203;
wire  _GEN5206 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5207 = io_x[14] ? _GEN3176 : _GEN5206;
wire  _GEN5208 = io_x[10] ? _GEN3183 : _GEN5207;
wire  _GEN5209 = io_x[24] ? _GEN5208 : _GEN5205;
wire  _GEN5210 = io_x[17] ? _GEN5209 : _GEN5200;
wire  _GEN5211 = io_x[12] ? _GEN5210 : _GEN5194;
wire  _GEN5212 = io_x[2] ? _GEN5211 : _GEN5182;
wire  _GEN5213 = io_x[24] ? _GEN3196 : _GEN3180;
wire  _GEN5214 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5215 = io_x[14] ? _GEN5214 : _GEN3176;
wire  _GEN5216 = io_x[10] ? _GEN5215 : _GEN3178;
wire  _GEN5217 = io_x[24] ? _GEN3180 : _GEN5216;
wire  _GEN5218 = io_x[17] ? _GEN5217 : _GEN5213;
wire  _GEN5219 = io_x[24] ? _GEN3180 : _GEN3196;
wire  _GEN5220 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5221 = io_x[14] ? _GEN5220 : _GEN3175;
wire  _GEN5222 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5223 = io_x[14] ? _GEN5222 : _GEN3176;
wire  _GEN5224 = io_x[10] ? _GEN5223 : _GEN5221;
wire  _GEN5225 = io_x[24] ? _GEN5224 : _GEN3196;
wire  _GEN5226 = io_x[17] ? _GEN5225 : _GEN5219;
wire  _GEN5227 = io_x[12] ? _GEN5226 : _GEN5218;
wire  _GEN5228 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5229 = io_x[14] ? _GEN3175 : _GEN5228;
wire  _GEN5230 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5231 = io_x[14] ? _GEN5230 : _GEN3176;
wire  _GEN5232 = io_x[10] ? _GEN5231 : _GEN5229;
wire  _GEN5233 = io_x[24] ? _GEN3180 : _GEN5232;
wire  _GEN5234 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5235 = io_x[14] ? _GEN5234 : _GEN3176;
wire  _GEN5236 = io_x[10] ? _GEN5235 : _GEN3178;
wire  _GEN5237 = io_x[24] ? _GEN3196 : _GEN5236;
wire  _GEN5238 = io_x[17] ? _GEN5237 : _GEN5233;
wire  _GEN5239 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5240 = io_x[10] ? _GEN3178 : _GEN5239;
wire  _GEN5241 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN5242 = io_x[24] ? _GEN5241 : _GEN5240;
wire  _GEN5243 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5244 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5245 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5246 = io_x[14] ? _GEN5245 : _GEN5244;
wire  _GEN5247 = io_x[10] ? _GEN5246 : _GEN5243;
wire  _GEN5248 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5249 = io_x[14] ? _GEN5248 : _GEN3176;
wire  _GEN5250 = io_x[10] ? _GEN5249 : _GEN3183;
wire  _GEN5251 = io_x[24] ? _GEN5250 : _GEN5247;
wire  _GEN5252 = io_x[17] ? _GEN5251 : _GEN5242;
wire  _GEN5253 = io_x[12] ? _GEN5252 : _GEN5238;
wire  _GEN5254 = io_x[2] ? _GEN5253 : _GEN5227;
wire  _GEN5255 = io_x[9] ? _GEN5254 : _GEN5212;
wire  _GEN5256 = io_x[13] ? _GEN5255 : _GEN5169;
wire  _GEN5257 = io_x[17] ? _GEN3243 : _GEN3174;
wire  _GEN5258 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5259 = io_x[14] ? _GEN5258 : _GEN3176;
wire  _GEN5260 = io_x[10] ? _GEN3178 : _GEN5259;
wire  _GEN5261 = io_x[24] ? _GEN3196 : _GEN5260;
wire  _GEN5262 = io_x[17] ? _GEN3174 : _GEN5261;
wire  _GEN5263 = io_x[12] ? _GEN5262 : _GEN5257;
wire  _GEN5264 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5265 = io_x[10] ? _GEN3178 : _GEN5264;
wire  _GEN5266 = io_x[24] ? _GEN3180 : _GEN5265;
wire  _GEN5267 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5268 = io_x[10] ? _GEN3178 : _GEN5267;
wire  _GEN5269 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5270 = io_x[14] ? _GEN5269 : _GEN3175;
wire  _GEN5271 = io_x[10] ? _GEN5270 : _GEN3183;
wire  _GEN5272 = io_x[24] ? _GEN5271 : _GEN5268;
wire  _GEN5273 = io_x[17] ? _GEN5272 : _GEN5266;
wire  _GEN5274 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5275 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5276 = io_x[14] ? _GEN5275 : _GEN5274;
wire  _GEN5277 = io_x[10] ? _GEN5276 : _GEN3178;
wire  _GEN5278 = io_x[24] ? _GEN5277 : _GEN3196;
wire  _GEN5279 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5280 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5281 = io_x[14] ? _GEN5280 : _GEN5279;
wire  _GEN5282 = io_x[10] ? _GEN5281 : _GEN3178;
wire  _GEN5283 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5284 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5285 = io_x[14] ? _GEN5284 : _GEN5283;
wire  _GEN5286 = io_x[10] ? _GEN5285 : _GEN3183;
wire  _GEN5287 = io_x[24] ? _GEN5286 : _GEN5282;
wire  _GEN5288 = io_x[17] ? _GEN5287 : _GEN5278;
wire  _GEN5289 = io_x[12] ? _GEN5288 : _GEN5273;
wire  _GEN5290 = io_x[2] ? _GEN5289 : _GEN5263;
wire  _GEN5291 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5292 = io_x[14] ? _GEN5291 : _GEN3175;
wire  _GEN5293 = io_x[10] ? _GEN5292 : _GEN3183;
wire  _GEN5294 = io_x[24] ? _GEN3196 : _GEN5293;
wire  _GEN5295 = io_x[17] ? _GEN5294 : _GEN3243;
wire  _GEN5296 = io_x[12] ? _GEN5295 : _GEN3370;
wire  _GEN5297 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN5298 = io_x[24] ? _GEN3180 : _GEN5297;
wire  _GEN5299 = io_x[17] ? _GEN3174 : _GEN5298;
wire  _GEN5300 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5301 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5302 = io_x[14] ? _GEN5301 : _GEN5300;
wire  _GEN5303 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5304 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5305 = io_x[14] ? _GEN5304 : _GEN5303;
wire  _GEN5306 = io_x[10] ? _GEN5305 : _GEN5302;
wire  _GEN5307 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5308 = io_x[14] ? _GEN5307 : _GEN3176;
wire  _GEN5309 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5310 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5311 = io_x[14] ? _GEN5310 : _GEN5309;
wire  _GEN5312 = io_x[10] ? _GEN5311 : _GEN5308;
wire  _GEN5313 = io_x[24] ? _GEN5312 : _GEN5306;
wire  _GEN5314 = io_x[17] ? _GEN5313 : _GEN3174;
wire  _GEN5315 = io_x[12] ? _GEN5314 : _GEN5299;
wire  _GEN5316 = io_x[2] ? _GEN5315 : _GEN5296;
wire  _GEN5317 = io_x[9] ? _GEN5316 : _GEN5290;
wire  _GEN5318 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5319 = io_x[14] ? _GEN5318 : _GEN3176;
wire  _GEN5320 = io_x[10] ? _GEN5319 : _GEN3178;
wire  _GEN5321 = io_x[24] ? _GEN5320 : _GEN3180;
wire  _GEN5322 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5323 = io_x[14] ? _GEN5322 : _GEN3175;
wire  _GEN5324 = io_x[10] ? _GEN5323 : _GEN3178;
wire  _GEN5325 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5326 = io_x[14] ? _GEN5325 : _GEN3175;
wire  _GEN5327 = io_x[10] ? _GEN5326 : _GEN3178;
wire  _GEN5328 = io_x[24] ? _GEN5327 : _GEN5324;
wire  _GEN5329 = io_x[17] ? _GEN5328 : _GEN5321;
wire  _GEN5330 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5331 = io_x[10] ? _GEN5330 : _GEN3178;
wire  _GEN5332 = io_x[24] ? _GEN3196 : _GEN5331;
wire  _GEN5333 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5334 = io_x[14] ? _GEN3176 : _GEN5333;
wire  _GEN5335 = io_x[10] ? _GEN5334 : _GEN3178;
wire  _GEN5336 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5337 = io_x[14] ? _GEN3176 : _GEN5336;
wire  _GEN5338 = io_x[10] ? _GEN5337 : _GEN3178;
wire  _GEN5339 = io_x[24] ? _GEN5338 : _GEN5335;
wire  _GEN5340 = io_x[17] ? _GEN5339 : _GEN5332;
wire  _GEN5341 = io_x[12] ? _GEN5340 : _GEN5329;
wire  _GEN5342 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5343 = io_x[10] ? _GEN5342 : _GEN3178;
wire  _GEN5344 = io_x[24] ? _GEN3196 : _GEN5343;
wire  _GEN5345 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5346 = io_x[14] ? _GEN5345 : _GEN3176;
wire  _GEN5347 = io_x[10] ? _GEN5346 : _GEN3183;
wire  _GEN5348 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5349 = io_x[14] ? _GEN5348 : _GEN3175;
wire  _GEN5350 = io_x[10] ? _GEN5349 : _GEN3178;
wire  _GEN5351 = io_x[24] ? _GEN5350 : _GEN5347;
wire  _GEN5352 = io_x[17] ? _GEN5351 : _GEN5344;
wire  _GEN5353 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5354 = io_x[14] ? _GEN3176 : _GEN5353;
wire  _GEN5355 = io_x[10] ? _GEN5354 : _GEN3178;
wire  _GEN5356 = io_x[24] ? _GEN3196 : _GEN5355;
wire  _GEN5357 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5358 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5359 = io_x[14] ? _GEN5358 : _GEN5357;
wire  _GEN5360 = io_x[10] ? _GEN5359 : _GEN3178;
wire  _GEN5361 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5362 = io_x[14] ? _GEN3175 : _GEN5361;
wire  _GEN5363 = io_x[10] ? _GEN5362 : _GEN3178;
wire  _GEN5364 = io_x[24] ? _GEN5363 : _GEN5360;
wire  _GEN5365 = io_x[17] ? _GEN5364 : _GEN5356;
wire  _GEN5366 = io_x[12] ? _GEN5365 : _GEN5352;
wire  _GEN5367 = io_x[2] ? _GEN5366 : _GEN5341;
wire  _GEN5368 = io_x[24] ? _GEN3196 : _GEN3180;
wire  _GEN5369 = io_x[24] ? _GEN3196 : _GEN3180;
wire  _GEN5370 = io_x[17] ? _GEN5369 : _GEN5368;
wire  _GEN5371 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5372 = io_x[14] ? _GEN5371 : _GEN3176;
wire  _GEN5373 = io_x[10] ? _GEN5372 : _GEN3178;
wire  _GEN5374 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5375 = io_x[14] ? _GEN5374 : _GEN3176;
wire  _GEN5376 = io_x[10] ? _GEN5375 : _GEN3183;
wire  _GEN5377 = io_x[24] ? _GEN5376 : _GEN5373;
wire  _GEN5378 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5379 = io_x[10] ? _GEN3178 : _GEN5378;
wire  _GEN5380 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5381 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5382 = io_x[14] ? _GEN5381 : _GEN3176;
wire  _GEN5383 = io_x[10] ? _GEN5382 : _GEN5380;
wire  _GEN5384 = io_x[24] ? _GEN5383 : _GEN5379;
wire  _GEN5385 = io_x[17] ? _GEN5384 : _GEN5377;
wire  _GEN5386 = io_x[12] ? _GEN5385 : _GEN5370;
wire  _GEN5387 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5388 = io_x[14] ? _GEN3176 : _GEN5387;
wire  _GEN5389 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5390 = io_x[10] ? _GEN5389 : _GEN5388;
wire  _GEN5391 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5392 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5393 = io_x[14] ? _GEN5392 : _GEN5391;
wire  _GEN5394 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5395 = io_x[10] ? _GEN5394 : _GEN5393;
wire  _GEN5396 = io_x[24] ? _GEN5395 : _GEN5390;
wire  _GEN5397 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5398 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5399 = io_x[14] ? _GEN5398 : _GEN5397;
wire  _GEN5400 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5401 = io_x[10] ? _GEN5400 : _GEN5399;
wire  _GEN5402 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5403 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5404 = io_x[14] ? _GEN5403 : _GEN5402;
wire  _GEN5405 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5406 = io_x[10] ? _GEN5405 : _GEN5404;
wire  _GEN5407 = io_x[24] ? _GEN5406 : _GEN5401;
wire  _GEN5408 = io_x[17] ? _GEN5407 : _GEN5396;
wire  _GEN5409 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5410 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5411 = io_x[14] ? _GEN5410 : _GEN5409;
wire  _GEN5412 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5413 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5414 = io_x[14] ? _GEN5413 : _GEN5412;
wire  _GEN5415 = io_x[10] ? _GEN5414 : _GEN5411;
wire  _GEN5416 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5417 = io_x[14] ? _GEN5416 : _GEN3176;
wire  _GEN5418 = io_x[10] ? _GEN5417 : _GEN3183;
wire  _GEN5419 = io_x[24] ? _GEN5418 : _GEN5415;
wire  _GEN5420 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5421 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5422 = io_x[14] ? _GEN5421 : _GEN5420;
wire  _GEN5423 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5424 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5425 = io_x[14] ? _GEN5424 : _GEN5423;
wire  _GEN5426 = io_x[10] ? _GEN5425 : _GEN5422;
wire  _GEN5427 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5428 = io_x[14] ? _GEN3175 : _GEN5427;
wire  _GEN5429 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5430 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5431 = io_x[14] ? _GEN5430 : _GEN5429;
wire  _GEN5432 = io_x[10] ? _GEN5431 : _GEN5428;
wire  _GEN5433 = io_x[24] ? _GEN5432 : _GEN5426;
wire  _GEN5434 = io_x[17] ? _GEN5433 : _GEN5419;
wire  _GEN5435 = io_x[12] ? _GEN5434 : _GEN5408;
wire  _GEN5436 = io_x[2] ? _GEN5435 : _GEN5386;
wire  _GEN5437 = io_x[9] ? _GEN5436 : _GEN5367;
wire  _GEN5438 = io_x[13] ? _GEN5437 : _GEN5317;
wire  _GEN5439 = io_x[7] ? _GEN5438 : _GEN5256;
wire  _GEN5440 = io_x[15] ? _GEN5439 : _GEN5102;
wire  _GEN5441 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN5442 = io_x[24] ? _GEN3180 : _GEN5441;
wire  _GEN5443 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5444 = io_x[14] ? _GEN5443 : _GEN3175;
wire  _GEN5445 = io_x[10] ? _GEN3178 : _GEN5444;
wire  _GEN5446 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5447 = io_x[14] ? _GEN5446 : _GEN3176;
wire  _GEN5448 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5449 = io_x[10] ? _GEN5448 : _GEN5447;
wire  _GEN5450 = io_x[24] ? _GEN5449 : _GEN5445;
wire  _GEN5451 = io_x[17] ? _GEN5450 : _GEN5442;
wire  _GEN5452 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5453 = io_x[14] ? _GEN5452 : _GEN3175;
wire  _GEN5454 = io_x[10] ? _GEN5453 : _GEN3178;
wire  _GEN5455 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN5456 = io_x[24] ? _GEN5455 : _GEN5454;
wire  _GEN5457 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5458 = io_x[14] ? _GEN5457 : _GEN3175;
wire  _GEN5459 = io_x[10] ? _GEN5458 : _GEN3178;
wire  _GEN5460 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN5461 = io_x[24] ? _GEN5460 : _GEN5459;
wire  _GEN5462 = io_x[17] ? _GEN5461 : _GEN5456;
wire  _GEN5463 = io_x[12] ? _GEN5462 : _GEN5451;
wire  _GEN5464 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5465 = io_x[14] ? _GEN5464 : _GEN3176;
wire  _GEN5466 = io_x[10] ? _GEN3178 : _GEN5465;
wire  _GEN5467 = io_x[24] ? _GEN3180 : _GEN5466;
wire  _GEN5468 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5469 = io_x[14] ? _GEN5468 : _GEN3176;
wire  _GEN5470 = io_x[10] ? _GEN3178 : _GEN5469;
wire  _GEN5471 = io_x[24] ? _GEN3180 : _GEN5470;
wire  _GEN5472 = io_x[17] ? _GEN5471 : _GEN5467;
wire  _GEN5473 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5474 = io_x[14] ? _GEN5473 : _GEN3176;
wire  _GEN5475 = io_x[10] ? _GEN5474 : _GEN3183;
wire  _GEN5476 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5477 = io_x[14] ? _GEN5476 : _GEN3176;
wire  _GEN5478 = io_x[10] ? _GEN3178 : _GEN5477;
wire  _GEN5479 = io_x[24] ? _GEN5478 : _GEN5475;
wire  _GEN5480 = io_x[17] ? _GEN5479 : _GEN3174;
wire  _GEN5481 = io_x[12] ? _GEN5480 : _GEN5472;
wire  _GEN5482 = io_x[2] ? _GEN5481 : _GEN5463;
wire  _GEN5483 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5484 = io_x[10] ? _GEN5483 : _GEN3178;
wire  _GEN5485 = io_x[24] ? _GEN5484 : _GEN3196;
wire  _GEN5486 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5487 = io_x[10] ? _GEN5486 : _GEN3178;
wire  _GEN5488 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5489 = io_x[14] ? _GEN5488 : _GEN3176;
wire  _GEN5490 = io_x[10] ? _GEN5489 : _GEN3183;
wire  _GEN5491 = io_x[24] ? _GEN5490 : _GEN5487;
wire  _GEN5492 = io_x[17] ? _GEN5491 : _GEN5485;
wire  _GEN5493 = io_x[12] ? _GEN5492 : _GEN3370;
wire  _GEN5494 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5495 = io_x[14] ? _GEN5494 : _GEN3176;
wire  _GEN5496 = io_x[10] ? _GEN5495 : _GEN3178;
wire  _GEN5497 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5498 = io_x[10] ? _GEN5497 : _GEN3178;
wire  _GEN5499 = io_x[24] ? _GEN5498 : _GEN5496;
wire  _GEN5500 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5501 = io_x[14] ? _GEN5500 : _GEN3176;
wire  _GEN5502 = io_x[10] ? _GEN5501 : _GEN3183;
wire  _GEN5503 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN5504 = io_x[24] ? _GEN5503 : _GEN5502;
wire  _GEN5505 = io_x[17] ? _GEN5504 : _GEN5499;
wire  _GEN5506 = io_x[12] ? _GEN5505 : _GEN3958;
wire  _GEN5507 = io_x[2] ? _GEN5506 : _GEN5493;
wire  _GEN5508 = io_x[9] ? _GEN5507 : _GEN5482;
wire  _GEN5509 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5510 = io_x[10] ? _GEN5509 : _GEN3178;
wire  _GEN5511 = io_x[24] ? _GEN5510 : _GEN3180;
wire  _GEN5512 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5513 = io_x[14] ? _GEN5512 : _GEN3176;
wire  _GEN5514 = io_x[10] ? _GEN5513 : _GEN3178;
wire  _GEN5515 = io_x[24] ? _GEN3180 : _GEN5514;
wire  _GEN5516 = io_x[17] ? _GEN5515 : _GEN5511;
wire  _GEN5517 = io_x[24] ? _GEN3196 : _GEN3180;
wire  _GEN5518 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5519 = io_x[14] ? _GEN5518 : _GEN3175;
wire  _GEN5520 = io_x[10] ? _GEN3183 : _GEN5519;
wire  _GEN5521 = io_x[24] ? _GEN5520 : _GEN3180;
wire  _GEN5522 = io_x[17] ? _GEN5521 : _GEN5517;
wire  _GEN5523 = io_x[12] ? _GEN5522 : _GEN5516;
wire  _GEN5524 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5525 = io_x[14] ? _GEN3176 : _GEN5524;
wire  _GEN5526 = io_x[10] ? _GEN5525 : _GEN3178;
wire  _GEN5527 = io_x[24] ? _GEN3196 : _GEN5526;
wire  _GEN5528 = io_x[17] ? _GEN5527 : _GEN3243;
wire  _GEN5529 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5530 = io_x[10] ? _GEN5529 : _GEN3178;
wire  _GEN5531 = io_x[24] ? _GEN3180 : _GEN5530;
wire  _GEN5532 = io_x[17] ? _GEN5531 : _GEN3174;
wire  _GEN5533 = io_x[12] ? _GEN5532 : _GEN5528;
wire  _GEN5534 = io_x[2] ? _GEN5533 : _GEN5523;
wire  _GEN5535 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5536 = io_x[10] ? _GEN5535 : _GEN3178;
wire  _GEN5537 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5538 = io_x[10] ? _GEN5537 : _GEN3178;
wire  _GEN5539 = io_x[24] ? _GEN5538 : _GEN5536;
wire  _GEN5540 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5541 = io_x[14] ? _GEN5540 : _GEN3176;
wire  _GEN5542 = io_x[10] ? _GEN5541 : _GEN3178;
wire  _GEN5543 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5544 = io_x[14] ? _GEN5543 : _GEN3176;
wire  _GEN5545 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5546 = io_x[14] ? _GEN3175 : _GEN5545;
wire  _GEN5547 = io_x[10] ? _GEN5546 : _GEN5544;
wire  _GEN5548 = io_x[24] ? _GEN5547 : _GEN5542;
wire  _GEN5549 = io_x[17] ? _GEN5548 : _GEN5539;
wire  _GEN5550 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5551 = io_x[14] ? _GEN5550 : _GEN3175;
wire  _GEN5552 = io_x[10] ? _GEN5551 : _GEN3178;
wire  _GEN5553 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5554 = io_x[14] ? _GEN5553 : _GEN3176;
wire  _GEN5555 = io_x[10] ? _GEN5554 : _GEN3178;
wire  _GEN5556 = io_x[24] ? _GEN5555 : _GEN5552;
wire  _GEN5557 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5558 = io_x[14] ? _GEN5557 : _GEN3175;
wire  _GEN5559 = io_x[10] ? _GEN5558 : _GEN3178;
wire  _GEN5560 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5561 = io_x[14] ? _GEN5560 : _GEN3176;
wire  _GEN5562 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5563 = io_x[14] ? _GEN5562 : _GEN3176;
wire  _GEN5564 = io_x[10] ? _GEN5563 : _GEN5561;
wire  _GEN5565 = io_x[24] ? _GEN5564 : _GEN5559;
wire  _GEN5566 = io_x[17] ? _GEN5565 : _GEN5556;
wire  _GEN5567 = io_x[12] ? _GEN5566 : _GEN5549;
wire  _GEN5568 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5569 = io_x[14] ? _GEN3176 : _GEN5568;
wire  _GEN5570 = io_x[10] ? _GEN5569 : _GEN3178;
wire  _GEN5571 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5572 = io_x[14] ? _GEN5571 : _GEN3175;
wire  _GEN5573 = io_x[10] ? _GEN3178 : _GEN5572;
wire  _GEN5574 = io_x[24] ? _GEN5573 : _GEN5570;
wire  _GEN5575 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5576 = io_x[14] ? _GEN3176 : _GEN5575;
wire  _GEN5577 = io_x[10] ? _GEN5576 : _GEN3183;
wire  _GEN5578 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5579 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5580 = io_x[14] ? _GEN5579 : _GEN5578;
wire  _GEN5581 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5582 = io_x[14] ? _GEN3176 : _GEN5581;
wire  _GEN5583 = io_x[10] ? _GEN5582 : _GEN5580;
wire  _GEN5584 = io_x[24] ? _GEN5583 : _GEN5577;
wire  _GEN5585 = io_x[17] ? _GEN5584 : _GEN5574;
wire  _GEN5586 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN5587 = io_x[24] ? _GEN3180 : _GEN5586;
wire  _GEN5588 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN5589 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5590 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5591 = io_x[14] ? _GEN5590 : _GEN3176;
wire  _GEN5592 = io_x[10] ? _GEN5591 : _GEN5589;
wire  _GEN5593 = io_x[24] ? _GEN5592 : _GEN5588;
wire  _GEN5594 = io_x[17] ? _GEN5593 : _GEN5587;
wire  _GEN5595 = io_x[12] ? _GEN5594 : _GEN5585;
wire  _GEN5596 = io_x[2] ? _GEN5595 : _GEN5567;
wire  _GEN5597 = io_x[9] ? _GEN5596 : _GEN5534;
wire  _GEN5598 = io_x[13] ? _GEN5597 : _GEN5508;
wire  _GEN5599 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5600 = io_x[14] ? _GEN5599 : _GEN3176;
wire  _GEN5601 = io_x[10] ? _GEN5600 : _GEN3178;
wire  _GEN5602 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5603 = io_x[14] ? _GEN5602 : _GEN3176;
wire  _GEN5604 = io_x[10] ? _GEN5603 : _GEN3178;
wire  _GEN5605 = io_x[24] ? _GEN5604 : _GEN5601;
wire  _GEN5606 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5607 = io_x[14] ? _GEN5606 : _GEN3176;
wire  _GEN5608 = io_x[10] ? _GEN5607 : _GEN3178;
wire  _GEN5609 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5610 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5611 = io_x[14] ? _GEN5610 : _GEN3176;
wire  _GEN5612 = io_x[10] ? _GEN5611 : _GEN5609;
wire  _GEN5613 = io_x[24] ? _GEN5612 : _GEN5608;
wire  _GEN5614 = io_x[17] ? _GEN5613 : _GEN5605;
wire  _GEN5615 = io_x[12] ? _GEN5614 : _GEN3958;
wire  _GEN5616 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5617 = io_x[14] ? _GEN5616 : _GEN3176;
wire  _GEN5618 = io_x[10] ? _GEN5617 : _GEN3183;
wire  _GEN5619 = io_x[24] ? _GEN3180 : _GEN5618;
wire  _GEN5620 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5621 = io_x[14] ? _GEN5620 : _GEN3175;
wire  _GEN5622 = io_x[10] ? _GEN5621 : _GEN3178;
wire  _GEN5623 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5624 = io_x[14] ? _GEN5623 : _GEN3176;
wire  _GEN5625 = io_x[10] ? _GEN5624 : _GEN3178;
wire  _GEN5626 = io_x[24] ? _GEN5625 : _GEN5622;
wire  _GEN5627 = io_x[17] ? _GEN5626 : _GEN5619;
wire  _GEN5628 = io_x[12] ? _GEN5627 : _GEN3958;
wire  _GEN5629 = io_x[2] ? _GEN5628 : _GEN5615;
wire  _GEN5630 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5631 = io_x[14] ? _GEN5630 : _GEN3176;
wire  _GEN5632 = io_x[10] ? _GEN3178 : _GEN5631;
wire  _GEN5633 = io_x[24] ? _GEN5632 : _GEN3180;
wire  _GEN5634 = io_x[17] ? _GEN3174 : _GEN5633;
wire  _GEN5635 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN5636 = io_x[24] ? _GEN5635 : _GEN3196;
wire  _GEN5637 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5638 = io_x[14] ? _GEN5637 : _GEN3176;
wire  _GEN5639 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5640 = io_x[14] ? _GEN5639 : _GEN3176;
wire  _GEN5641 = io_x[10] ? _GEN5640 : _GEN5638;
wire  _GEN5642 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5643 = io_x[14] ? _GEN5642 : _GEN3175;
wire  _GEN5644 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5645 = io_x[10] ? _GEN5644 : _GEN5643;
wire  _GEN5646 = io_x[24] ? _GEN5645 : _GEN5641;
wire  _GEN5647 = io_x[17] ? _GEN5646 : _GEN5636;
wire  _GEN5648 = io_x[12] ? _GEN5647 : _GEN5634;
wire  _GEN5649 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5650 = io_x[14] ? _GEN5649 : _GEN3176;
wire  _GEN5651 = io_x[10] ? _GEN5650 : _GEN3183;
wire  _GEN5652 = io_x[24] ? _GEN3180 : _GEN5651;
wire  _GEN5653 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5654 = io_x[14] ? _GEN5653 : _GEN3176;
wire  _GEN5655 = io_x[10] ? _GEN5654 : _GEN3178;
wire  _GEN5656 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5657 = io_x[14] ? _GEN5656 : _GEN3176;
wire  _GEN5658 = io_x[10] ? _GEN3178 : _GEN5657;
wire  _GEN5659 = io_x[24] ? _GEN5658 : _GEN5655;
wire  _GEN5660 = io_x[17] ? _GEN5659 : _GEN5652;
wire  _GEN5661 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5662 = io_x[14] ? _GEN5661 : _GEN3176;
wire  _GEN5663 = io_x[10] ? _GEN3178 : _GEN5662;
wire  _GEN5664 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN5665 = io_x[24] ? _GEN5664 : _GEN5663;
wire  _GEN5666 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5667 = io_x[14] ? _GEN5666 : _GEN3176;
wire  _GEN5668 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5669 = io_x[10] ? _GEN5668 : _GEN5667;
wire  _GEN5670 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5671 = io_x[14] ? _GEN5670 : _GEN3176;
wire  _GEN5672 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5673 = io_x[14] ? _GEN5672 : _GEN3176;
wire  _GEN5674 = io_x[10] ? _GEN5673 : _GEN5671;
wire  _GEN5675 = io_x[24] ? _GEN5674 : _GEN5669;
wire  _GEN5676 = io_x[17] ? _GEN5675 : _GEN5665;
wire  _GEN5677 = io_x[12] ? _GEN5676 : _GEN5660;
wire  _GEN5678 = io_x[2] ? _GEN5677 : _GEN5648;
wire  _GEN5679 = io_x[9] ? _GEN5678 : _GEN5629;
wire  _GEN5680 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5681 = io_x[14] ? _GEN3176 : _GEN5680;
wire  _GEN5682 = io_x[10] ? _GEN5681 : _GEN3178;
wire  _GEN5683 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5684 = io_x[14] ? _GEN3176 : _GEN5683;
wire  _GEN5685 = io_x[10] ? _GEN5684 : _GEN3178;
wire  _GEN5686 = io_x[24] ? _GEN5685 : _GEN5682;
wire  _GEN5687 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5688 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5689 = io_x[14] ? _GEN5688 : _GEN5687;
wire  _GEN5690 = io_x[10] ? _GEN5689 : _GEN3178;
wire  _GEN5691 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5692 = io_x[14] ? _GEN3176 : _GEN5691;
wire  _GEN5693 = io_x[10] ? _GEN5692 : _GEN3178;
wire  _GEN5694 = io_x[24] ? _GEN5693 : _GEN5690;
wire  _GEN5695 = io_x[17] ? _GEN5694 : _GEN5686;
wire  _GEN5696 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5697 = io_x[14] ? _GEN5696 : _GEN3176;
wire  _GEN5698 = io_x[10] ? _GEN3183 : _GEN5697;
wire  _GEN5699 = io_x[24] ? _GEN3196 : _GEN5698;
wire  _GEN5700 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN5701 = io_x[24] ? _GEN3196 : _GEN5700;
wire  _GEN5702 = io_x[17] ? _GEN5701 : _GEN5699;
wire  _GEN5703 = io_x[12] ? _GEN5702 : _GEN5695;
wire  _GEN5704 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5705 = io_x[14] ? _GEN3176 : _GEN5704;
wire  _GEN5706 = io_x[10] ? _GEN5705 : _GEN3178;
wire  _GEN5707 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN5708 = io_x[24] ? _GEN5707 : _GEN5706;
wire  _GEN5709 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5710 = io_x[14] ? _GEN3176 : _GEN5709;
wire  _GEN5711 = io_x[10] ? _GEN5710 : _GEN3183;
wire  _GEN5712 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN5713 = io_x[24] ? _GEN5712 : _GEN5711;
wire  _GEN5714 = io_x[17] ? _GEN5713 : _GEN5708;
wire  _GEN5715 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN5716 = io_x[24] ? _GEN5715 : _GEN3180;
wire  _GEN5717 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5718 = io_x[10] ? _GEN3178 : _GEN5717;
wire  _GEN5719 = io_x[24] ? _GEN5718 : _GEN3180;
wire  _GEN5720 = io_x[17] ? _GEN5719 : _GEN5716;
wire  _GEN5721 = io_x[12] ? _GEN5720 : _GEN5714;
wire  _GEN5722 = io_x[2] ? _GEN5721 : _GEN5703;
wire  _GEN5723 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5724 = io_x[14] ? _GEN5723 : _GEN3175;
wire  _GEN5725 = io_x[10] ? _GEN3178 : _GEN5724;
wire  _GEN5726 = io_x[24] ? _GEN5725 : _GEN3180;
wire  _GEN5727 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5728 = io_x[14] ? _GEN5727 : _GEN3176;
wire  _GEN5729 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5730 = io_x[14] ? _GEN3175 : _GEN5729;
wire  _GEN5731 = io_x[10] ? _GEN5730 : _GEN5728;
wire  _GEN5732 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5733 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5734 = io_x[14] ? _GEN5733 : _GEN5732;
wire  _GEN5735 = io_x[10] ? _GEN3178 : _GEN5734;
wire  _GEN5736 = io_x[24] ? _GEN5735 : _GEN5731;
wire  _GEN5737 = io_x[17] ? _GEN5736 : _GEN5726;
wire  _GEN5738 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5739 = io_x[14] ? _GEN5738 : _GEN3176;
wire  _GEN5740 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5741 = io_x[14] ? _GEN5740 : _GEN3176;
wire  _GEN5742 = io_x[10] ? _GEN5741 : _GEN5739;
wire  _GEN5743 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5744 = io_x[14] ? _GEN5743 : _GEN3176;
wire  _GEN5745 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5746 = io_x[14] ? _GEN5745 : _GEN3175;
wire  _GEN5747 = io_x[10] ? _GEN5746 : _GEN5744;
wire  _GEN5748 = io_x[24] ? _GEN5747 : _GEN5742;
wire  _GEN5749 = io_x[17] ? _GEN5748 : _GEN3174;
wire  _GEN5750 = io_x[12] ? _GEN5749 : _GEN5737;
wire  _GEN5751 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5752 = io_x[14] ? _GEN5751 : _GEN3176;
wire  _GEN5753 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5754 = io_x[14] ? _GEN3176 : _GEN5753;
wire  _GEN5755 = io_x[10] ? _GEN5754 : _GEN5752;
wire  _GEN5756 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5757 = io_x[10] ? _GEN3183 : _GEN5756;
wire  _GEN5758 = io_x[24] ? _GEN5757 : _GEN5755;
wire  _GEN5759 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5760 = io_x[14] ? _GEN5759 : _GEN3175;
wire  _GEN5761 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5762 = io_x[10] ? _GEN5761 : _GEN5760;
wire  _GEN5763 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5764 = io_x[14] ? _GEN5763 : _GEN3176;
wire  _GEN5765 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5766 = io_x[10] ? _GEN5765 : _GEN5764;
wire  _GEN5767 = io_x[24] ? _GEN5766 : _GEN5762;
wire  _GEN5768 = io_x[17] ? _GEN5767 : _GEN5758;
wire  _GEN5769 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5770 = io_x[14] ? _GEN3175 : _GEN5769;
wire  _GEN5771 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5772 = io_x[14] ? _GEN5771 : _GEN3176;
wire  _GEN5773 = io_x[10] ? _GEN5772 : _GEN5770;
wire  _GEN5774 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5775 = io_x[14] ? _GEN5774 : _GEN3176;
wire  _GEN5776 = io_x[10] ? _GEN5775 : _GEN3178;
wire  _GEN5777 = io_x[24] ? _GEN5776 : _GEN5773;
wire  _GEN5778 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5779 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5780 = io_x[14] ? _GEN5779 : _GEN5778;
wire  _GEN5781 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5782 = io_x[14] ? _GEN5781 : _GEN3175;
wire  _GEN5783 = io_x[10] ? _GEN5782 : _GEN5780;
wire  _GEN5784 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5785 = io_x[14] ? _GEN5784 : _GEN3176;
wire  _GEN5786 = io_x[10] ? _GEN5785 : _GEN3183;
wire  _GEN5787 = io_x[24] ? _GEN5786 : _GEN5783;
wire  _GEN5788 = io_x[17] ? _GEN5787 : _GEN5777;
wire  _GEN5789 = io_x[12] ? _GEN5788 : _GEN5768;
wire  _GEN5790 = io_x[2] ? _GEN5789 : _GEN5750;
wire  _GEN5791 = io_x[9] ? _GEN5790 : _GEN5722;
wire  _GEN5792 = io_x[13] ? _GEN5791 : _GEN5679;
wire  _GEN5793 = io_x[7] ? _GEN5792 : _GEN5598;
wire  _GEN5794 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5795 = io_x[14] ? _GEN5794 : _GEN3176;
wire  _GEN5796 = io_x[10] ? _GEN3178 : _GEN5795;
wire  _GEN5797 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5798 = io_x[14] ? _GEN5797 : _GEN3176;
wire  _GEN5799 = io_x[10] ? _GEN3178 : _GEN5798;
wire  _GEN5800 = io_x[24] ? _GEN5799 : _GEN5796;
wire  _GEN5801 = io_x[17] ? _GEN5800 : _GEN3174;
wire  _GEN5802 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5803 = io_x[14] ? _GEN3176 : _GEN5802;
wire  _GEN5804 = io_x[10] ? _GEN5803 : _GEN3178;
wire  _GEN5805 = io_x[24] ? _GEN3196 : _GEN5804;
wire  _GEN5806 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5807 = io_x[14] ? _GEN3176 : _GEN5806;
wire  _GEN5808 = io_x[10] ? _GEN5807 : _GEN3178;
wire  _GEN5809 = io_x[24] ? _GEN3196 : _GEN5808;
wire  _GEN5810 = io_x[17] ? _GEN5809 : _GEN5805;
wire  _GEN5811 = io_x[12] ? _GEN5810 : _GEN5801;
wire  _GEN5812 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5813 = io_x[14] ? _GEN5812 : _GEN3176;
wire  _GEN5814 = io_x[10] ? _GEN3178 : _GEN5813;
wire  _GEN5815 = io_x[24] ? _GEN3180 : _GEN5814;
wire  _GEN5816 = io_x[10] ? _GEN3178 : _GEN5469;
wire  _GEN5817 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN5818 = io_x[24] ? _GEN5817 : _GEN5816;
wire  _GEN5819 = io_x[17] ? _GEN5818 : _GEN5815;
wire  _GEN5820 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5821 = io_x[14] ? _GEN3176 : _GEN5820;
wire  _GEN5822 = io_x[10] ? _GEN5821 : _GEN3178;
wire  _GEN5823 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5824 = io_x[10] ? _GEN5823 : _GEN3178;
wire  _GEN5825 = io_x[24] ? _GEN5824 : _GEN5822;
wire  _GEN5826 = io_x[17] ? _GEN5825 : _GEN3174;
wire  _GEN5827 = io_x[12] ? _GEN5826 : _GEN5819;
wire  _GEN5828 = io_x[2] ? _GEN5827 : _GEN5811;
wire  _GEN5829 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5830 = io_x[10] ? _GEN3178 : _GEN5829;
wire  _GEN5831 = io_x[24] ? _GEN5830 : _GEN3180;
wire  _GEN5832 = io_x[17] ? _GEN5831 : _GEN3174;
wire  _GEN5833 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5834 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5835 = io_x[10] ? _GEN5834 : _GEN5833;
wire  _GEN5836 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5837 = io_x[10] ? _GEN5836 : _GEN3183;
wire  _GEN5838 = io_x[24] ? _GEN5837 : _GEN5835;
wire  _GEN5839 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5840 = io_x[14] ? _GEN5839 : _GEN3176;
wire  _GEN5841 = io_x[10] ? _GEN5840 : _GEN3183;
wire  _GEN5842 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5843 = io_x[14] ? _GEN5842 : _GEN3175;
wire  _GEN5844 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5845 = io_x[10] ? _GEN5844 : _GEN5843;
wire  _GEN5846 = io_x[24] ? _GEN5845 : _GEN5841;
wire  _GEN5847 = io_x[17] ? _GEN5846 : _GEN5838;
wire  _GEN5848 = io_x[12] ? _GEN5847 : _GEN5832;
wire  _GEN5849 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5850 = io_x[14] ? _GEN5849 : _GEN3175;
wire  _GEN5851 = io_x[10] ? _GEN3178 : _GEN5850;
wire  _GEN5852 = io_x[24] ? _GEN5851 : _GEN3196;
wire  _GEN5853 = io_x[17] ? _GEN5852 : _GEN3243;
wire  _GEN5854 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5855 = io_x[14] ? _GEN5854 : _GEN3175;
wire  _GEN5856 = io_x[10] ? _GEN5855 : _GEN3178;
wire  _GEN5857 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5858 = io_x[10] ? _GEN3183 : _GEN5857;
wire  _GEN5859 = io_x[24] ? _GEN5858 : _GEN5856;
wire  _GEN5860 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5861 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5862 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5863 = io_x[14] ? _GEN5862 : _GEN5861;
wire  _GEN5864 = io_x[10] ? _GEN5863 : _GEN5860;
wire  _GEN5865 = io_x[24] ? _GEN3180 : _GEN5864;
wire  _GEN5866 = io_x[17] ? _GEN5865 : _GEN5859;
wire  _GEN5867 = io_x[12] ? _GEN5866 : _GEN5853;
wire  _GEN5868 = io_x[2] ? _GEN5867 : _GEN5848;
wire  _GEN5869 = io_x[9] ? _GEN5868 : _GEN5828;
wire  _GEN5870 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5871 = io_x[14] ? _GEN3175 : _GEN5870;
wire  _GEN5872 = io_x[10] ? _GEN5871 : _GEN3178;
wire  _GEN5873 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5874 = io_x[10] ? _GEN5873 : _GEN3183;
wire  _GEN5875 = io_x[24] ? _GEN5874 : _GEN5872;
wire  _GEN5876 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5877 = io_x[14] ? _GEN3175 : _GEN5876;
wire  _GEN5878 = io_x[10] ? _GEN5877 : _GEN3178;
wire  _GEN5879 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5880 = io_x[10] ? _GEN5879 : _GEN3183;
wire  _GEN5881 = io_x[24] ? _GEN5880 : _GEN5878;
wire  _GEN5882 = io_x[17] ? _GEN5881 : _GEN5875;
wire  _GEN5883 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5884 = io_x[14] ? _GEN3176 : _GEN5883;
wire  _GEN5885 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5886 = io_x[10] ? _GEN5885 : _GEN5884;
wire  _GEN5887 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5888 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5889 = io_x[14] ? _GEN5888 : _GEN5887;
wire  _GEN5890 = io_x[10] ? _GEN3178 : _GEN5889;
wire  _GEN5891 = io_x[24] ? _GEN5890 : _GEN5886;
wire  _GEN5892 = io_x[17] ? _GEN5891 : _GEN3243;
wire  _GEN5893 = io_x[12] ? _GEN5892 : _GEN5882;
wire  _GEN5894 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5895 = io_x[10] ? _GEN5894 : _GEN3178;
wire  _GEN5896 = io_x[24] ? _GEN3180 : _GEN5895;
wire  _GEN5897 = io_x[17] ? _GEN5896 : _GEN3243;
wire  _GEN5898 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5899 = io_x[14] ? _GEN3175 : _GEN5898;
wire  _GEN5900 = io_x[10] ? _GEN3183 : _GEN5899;
wire  _GEN5901 = io_x[24] ? _GEN3196 : _GEN5900;
wire  _GEN5902 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5903 = io_x[14] ? _GEN3175 : _GEN5902;
wire  _GEN5904 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN5905 = io_x[10] ? _GEN5904 : _GEN5903;
wire  _GEN5906 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5907 = io_x[14] ? _GEN5906 : _GEN3176;
wire  _GEN5908 = io_x[10] ? _GEN3183 : _GEN5907;
wire  _GEN5909 = io_x[24] ? _GEN5908 : _GEN5905;
wire  _GEN5910 = io_x[17] ? _GEN5909 : _GEN5901;
wire  _GEN5911 = io_x[12] ? _GEN5910 : _GEN5897;
wire  _GEN5912 = io_x[2] ? _GEN5911 : _GEN5893;
wire  _GEN5913 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5914 = io_x[10] ? _GEN3178 : _GEN5913;
wire  _GEN5915 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5916 = io_x[14] ? _GEN3176 : _GEN5915;
wire  _GEN5917 = io_x[10] ? _GEN5916 : _GEN3183;
wire  _GEN5918 = io_x[24] ? _GEN5917 : _GEN5914;
wire  _GEN5919 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5920 = io_x[14] ? _GEN5919 : _GEN3176;
wire  _GEN5921 = io_x[10] ? _GEN5920 : _GEN3178;
wire  _GEN5922 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5923 = io_x[14] ? _GEN3175 : _GEN5922;
wire  _GEN5924 = io_x[10] ? _GEN5923 : _GEN3183;
wire  _GEN5925 = io_x[24] ? _GEN5924 : _GEN5921;
wire  _GEN5926 = io_x[17] ? _GEN5925 : _GEN5918;
wire  _GEN5927 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5928 = io_x[14] ? _GEN3176 : _GEN5927;
wire  _GEN5929 = io_x[10] ? _GEN5928 : _GEN3178;
wire  _GEN5930 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5931 = io_x[10] ? _GEN5930 : _GEN3178;
wire  _GEN5932 = io_x[24] ? _GEN5931 : _GEN5929;
wire  _GEN5933 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5934 = io_x[14] ? _GEN5933 : _GEN3175;
wire  _GEN5935 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5936 = io_x[14] ? _GEN5935 : _GEN3176;
wire  _GEN5937 = io_x[10] ? _GEN5936 : _GEN5934;
wire  _GEN5938 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5939 = io_x[10] ? _GEN5938 : _GEN3178;
wire  _GEN5940 = io_x[24] ? _GEN5939 : _GEN5937;
wire  _GEN5941 = io_x[17] ? _GEN5940 : _GEN5932;
wire  _GEN5942 = io_x[12] ? _GEN5941 : _GEN5926;
wire  _GEN5943 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5944 = io_x[14] ? _GEN5943 : _GEN3175;
wire  _GEN5945 = io_x[10] ? _GEN5944 : _GEN3178;
wire  _GEN5946 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5947 = io_x[14] ? _GEN3176 : _GEN5946;
wire  _GEN5948 = io_x[10] ? _GEN3183 : _GEN5947;
wire  _GEN5949 = io_x[24] ? _GEN5948 : _GEN5945;
wire  _GEN5950 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5951 = io_x[14] ? _GEN5950 : _GEN3175;
wire  _GEN5952 = io_x[10] ? _GEN5951 : _GEN3183;
wire  _GEN5953 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5954 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5955 = io_x[14] ? _GEN5954 : _GEN5953;
wire  _GEN5956 = io_x[10] ? _GEN3183 : _GEN5955;
wire  _GEN5957 = io_x[24] ? _GEN5956 : _GEN5952;
wire  _GEN5958 = io_x[17] ? _GEN5957 : _GEN5949;
wire  _GEN5959 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5960 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5961 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5962 = io_x[14] ? _GEN5961 : _GEN5960;
wire  _GEN5963 = io_x[10] ? _GEN5962 : _GEN5959;
wire  _GEN5964 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5965 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5966 = io_x[14] ? _GEN5965 : _GEN5964;
wire  _GEN5967 = io_x[10] ? _GEN5966 : _GEN3178;
wire  _GEN5968 = io_x[24] ? _GEN5967 : _GEN5963;
wire  _GEN5969 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN5970 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5971 = io_x[14] ? _GEN5970 : _GEN3176;
wire  _GEN5972 = io_x[10] ? _GEN5971 : _GEN5969;
wire  _GEN5973 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5974 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5975 = io_x[14] ? _GEN5974 : _GEN5973;
wire  _GEN5976 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5977 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN5978 = io_x[14] ? _GEN5977 : _GEN5976;
wire  _GEN5979 = io_x[10] ? _GEN5978 : _GEN5975;
wire  _GEN5980 = io_x[24] ? _GEN5979 : _GEN5972;
wire  _GEN5981 = io_x[17] ? _GEN5980 : _GEN5968;
wire  _GEN5982 = io_x[12] ? _GEN5981 : _GEN5958;
wire  _GEN5983 = io_x[2] ? _GEN5982 : _GEN5942;
wire  _GEN5984 = io_x[9] ? _GEN5983 : _GEN5912;
wire  _GEN5985 = io_x[13] ? _GEN5984 : _GEN5869;
wire  _GEN5986 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5987 = io_x[14] ? _GEN5986 : _GEN3176;
wire  _GEN5988 = io_x[10] ? _GEN5987 : _GEN3178;
wire  _GEN5989 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN5990 = io_x[24] ? _GEN5989 : _GEN5988;
wire  _GEN5991 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5992 = io_x[14] ? _GEN5991 : _GEN3176;
wire  _GEN5993 = io_x[10] ? _GEN5992 : _GEN3183;
wire  _GEN5994 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN5995 = io_x[14] ? _GEN5994 : _GEN3176;
wire  _GEN5996 = io_x[10] ? _GEN5995 : _GEN3183;
wire  _GEN5997 = io_x[24] ? _GEN5996 : _GEN5993;
wire  _GEN5998 = io_x[17] ? _GEN5997 : _GEN5990;
wire  _GEN5999 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6000 = io_x[14] ? _GEN5999 : _GEN3176;
wire  _GEN6001 = io_x[10] ? _GEN6000 : _GEN3183;
wire  _GEN6002 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6003 = io_x[14] ? _GEN6002 : _GEN3176;
wire  _GEN6004 = io_x[10] ? _GEN6003 : _GEN3178;
wire  _GEN6005 = io_x[24] ? _GEN6004 : _GEN6001;
wire  _GEN6006 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6007 = io_x[14] ? _GEN6006 : _GEN3175;
wire  _GEN6008 = io_x[10] ? _GEN6007 : _GEN3183;
wire  _GEN6009 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6010 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6011 = io_x[14] ? _GEN6010 : _GEN6009;
wire  _GEN6012 = io_x[10] ? _GEN6011 : _GEN3178;
wire  _GEN6013 = io_x[24] ? _GEN6012 : _GEN6008;
wire  _GEN6014 = io_x[17] ? _GEN6013 : _GEN6005;
wire  _GEN6015 = io_x[12] ? _GEN6014 : _GEN5998;
wire  _GEN6016 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6017 = io_x[14] ? _GEN6016 : _GEN3175;
wire  _GEN6018 = io_x[10] ? _GEN6017 : _GEN3183;
wire  _GEN6019 = io_x[24] ? _GEN6018 : _GEN3180;
wire  _GEN6020 = io_x[17] ? _GEN6019 : _GEN3243;
wire  _GEN6021 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6022 = io_x[14] ? _GEN6021 : _GEN3176;
wire  _GEN6023 = io_x[10] ? _GEN6022 : _GEN3178;
wire  _GEN6024 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN6025 = io_x[24] ? _GEN6024 : _GEN6023;
wire  _GEN6026 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6027 = io_x[14] ? _GEN3176 : _GEN6026;
wire  _GEN6028 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6029 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6030 = io_x[14] ? _GEN6029 : _GEN6028;
wire  _GEN6031 = io_x[10] ? _GEN6030 : _GEN6027;
wire  _GEN6032 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6033 = io_x[14] ? _GEN6032 : _GEN3175;
wire  _GEN6034 = io_x[10] ? _GEN6033 : _GEN3183;
wire  _GEN6035 = io_x[24] ? _GEN6034 : _GEN6031;
wire  _GEN6036 = io_x[17] ? _GEN6035 : _GEN6025;
wire  _GEN6037 = io_x[12] ? _GEN6036 : _GEN6020;
wire  _GEN6038 = io_x[2] ? _GEN6037 : _GEN6015;
wire  _GEN6039 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6040 = io_x[14] ? _GEN6039 : _GEN3175;
wire  _GEN6041 = io_x[10] ? _GEN3178 : _GEN6040;
wire  _GEN6042 = io_x[24] ? _GEN3180 : _GEN6041;
wire  _GEN6043 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6044 = io_x[14] ? _GEN6043 : _GEN3175;
wire  _GEN6045 = io_x[10] ? _GEN3178 : _GEN6044;
wire  _GEN6046 = io_x[24] ? _GEN3180 : _GEN6045;
wire  _GEN6047 = io_x[17] ? _GEN6046 : _GEN6042;
wire  _GEN6048 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6049 = io_x[14] ? _GEN3176 : _GEN6048;
wire  _GEN6050 = io_x[10] ? _GEN3183 : _GEN6049;
wire  _GEN6051 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6052 = io_x[14] ? _GEN6051 : _GEN3176;
wire  _GEN6053 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6054 = io_x[14] ? _GEN6053 : _GEN3175;
wire  _GEN6055 = io_x[10] ? _GEN6054 : _GEN6052;
wire  _GEN6056 = io_x[24] ? _GEN6055 : _GEN6050;
wire  _GEN6057 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN6058 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6059 = io_x[14] ? _GEN3175 : _GEN6058;
wire  _GEN6060 = io_x[10] ? _GEN6059 : _GEN6057;
wire  _GEN6061 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN6062 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN6063 = io_x[10] ? _GEN6062 : _GEN6061;
wire  _GEN6064 = io_x[24] ? _GEN6063 : _GEN6060;
wire  _GEN6065 = io_x[17] ? _GEN6064 : _GEN6056;
wire  _GEN6066 = io_x[12] ? _GEN6065 : _GEN6047;
wire  _GEN6067 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6068 = io_x[14] ? _GEN6067 : _GEN3176;
wire  _GEN6069 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6070 = io_x[14] ? _GEN6069 : _GEN3176;
wire  _GEN6071 = io_x[10] ? _GEN6070 : _GEN6068;
wire  _GEN6072 = io_x[24] ? _GEN3180 : _GEN6071;
wire  _GEN6073 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6074 = io_x[14] ? _GEN6073 : _GEN3176;
wire  _GEN6075 = io_x[14] ? _GEN3176 : _GEN3175;
wire  _GEN6076 = io_x[10] ? _GEN6075 : _GEN6074;
wire  _GEN6077 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6078 = io_x[14] ? _GEN6077 : _GEN3176;
wire  _GEN6079 = io_x[10] ? _GEN3183 : _GEN6078;
wire  _GEN6080 = io_x[24] ? _GEN6079 : _GEN6076;
wire  _GEN6081 = io_x[17] ? _GEN6080 : _GEN6072;
wire  _GEN6082 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6083 = io_x[14] ? _GEN6082 : _GEN3175;
wire  _GEN6084 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6085 = io_x[14] ? _GEN3176 : _GEN6084;
wire  _GEN6086 = io_x[10] ? _GEN6085 : _GEN6083;
wire  _GEN6087 = io_x[24] ? _GEN3196 : _GEN6086;
wire  _GEN6088 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6089 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6090 = io_x[14] ? _GEN6089 : _GEN6088;
wire  _GEN6091 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6092 = io_x[14] ? _GEN3176 : _GEN6091;
wire  _GEN6093 = io_x[10] ? _GEN6092 : _GEN6090;
wire  _GEN6094 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6095 = io_x[14] ? _GEN3175 : _GEN6094;
wire  _GEN6096 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6097 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6098 = io_x[14] ? _GEN6097 : _GEN6096;
wire  _GEN6099 = io_x[10] ? _GEN6098 : _GEN6095;
wire  _GEN6100 = io_x[24] ? _GEN6099 : _GEN6093;
wire  _GEN6101 = io_x[17] ? _GEN6100 : _GEN6087;
wire  _GEN6102 = io_x[12] ? _GEN6101 : _GEN6081;
wire  _GEN6103 = io_x[2] ? _GEN6102 : _GEN6066;
wire  _GEN6104 = io_x[9] ? _GEN6103 : _GEN6038;
wire  _GEN6105 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6106 = io_x[14] ? _GEN6105 : _GEN3175;
wire  _GEN6107 = io_x[10] ? _GEN6106 : _GEN3178;
wire  _GEN6108 = io_x[24] ? _GEN6107 : _GEN3196;
wire  _GEN6109 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6110 = io_x[14] ? _GEN6109 : _GEN3175;
wire  _GEN6111 = io_x[10] ? _GEN6110 : _GEN3178;
wire  _GEN6112 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6113 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6114 = io_x[14] ? _GEN6113 : _GEN6112;
wire  _GEN6115 = io_x[10] ? _GEN6114 : _GEN3183;
wire  _GEN6116 = io_x[24] ? _GEN6115 : _GEN6111;
wire  _GEN6117 = io_x[17] ? _GEN6116 : _GEN6108;
wire  _GEN6118 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6119 = io_x[14] ? _GEN3176 : _GEN6118;
wire  _GEN6120 = io_x[10] ? _GEN6119 : _GEN3178;
wire  _GEN6121 = io_x[24] ? _GEN6120 : _GEN3180;
wire  _GEN6122 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6123 = io_x[14] ? _GEN3175 : _GEN6122;
wire  _GEN6124 = io_x[10] ? _GEN6123 : _GEN3178;
wire  _GEN6125 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6126 = io_x[14] ? _GEN3176 : _GEN6125;
wire  _GEN6127 = io_x[10] ? _GEN6126 : _GEN3178;
wire  _GEN6128 = io_x[24] ? _GEN6127 : _GEN6124;
wire  _GEN6129 = io_x[17] ? _GEN6128 : _GEN6121;
wire  _GEN6130 = io_x[12] ? _GEN6129 : _GEN6117;
wire  _GEN6131 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6132 = io_x[14] ? _GEN6131 : _GEN3176;
wire  _GEN6133 = io_x[10] ? _GEN6132 : _GEN3178;
wire  _GEN6134 = io_x[10] ? _GEN3178 : _GEN3183;
wire  _GEN6135 = io_x[24] ? _GEN6134 : _GEN6133;
wire  _GEN6136 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6137 = io_x[14] ? _GEN3176 : _GEN6136;
wire  _GEN6138 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6139 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6140 = io_x[14] ? _GEN6139 : _GEN6138;
wire  _GEN6141 = io_x[10] ? _GEN6140 : _GEN6137;
wire  _GEN6142 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6143 = io_x[14] ? _GEN6142 : _GEN3176;
wire  _GEN6144 = io_x[10] ? _GEN6143 : _GEN3178;
wire  _GEN6145 = io_x[24] ? _GEN6144 : _GEN6141;
wire  _GEN6146 = io_x[17] ? _GEN6145 : _GEN6135;
wire  _GEN6147 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6148 = io_x[14] ? _GEN6147 : _GEN3176;
wire  _GEN6149 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6150 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6151 = io_x[14] ? _GEN6150 : _GEN6149;
wire  _GEN6152 = io_x[10] ? _GEN6151 : _GEN6148;
wire  _GEN6153 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6154 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6155 = io_x[14] ? _GEN6154 : _GEN6153;
wire  _GEN6156 = io_x[10] ? _GEN6155 : _GEN3178;
wire  _GEN6157 = io_x[24] ? _GEN6156 : _GEN6152;
wire  _GEN6158 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN6159 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6160 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6161 = io_x[14] ? _GEN6160 : _GEN6159;
wire  _GEN6162 = io_x[10] ? _GEN6161 : _GEN6158;
wire  _GEN6163 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6164 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6165 = io_x[14] ? _GEN6164 : _GEN6163;
wire  _GEN6166 = io_x[10] ? _GEN6165 : _GEN3183;
wire  _GEN6167 = io_x[24] ? _GEN6166 : _GEN6162;
wire  _GEN6168 = io_x[17] ? _GEN6167 : _GEN6157;
wire  _GEN6169 = io_x[12] ? _GEN6168 : _GEN6146;
wire  _GEN6170 = io_x[2] ? _GEN6169 : _GEN6130;
wire  _GEN6171 = io_x[14] ? _GEN3175 : _GEN3176;
wire  _GEN6172 = io_x[10] ? _GEN3183 : _GEN6171;
wire  _GEN6173 = io_x[24] ? _GEN6172 : _GEN3196;
wire  _GEN6174 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6175 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6176 = io_x[14] ? _GEN6175 : _GEN6174;
wire  _GEN6177 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6178 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6179 = io_x[14] ? _GEN6178 : _GEN6177;
wire  _GEN6180 = io_x[10] ? _GEN6179 : _GEN6176;
wire  _GEN6181 = io_x[10] ? _GEN3183 : _GEN3178;
wire  _GEN6182 = io_x[24] ? _GEN6181 : _GEN6180;
wire  _GEN6183 = io_x[17] ? _GEN6182 : _GEN6173;
wire  _GEN6184 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6185 = io_x[14] ? _GEN6184 : _GEN3176;
wire  _GEN6186 = io_x[10] ? _GEN6185 : _GEN3183;
wire  _GEN6187 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6188 = io_x[14] ? _GEN3176 : _GEN6187;
wire  _GEN6189 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6190 = io_x[14] ? _GEN6189 : _GEN3175;
wire  _GEN6191 = io_x[10] ? _GEN6190 : _GEN6188;
wire  _GEN6192 = io_x[24] ? _GEN6191 : _GEN6186;
wire  _GEN6193 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6194 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6195 = io_x[14] ? _GEN6194 : _GEN6193;
wire  _GEN6196 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6197 = io_x[14] ? _GEN6196 : _GEN3176;
wire  _GEN6198 = io_x[10] ? _GEN6197 : _GEN6195;
wire  _GEN6199 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6200 = io_x[14] ? _GEN3175 : _GEN6199;
wire  _GEN6201 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6202 = io_x[14] ? _GEN6201 : _GEN3175;
wire  _GEN6203 = io_x[10] ? _GEN6202 : _GEN6200;
wire  _GEN6204 = io_x[24] ? _GEN6203 : _GEN6198;
wire  _GEN6205 = io_x[17] ? _GEN6204 : _GEN6192;
wire  _GEN6206 = io_x[12] ? _GEN6205 : _GEN6183;
wire  _GEN6207 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6208 = io_x[14] ? _GEN6207 : _GEN3175;
wire  _GEN6209 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6210 = io_x[14] ? _GEN6209 : _GEN3176;
wire  _GEN6211 = io_x[10] ? _GEN6210 : _GEN6208;
wire  _GEN6212 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6213 = io_x[14] ? _GEN3175 : _GEN6212;
wire  _GEN6214 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6215 = io_x[14] ? _GEN3176 : _GEN6214;
wire  _GEN6216 = io_x[10] ? _GEN6215 : _GEN6213;
wire  _GEN6217 = io_x[24] ? _GEN6216 : _GEN6211;
wire  _GEN6218 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6219 = io_x[14] ? _GEN3176 : _GEN6218;
wire  _GEN6220 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6221 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6222 = io_x[14] ? _GEN6221 : _GEN6220;
wire  _GEN6223 = io_x[10] ? _GEN6222 : _GEN6219;
wire  _GEN6224 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6225 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6226 = io_x[14] ? _GEN6225 : _GEN6224;
wire  _GEN6227 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6228 = io_x[14] ? _GEN6227 : _GEN3176;
wire  _GEN6229 = io_x[10] ? _GEN6228 : _GEN6226;
wire  _GEN6230 = io_x[24] ? _GEN6229 : _GEN6223;
wire  _GEN6231 = io_x[17] ? _GEN6230 : _GEN6217;
wire  _GEN6232 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6233 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6234 = io_x[14] ? _GEN6233 : _GEN6232;
wire  _GEN6235 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6236 = io_x[14] ? _GEN6235 : _GEN3175;
wire  _GEN6237 = io_x[10] ? _GEN6236 : _GEN6234;
wire  _GEN6238 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6239 = io_x[14] ? _GEN3175 : _GEN6238;
wire  _GEN6240 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6241 = io_x[14] ? _GEN6240 : _GEN3175;
wire  _GEN6242 = io_x[10] ? _GEN6241 : _GEN6239;
wire  _GEN6243 = io_x[24] ? _GEN6242 : _GEN6237;
wire  _GEN6244 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6245 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6246 = io_x[14] ? _GEN6245 : _GEN6244;
wire  _GEN6247 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6248 = io_x[14] ? _GEN6247 : _GEN3175;
wire  _GEN6249 = io_x[10] ? _GEN6248 : _GEN6246;
wire  _GEN6250 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6251 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6252 = io_x[14] ? _GEN6251 : _GEN6250;
wire  _GEN6253 = io_x[6] ? _GEN3184 : _GEN3185;
wire  _GEN6254 = io_x[6] ? _GEN3185 : _GEN3184;
wire  _GEN6255 = io_x[14] ? _GEN6254 : _GEN6253;
wire  _GEN6256 = io_x[10] ? _GEN6255 : _GEN6252;
wire  _GEN6257 = io_x[24] ? _GEN6256 : _GEN6249;
wire  _GEN6258 = io_x[17] ? _GEN6257 : _GEN6243;
wire  _GEN6259 = io_x[12] ? _GEN6258 : _GEN6231;
wire  _GEN6260 = io_x[2] ? _GEN6259 : _GEN6206;
wire  _GEN6261 = io_x[9] ? _GEN6260 : _GEN6170;
wire  _GEN6262 = io_x[13] ? _GEN6261 : _GEN6104;
wire  _GEN6263 = io_x[7] ? _GEN6262 : _GEN5985;
wire  _GEN6264 = io_x[15] ? _GEN6263 : _GEN5793;
wire  _GEN6265 = io_x[3] ? _GEN6264 : _GEN5440;
wire  _GEN6266 = io_x[27] ? _GEN6265 : _GEN4829;
assign io_y[7] = _GEN6266;
wire  _GEN6267 = 1'b0;
wire  _GEN6268 = 1'b1;
wire  _GEN6269 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6270 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6271 = io_x[9] ? _GEN6270 : _GEN6269;
wire  _GEN6272 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6273 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6274 = io_x[9] ? _GEN6273 : _GEN6272;
wire  _GEN6275 = io_x[24] ? _GEN6274 : _GEN6271;
wire  _GEN6276 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6277 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6278 = io_x[9] ? _GEN6277 : _GEN6276;
wire  _GEN6279 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6280 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6281 = io_x[9] ? _GEN6280 : _GEN6279;
wire  _GEN6282 = io_x[24] ? _GEN6281 : _GEN6278;
wire  _GEN6283 = io_x[26] ? _GEN6282 : _GEN6275;
wire  _GEN6284 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6285 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6286 = io_x[9] ? _GEN6285 : _GEN6284;
wire  _GEN6287 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6288 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6289 = io_x[9] ? _GEN6288 : _GEN6287;
wire  _GEN6290 = io_x[24] ? _GEN6289 : _GEN6286;
wire  _GEN6291 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6292 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6293 = io_x[9] ? _GEN6292 : _GEN6291;
wire  _GEN6294 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6295 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6296 = io_x[9] ? _GEN6295 : _GEN6294;
wire  _GEN6297 = io_x[24] ? _GEN6296 : _GEN6293;
wire  _GEN6298 = io_x[26] ? _GEN6297 : _GEN6290;
wire  _GEN6299 = io_x[5] ? _GEN6298 : _GEN6283;
wire  _GEN6300 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6301 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6302 = io_x[9] ? _GEN6301 : _GEN6300;
wire  _GEN6303 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6304 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6305 = io_x[9] ? _GEN6304 : _GEN6303;
wire  _GEN6306 = io_x[24] ? _GEN6305 : _GEN6302;
wire  _GEN6307 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6308 = 1'b1;
wire  _GEN6309 = io_x[9] ? _GEN6308 : _GEN6307;
wire  _GEN6310 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6311 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6312 = io_x[9] ? _GEN6311 : _GEN6310;
wire  _GEN6313 = io_x[24] ? _GEN6312 : _GEN6309;
wire  _GEN6314 = io_x[26] ? _GEN6313 : _GEN6306;
wire  _GEN6315 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6316 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6317 = io_x[9] ? _GEN6316 : _GEN6315;
wire  _GEN6318 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6319 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6320 = io_x[9] ? _GEN6319 : _GEN6318;
wire  _GEN6321 = io_x[24] ? _GEN6320 : _GEN6317;
wire  _GEN6322 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6323 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6324 = io_x[9] ? _GEN6323 : _GEN6322;
wire  _GEN6325 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6326 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6327 = io_x[9] ? _GEN6326 : _GEN6325;
wire  _GEN6328 = io_x[24] ? _GEN6327 : _GEN6324;
wire  _GEN6329 = io_x[26] ? _GEN6328 : _GEN6321;
wire  _GEN6330 = io_x[5] ? _GEN6329 : _GEN6314;
wire  _GEN6331 = io_x[22] ? _GEN6330 : _GEN6299;
wire  _GEN6332 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6333 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6334 = io_x[9] ? _GEN6333 : _GEN6332;
wire  _GEN6335 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6336 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6337 = io_x[9] ? _GEN6336 : _GEN6335;
wire  _GEN6338 = io_x[24] ? _GEN6337 : _GEN6334;
wire  _GEN6339 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6340 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6341 = io_x[9] ? _GEN6340 : _GEN6339;
wire  _GEN6342 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6343 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6344 = io_x[9] ? _GEN6343 : _GEN6342;
wire  _GEN6345 = io_x[24] ? _GEN6344 : _GEN6341;
wire  _GEN6346 = io_x[26] ? _GEN6345 : _GEN6338;
wire  _GEN6347 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6348 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6349 = io_x[9] ? _GEN6348 : _GEN6347;
wire  _GEN6350 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6351 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6352 = io_x[9] ? _GEN6351 : _GEN6350;
wire  _GEN6353 = io_x[24] ? _GEN6352 : _GEN6349;
wire  _GEN6354 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6355 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6356 = io_x[9] ? _GEN6355 : _GEN6354;
wire  _GEN6357 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6358 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6359 = io_x[9] ? _GEN6358 : _GEN6357;
wire  _GEN6360 = io_x[24] ? _GEN6359 : _GEN6356;
wire  _GEN6361 = io_x[26] ? _GEN6360 : _GEN6353;
wire  _GEN6362 = io_x[5] ? _GEN6361 : _GEN6346;
wire  _GEN6363 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6364 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6365 = io_x[9] ? _GEN6364 : _GEN6363;
wire  _GEN6366 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6367 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6368 = io_x[9] ? _GEN6367 : _GEN6366;
wire  _GEN6369 = io_x[24] ? _GEN6368 : _GEN6365;
wire  _GEN6370 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6371 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6372 = io_x[9] ? _GEN6371 : _GEN6370;
wire  _GEN6373 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6374 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6375 = io_x[9] ? _GEN6374 : _GEN6373;
wire  _GEN6376 = io_x[24] ? _GEN6375 : _GEN6372;
wire  _GEN6377 = io_x[26] ? _GEN6376 : _GEN6369;
wire  _GEN6378 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6379 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6380 = io_x[9] ? _GEN6379 : _GEN6378;
wire  _GEN6381 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6382 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6383 = io_x[9] ? _GEN6382 : _GEN6381;
wire  _GEN6384 = io_x[24] ? _GEN6383 : _GEN6380;
wire  _GEN6385 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6386 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6387 = io_x[9] ? _GEN6386 : _GEN6385;
wire  _GEN6388 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6389 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6390 = io_x[9] ? _GEN6389 : _GEN6388;
wire  _GEN6391 = io_x[24] ? _GEN6390 : _GEN6387;
wire  _GEN6392 = io_x[26] ? _GEN6391 : _GEN6384;
wire  _GEN6393 = io_x[5] ? _GEN6392 : _GEN6377;
wire  _GEN6394 = io_x[22] ? _GEN6393 : _GEN6362;
wire  _GEN6395 = io_x[13] ? _GEN6394 : _GEN6331;
wire  _GEN6396 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6397 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6398 = io_x[9] ? _GEN6397 : _GEN6396;
wire  _GEN6399 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6400 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6401 = io_x[9] ? _GEN6400 : _GEN6399;
wire  _GEN6402 = io_x[24] ? _GEN6401 : _GEN6398;
wire  _GEN6403 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6404 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6405 = io_x[9] ? _GEN6404 : _GEN6403;
wire  _GEN6406 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6407 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6408 = io_x[9] ? _GEN6407 : _GEN6406;
wire  _GEN6409 = io_x[24] ? _GEN6408 : _GEN6405;
wire  _GEN6410 = io_x[26] ? _GEN6409 : _GEN6402;
wire  _GEN6411 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6412 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6413 = io_x[9] ? _GEN6412 : _GEN6411;
wire  _GEN6414 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6415 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6416 = io_x[9] ? _GEN6415 : _GEN6414;
wire  _GEN6417 = io_x[24] ? _GEN6416 : _GEN6413;
wire  _GEN6418 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6419 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6420 = io_x[9] ? _GEN6419 : _GEN6418;
wire  _GEN6421 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6422 = io_x[9] ? _GEN6421 : _GEN6308;
wire  _GEN6423 = io_x[24] ? _GEN6422 : _GEN6420;
wire  _GEN6424 = io_x[26] ? _GEN6423 : _GEN6417;
wire  _GEN6425 = io_x[5] ? _GEN6424 : _GEN6410;
wire  _GEN6426 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6427 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6428 = io_x[9] ? _GEN6427 : _GEN6426;
wire  _GEN6429 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6430 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6431 = io_x[9] ? _GEN6430 : _GEN6429;
wire  _GEN6432 = io_x[24] ? _GEN6431 : _GEN6428;
wire  _GEN6433 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6434 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6435 = io_x[9] ? _GEN6434 : _GEN6433;
wire  _GEN6436 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6437 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6438 = io_x[9] ? _GEN6437 : _GEN6436;
wire  _GEN6439 = io_x[24] ? _GEN6438 : _GEN6435;
wire  _GEN6440 = io_x[26] ? _GEN6439 : _GEN6432;
wire  _GEN6441 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6442 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6443 = io_x[9] ? _GEN6442 : _GEN6441;
wire  _GEN6444 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6445 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6446 = io_x[9] ? _GEN6445 : _GEN6444;
wire  _GEN6447 = io_x[24] ? _GEN6446 : _GEN6443;
wire  _GEN6448 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6449 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6450 = io_x[9] ? _GEN6449 : _GEN6448;
wire  _GEN6451 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6452 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6453 = io_x[9] ? _GEN6452 : _GEN6451;
wire  _GEN6454 = io_x[24] ? _GEN6453 : _GEN6450;
wire  _GEN6455 = io_x[26] ? _GEN6454 : _GEN6447;
wire  _GEN6456 = io_x[5] ? _GEN6455 : _GEN6440;
wire  _GEN6457 = io_x[22] ? _GEN6456 : _GEN6425;
wire  _GEN6458 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6459 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6460 = io_x[9] ? _GEN6459 : _GEN6458;
wire  _GEN6461 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6462 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6463 = io_x[9] ? _GEN6462 : _GEN6461;
wire  _GEN6464 = io_x[24] ? _GEN6463 : _GEN6460;
wire  _GEN6465 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6466 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6467 = io_x[9] ? _GEN6466 : _GEN6465;
wire  _GEN6468 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6469 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6470 = io_x[9] ? _GEN6469 : _GEN6468;
wire  _GEN6471 = io_x[24] ? _GEN6470 : _GEN6467;
wire  _GEN6472 = io_x[26] ? _GEN6471 : _GEN6464;
wire  _GEN6473 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6474 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6475 = io_x[9] ? _GEN6474 : _GEN6473;
wire  _GEN6476 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6477 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6478 = io_x[9] ? _GEN6477 : _GEN6476;
wire  _GEN6479 = io_x[24] ? _GEN6478 : _GEN6475;
wire  _GEN6480 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6481 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6482 = io_x[9] ? _GEN6481 : _GEN6480;
wire  _GEN6483 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6484 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6485 = io_x[9] ? _GEN6484 : _GEN6483;
wire  _GEN6486 = io_x[24] ? _GEN6485 : _GEN6482;
wire  _GEN6487 = io_x[26] ? _GEN6486 : _GEN6479;
wire  _GEN6488 = io_x[5] ? _GEN6487 : _GEN6472;
wire  _GEN6489 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6490 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6491 = io_x[9] ? _GEN6490 : _GEN6489;
wire  _GEN6492 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6493 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6494 = io_x[9] ? _GEN6493 : _GEN6492;
wire  _GEN6495 = io_x[24] ? _GEN6494 : _GEN6491;
wire  _GEN6496 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6497 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6498 = io_x[9] ? _GEN6497 : _GEN6496;
wire  _GEN6499 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6500 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6501 = io_x[9] ? _GEN6500 : _GEN6499;
wire  _GEN6502 = io_x[24] ? _GEN6501 : _GEN6498;
wire  _GEN6503 = io_x[26] ? _GEN6502 : _GEN6495;
wire  _GEN6504 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6505 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6506 = io_x[9] ? _GEN6505 : _GEN6504;
wire  _GEN6507 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6508 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6509 = io_x[9] ? _GEN6508 : _GEN6507;
wire  _GEN6510 = io_x[24] ? _GEN6509 : _GEN6506;
wire  _GEN6511 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6512 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6513 = io_x[9] ? _GEN6512 : _GEN6511;
wire  _GEN6514 = io_x[1] ? _GEN6267 : _GEN6268;
wire  _GEN6515 = io_x[1] ? _GEN6268 : _GEN6267;
wire  _GEN6516 = io_x[9] ? _GEN6515 : _GEN6514;
wire  _GEN6517 = io_x[24] ? _GEN6516 : _GEN6513;
wire  _GEN6518 = io_x[26] ? _GEN6517 : _GEN6510;
wire  _GEN6519 = io_x[5] ? _GEN6518 : _GEN6503;
wire  _GEN6520 = io_x[22] ? _GEN6519 : _GEN6488;
wire  _GEN6521 = io_x[13] ? _GEN6520 : _GEN6457;
wire  _GEN6522 = io_x[30] ? _GEN6521 : _GEN6395;
assign io_y[6] = _GEN6522;
wire  _GEN6523 = 1'b0;
wire  _GEN6524 = 1'b1;
wire  _GEN6525 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6526 = 1'b0;
wire  _GEN6527 = io_x[8] ? _GEN6526 : _GEN6525;
wire  _GEN6528 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6529 = io_x[8] ? _GEN6528 : _GEN6526;
wire  _GEN6530 = io_x[25] ? _GEN6529 : _GEN6527;
wire  _GEN6531 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6532 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6533 = io_x[8] ? _GEN6532 : _GEN6531;
wire  _GEN6534 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6535 = io_x[8] ? _GEN6534 : _GEN6526;
wire  _GEN6536 = io_x[25] ? _GEN6535 : _GEN6533;
wire  _GEN6537 = io_x[3] ? _GEN6536 : _GEN6530;
wire  _GEN6538 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6539 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6540 = io_x[8] ? _GEN6539 : _GEN6538;
wire  _GEN6541 = 1'b1;
wire  _GEN6542 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6543 = io_x[8] ? _GEN6542 : _GEN6541;
wire  _GEN6544 = io_x[25] ? _GEN6543 : _GEN6540;
wire  _GEN6545 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6546 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6547 = io_x[8] ? _GEN6546 : _GEN6545;
wire  _GEN6548 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6549 = io_x[8] ? _GEN6548 : _GEN6541;
wire  _GEN6550 = io_x[25] ? _GEN6549 : _GEN6547;
wire  _GEN6551 = io_x[3] ? _GEN6550 : _GEN6544;
wire  _GEN6552 = io_x[5] ? _GEN6551 : _GEN6537;
wire  _GEN6553 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6554 = io_x[8] ? _GEN6526 : _GEN6553;
wire  _GEN6555 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6556 = io_x[8] ? _GEN6541 : _GEN6555;
wire  _GEN6557 = io_x[25] ? _GEN6556 : _GEN6554;
wire  _GEN6558 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6559 = io_x[8] ? _GEN6558 : _GEN6526;
wire  _GEN6560 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6561 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6562 = io_x[8] ? _GEN6561 : _GEN6560;
wire  _GEN6563 = io_x[25] ? _GEN6562 : _GEN6559;
wire  _GEN6564 = io_x[3] ? _GEN6563 : _GEN6557;
wire  _GEN6565 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6566 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6567 = io_x[8] ? _GEN6566 : _GEN6565;
wire  _GEN6568 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6569 = io_x[8] ? _GEN6526 : _GEN6568;
wire  _GEN6570 = io_x[25] ? _GEN6569 : _GEN6567;
wire  _GEN6571 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6572 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6573 = io_x[8] ? _GEN6572 : _GEN6571;
wire  _GEN6574 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6575 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6576 = io_x[8] ? _GEN6575 : _GEN6574;
wire  _GEN6577 = io_x[25] ? _GEN6576 : _GEN6573;
wire  _GEN6578 = io_x[3] ? _GEN6577 : _GEN6570;
wire  _GEN6579 = io_x[5] ? _GEN6578 : _GEN6564;
wire  _GEN6580 = io_x[7] ? _GEN6579 : _GEN6552;
wire  _GEN6581 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6582 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6583 = io_x[8] ? _GEN6582 : _GEN6581;
wire  _GEN6584 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6585 = io_x[8] ? _GEN6541 : _GEN6584;
wire  _GEN6586 = io_x[25] ? _GEN6585 : _GEN6583;
wire  _GEN6587 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6588 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6589 = io_x[8] ? _GEN6588 : _GEN6587;
wire  _GEN6590 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6591 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6592 = io_x[8] ? _GEN6591 : _GEN6590;
wire  _GEN6593 = io_x[25] ? _GEN6592 : _GEN6589;
wire  _GEN6594 = io_x[3] ? _GEN6593 : _GEN6586;
wire  _GEN6595 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6596 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6597 = io_x[8] ? _GEN6596 : _GEN6595;
wire  _GEN6598 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6599 = io_x[8] ? _GEN6598 : _GEN6541;
wire  _GEN6600 = io_x[25] ? _GEN6599 : _GEN6597;
wire  _GEN6601 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6602 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6603 = io_x[8] ? _GEN6602 : _GEN6601;
wire  _GEN6604 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6605 = io_x[8] ? _GEN6604 : _GEN6541;
wire  _GEN6606 = io_x[25] ? _GEN6605 : _GEN6603;
wire  _GEN6607 = io_x[3] ? _GEN6606 : _GEN6600;
wire  _GEN6608 = io_x[5] ? _GEN6607 : _GEN6594;
wire  _GEN6609 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6610 = io_x[8] ? _GEN6609 : _GEN6526;
wire  _GEN6611 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6612 = io_x[8] ? _GEN6541 : _GEN6611;
wire  _GEN6613 = io_x[25] ? _GEN6612 : _GEN6610;
wire  _GEN6614 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6615 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6616 = io_x[8] ? _GEN6615 : _GEN6614;
wire  _GEN6617 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6618 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6619 = io_x[8] ? _GEN6618 : _GEN6617;
wire  _GEN6620 = io_x[25] ? _GEN6619 : _GEN6616;
wire  _GEN6621 = io_x[3] ? _GEN6620 : _GEN6613;
wire  _GEN6622 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6623 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6624 = io_x[8] ? _GEN6623 : _GEN6622;
wire  _GEN6625 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6626 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6627 = io_x[8] ? _GEN6626 : _GEN6625;
wire  _GEN6628 = io_x[25] ? _GEN6627 : _GEN6624;
wire  _GEN6629 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6630 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6631 = io_x[8] ? _GEN6630 : _GEN6629;
wire  _GEN6632 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6633 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6634 = io_x[8] ? _GEN6633 : _GEN6632;
wire  _GEN6635 = io_x[25] ? _GEN6634 : _GEN6631;
wire  _GEN6636 = io_x[3] ? _GEN6635 : _GEN6628;
wire  _GEN6637 = io_x[5] ? _GEN6636 : _GEN6621;
wire  _GEN6638 = io_x[7] ? _GEN6637 : _GEN6608;
wire  _GEN6639 = io_x[9] ? _GEN6638 : _GEN6580;
wire  _GEN6640 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6641 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6642 = io_x[8] ? _GEN6641 : _GEN6640;
wire  _GEN6643 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6644 = io_x[8] ? _GEN6526 : _GEN6643;
wire  _GEN6645 = io_x[25] ? _GEN6644 : _GEN6642;
wire  _GEN6646 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6647 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6648 = io_x[8] ? _GEN6647 : _GEN6646;
wire  _GEN6649 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6650 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6651 = io_x[8] ? _GEN6650 : _GEN6649;
wire  _GEN6652 = io_x[25] ? _GEN6651 : _GEN6648;
wire  _GEN6653 = io_x[3] ? _GEN6652 : _GEN6645;
wire  _GEN6654 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6655 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6656 = io_x[8] ? _GEN6655 : _GEN6654;
wire  _GEN6657 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6658 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6659 = io_x[8] ? _GEN6658 : _GEN6657;
wire  _GEN6660 = io_x[25] ? _GEN6659 : _GEN6656;
wire  _GEN6661 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6662 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6663 = io_x[8] ? _GEN6662 : _GEN6661;
wire  _GEN6664 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6665 = io_x[8] ? _GEN6664 : _GEN6541;
wire  _GEN6666 = io_x[25] ? _GEN6665 : _GEN6663;
wire  _GEN6667 = io_x[3] ? _GEN6666 : _GEN6660;
wire  _GEN6668 = io_x[5] ? _GEN6667 : _GEN6653;
wire  _GEN6669 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6670 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6671 = io_x[8] ? _GEN6670 : _GEN6669;
wire  _GEN6672 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6673 = io_x[8] ? _GEN6526 : _GEN6672;
wire  _GEN6674 = io_x[25] ? _GEN6673 : _GEN6671;
wire  _GEN6675 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6676 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6677 = io_x[8] ? _GEN6676 : _GEN6675;
wire  _GEN6678 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6679 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6680 = io_x[8] ? _GEN6679 : _GEN6678;
wire  _GEN6681 = io_x[25] ? _GEN6680 : _GEN6677;
wire  _GEN6682 = io_x[3] ? _GEN6681 : _GEN6674;
wire  _GEN6683 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6684 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6685 = io_x[8] ? _GEN6684 : _GEN6683;
wire  _GEN6686 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6687 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6688 = io_x[8] ? _GEN6687 : _GEN6686;
wire  _GEN6689 = io_x[25] ? _GEN6688 : _GEN6685;
wire  _GEN6690 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6691 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6692 = io_x[8] ? _GEN6691 : _GEN6690;
wire  _GEN6693 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6694 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6695 = io_x[8] ? _GEN6694 : _GEN6693;
wire  _GEN6696 = io_x[25] ? _GEN6695 : _GEN6692;
wire  _GEN6697 = io_x[3] ? _GEN6696 : _GEN6689;
wire  _GEN6698 = io_x[5] ? _GEN6697 : _GEN6682;
wire  _GEN6699 = io_x[7] ? _GEN6698 : _GEN6668;
wire  _GEN6700 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6701 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6702 = io_x[8] ? _GEN6701 : _GEN6700;
wire  _GEN6703 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6704 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6705 = io_x[8] ? _GEN6704 : _GEN6703;
wire  _GEN6706 = io_x[25] ? _GEN6705 : _GEN6702;
wire  _GEN6707 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6708 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6709 = io_x[8] ? _GEN6708 : _GEN6707;
wire  _GEN6710 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6711 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6712 = io_x[8] ? _GEN6711 : _GEN6710;
wire  _GEN6713 = io_x[25] ? _GEN6712 : _GEN6709;
wire  _GEN6714 = io_x[3] ? _GEN6713 : _GEN6706;
wire  _GEN6715 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6716 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6717 = io_x[8] ? _GEN6716 : _GEN6715;
wire  _GEN6718 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6719 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6720 = io_x[8] ? _GEN6719 : _GEN6718;
wire  _GEN6721 = io_x[25] ? _GEN6720 : _GEN6717;
wire  _GEN6722 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6723 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6724 = io_x[8] ? _GEN6723 : _GEN6722;
wire  _GEN6725 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6726 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6727 = io_x[8] ? _GEN6726 : _GEN6725;
wire  _GEN6728 = io_x[25] ? _GEN6727 : _GEN6724;
wire  _GEN6729 = io_x[3] ? _GEN6728 : _GEN6721;
wire  _GEN6730 = io_x[5] ? _GEN6729 : _GEN6714;
wire  _GEN6731 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6732 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6733 = io_x[8] ? _GEN6732 : _GEN6731;
wire  _GEN6734 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6735 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6736 = io_x[8] ? _GEN6735 : _GEN6734;
wire  _GEN6737 = io_x[25] ? _GEN6736 : _GEN6733;
wire  _GEN6738 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6739 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6740 = io_x[8] ? _GEN6739 : _GEN6738;
wire  _GEN6741 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6742 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6743 = io_x[8] ? _GEN6742 : _GEN6741;
wire  _GEN6744 = io_x[25] ? _GEN6743 : _GEN6740;
wire  _GEN6745 = io_x[3] ? _GEN6744 : _GEN6737;
wire  _GEN6746 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6747 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6748 = io_x[8] ? _GEN6747 : _GEN6746;
wire  _GEN6749 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6750 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6751 = io_x[8] ? _GEN6750 : _GEN6749;
wire  _GEN6752 = io_x[25] ? _GEN6751 : _GEN6748;
wire  _GEN6753 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6754 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6755 = io_x[8] ? _GEN6754 : _GEN6753;
wire  _GEN6756 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6757 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6758 = io_x[8] ? _GEN6757 : _GEN6756;
wire  _GEN6759 = io_x[25] ? _GEN6758 : _GEN6755;
wire  _GEN6760 = io_x[3] ? _GEN6759 : _GEN6752;
wire  _GEN6761 = io_x[5] ? _GEN6760 : _GEN6745;
wire  _GEN6762 = io_x[7] ? _GEN6761 : _GEN6730;
wire  _GEN6763 = io_x[9] ? _GEN6762 : _GEN6699;
wire  _GEN6764 = io_x[0] ? _GEN6763 : _GEN6639;
wire  _GEN6765 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6766 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6767 = io_x[8] ? _GEN6766 : _GEN6765;
wire  _GEN6768 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6769 = io_x[8] ? _GEN6768 : _GEN6541;
wire  _GEN6770 = io_x[25] ? _GEN6769 : _GEN6767;
wire  _GEN6771 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6772 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6773 = io_x[8] ? _GEN6772 : _GEN6771;
wire  _GEN6774 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6775 = io_x[8] ? _GEN6774 : _GEN6541;
wire  _GEN6776 = io_x[25] ? _GEN6775 : _GEN6773;
wire  _GEN6777 = io_x[3] ? _GEN6776 : _GEN6770;
wire  _GEN6778 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6779 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6780 = io_x[8] ? _GEN6779 : _GEN6778;
wire  _GEN6781 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6782 = io_x[8] ? _GEN6781 : _GEN6541;
wire  _GEN6783 = io_x[25] ? _GEN6782 : _GEN6780;
wire  _GEN6784 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6785 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6786 = io_x[8] ? _GEN6785 : _GEN6784;
wire  _GEN6787 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6788 = io_x[8] ? _GEN6787 : _GEN6541;
wire  _GEN6789 = io_x[25] ? _GEN6788 : _GEN6786;
wire  _GEN6790 = io_x[3] ? _GEN6789 : _GEN6783;
wire  _GEN6791 = io_x[5] ? _GEN6790 : _GEN6777;
wire  _GEN6792 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6793 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6794 = io_x[8] ? _GEN6793 : _GEN6792;
wire  _GEN6795 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6796 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6797 = io_x[8] ? _GEN6796 : _GEN6795;
wire  _GEN6798 = io_x[25] ? _GEN6797 : _GEN6794;
wire  _GEN6799 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6800 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6801 = io_x[8] ? _GEN6800 : _GEN6799;
wire  _GEN6802 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6803 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6804 = io_x[8] ? _GEN6803 : _GEN6802;
wire  _GEN6805 = io_x[25] ? _GEN6804 : _GEN6801;
wire  _GEN6806 = io_x[3] ? _GEN6805 : _GEN6798;
wire  _GEN6807 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6808 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6809 = io_x[8] ? _GEN6808 : _GEN6807;
wire  _GEN6810 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6811 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6812 = io_x[8] ? _GEN6811 : _GEN6810;
wire  _GEN6813 = io_x[25] ? _GEN6812 : _GEN6809;
wire  _GEN6814 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6815 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6816 = io_x[8] ? _GEN6815 : _GEN6814;
wire  _GEN6817 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6818 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6819 = io_x[8] ? _GEN6818 : _GEN6817;
wire  _GEN6820 = io_x[25] ? _GEN6819 : _GEN6816;
wire  _GEN6821 = io_x[3] ? _GEN6820 : _GEN6813;
wire  _GEN6822 = io_x[5] ? _GEN6821 : _GEN6806;
wire  _GEN6823 = io_x[7] ? _GEN6822 : _GEN6791;
wire  _GEN6824 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6825 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6826 = io_x[8] ? _GEN6825 : _GEN6824;
wire  _GEN6827 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6828 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6829 = io_x[8] ? _GEN6828 : _GEN6827;
wire  _GEN6830 = io_x[25] ? _GEN6829 : _GEN6826;
wire  _GEN6831 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6832 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6833 = io_x[8] ? _GEN6832 : _GEN6831;
wire  _GEN6834 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6835 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6836 = io_x[8] ? _GEN6835 : _GEN6834;
wire  _GEN6837 = io_x[25] ? _GEN6836 : _GEN6833;
wire  _GEN6838 = io_x[3] ? _GEN6837 : _GEN6830;
wire  _GEN6839 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6840 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6841 = io_x[8] ? _GEN6840 : _GEN6839;
wire  _GEN6842 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6843 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6844 = io_x[8] ? _GEN6843 : _GEN6842;
wire  _GEN6845 = io_x[25] ? _GEN6844 : _GEN6841;
wire  _GEN6846 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6847 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6848 = io_x[8] ? _GEN6847 : _GEN6846;
wire  _GEN6849 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6850 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6851 = io_x[8] ? _GEN6850 : _GEN6849;
wire  _GEN6852 = io_x[25] ? _GEN6851 : _GEN6848;
wire  _GEN6853 = io_x[3] ? _GEN6852 : _GEN6845;
wire  _GEN6854 = io_x[5] ? _GEN6853 : _GEN6838;
wire  _GEN6855 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6856 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6857 = io_x[8] ? _GEN6856 : _GEN6855;
wire  _GEN6858 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6859 = io_x[8] ? _GEN6858 : _GEN6541;
wire  _GEN6860 = io_x[25] ? _GEN6859 : _GEN6857;
wire  _GEN6861 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6862 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6863 = io_x[8] ? _GEN6862 : _GEN6861;
wire  _GEN6864 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6865 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6866 = io_x[8] ? _GEN6865 : _GEN6864;
wire  _GEN6867 = io_x[25] ? _GEN6866 : _GEN6863;
wire  _GEN6868 = io_x[3] ? _GEN6867 : _GEN6860;
wire  _GEN6869 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6870 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6871 = io_x[8] ? _GEN6870 : _GEN6869;
wire  _GEN6872 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6873 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6874 = io_x[8] ? _GEN6873 : _GEN6872;
wire  _GEN6875 = io_x[25] ? _GEN6874 : _GEN6871;
wire  _GEN6876 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6877 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6878 = io_x[8] ? _GEN6877 : _GEN6876;
wire  _GEN6879 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6880 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6881 = io_x[8] ? _GEN6880 : _GEN6879;
wire  _GEN6882 = io_x[25] ? _GEN6881 : _GEN6878;
wire  _GEN6883 = io_x[3] ? _GEN6882 : _GEN6875;
wire  _GEN6884 = io_x[5] ? _GEN6883 : _GEN6868;
wire  _GEN6885 = io_x[7] ? _GEN6884 : _GEN6854;
wire  _GEN6886 = io_x[9] ? _GEN6885 : _GEN6823;
wire  _GEN6887 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6888 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6889 = io_x[8] ? _GEN6888 : _GEN6887;
wire  _GEN6890 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6891 = io_x[8] ? _GEN6890 : _GEN6526;
wire  _GEN6892 = io_x[25] ? _GEN6891 : _GEN6889;
wire  _GEN6893 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6894 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6895 = io_x[8] ? _GEN6894 : _GEN6893;
wire  _GEN6896 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6897 = io_x[8] ? _GEN6896 : _GEN6541;
wire  _GEN6898 = io_x[25] ? _GEN6897 : _GEN6895;
wire  _GEN6899 = io_x[3] ? _GEN6898 : _GEN6892;
wire  _GEN6900 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6901 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6902 = io_x[8] ? _GEN6901 : _GEN6900;
wire  _GEN6903 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6904 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6905 = io_x[8] ? _GEN6904 : _GEN6903;
wire  _GEN6906 = io_x[25] ? _GEN6905 : _GEN6902;
wire  _GEN6907 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6908 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6909 = io_x[8] ? _GEN6908 : _GEN6907;
wire  _GEN6910 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6911 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6912 = io_x[8] ? _GEN6911 : _GEN6910;
wire  _GEN6913 = io_x[25] ? _GEN6912 : _GEN6909;
wire  _GEN6914 = io_x[3] ? _GEN6913 : _GEN6906;
wire  _GEN6915 = io_x[5] ? _GEN6914 : _GEN6899;
wire  _GEN6916 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6917 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6918 = io_x[8] ? _GEN6917 : _GEN6916;
wire  _GEN6919 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6920 = io_x[8] ? _GEN6541 : _GEN6919;
wire  _GEN6921 = io_x[25] ? _GEN6920 : _GEN6918;
wire  _GEN6922 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6923 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6924 = io_x[8] ? _GEN6923 : _GEN6922;
wire  _GEN6925 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6926 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6927 = io_x[8] ? _GEN6926 : _GEN6925;
wire  _GEN6928 = io_x[25] ? _GEN6927 : _GEN6924;
wire  _GEN6929 = io_x[3] ? _GEN6928 : _GEN6921;
wire  _GEN6930 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6931 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6932 = io_x[8] ? _GEN6931 : _GEN6930;
wire  _GEN6933 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6934 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6935 = io_x[8] ? _GEN6934 : _GEN6933;
wire  _GEN6936 = io_x[25] ? _GEN6935 : _GEN6932;
wire  _GEN6937 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6938 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6939 = io_x[8] ? _GEN6938 : _GEN6937;
wire  _GEN6940 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6941 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6942 = io_x[8] ? _GEN6941 : _GEN6940;
wire  _GEN6943 = io_x[25] ? _GEN6942 : _GEN6939;
wire  _GEN6944 = io_x[3] ? _GEN6943 : _GEN6936;
wire  _GEN6945 = io_x[5] ? _GEN6944 : _GEN6929;
wire  _GEN6946 = io_x[7] ? _GEN6945 : _GEN6915;
wire  _GEN6947 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6948 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6949 = io_x[8] ? _GEN6948 : _GEN6947;
wire  _GEN6950 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6951 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6952 = io_x[8] ? _GEN6951 : _GEN6950;
wire  _GEN6953 = io_x[25] ? _GEN6952 : _GEN6949;
wire  _GEN6954 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6955 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6956 = io_x[8] ? _GEN6955 : _GEN6954;
wire  _GEN6957 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6958 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6959 = io_x[8] ? _GEN6958 : _GEN6957;
wire  _GEN6960 = io_x[25] ? _GEN6959 : _GEN6956;
wire  _GEN6961 = io_x[3] ? _GEN6960 : _GEN6953;
wire  _GEN6962 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6963 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6964 = io_x[8] ? _GEN6963 : _GEN6962;
wire  _GEN6965 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6966 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6967 = io_x[8] ? _GEN6966 : _GEN6965;
wire  _GEN6968 = io_x[25] ? _GEN6967 : _GEN6964;
wire  _GEN6969 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6970 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6971 = io_x[8] ? _GEN6970 : _GEN6969;
wire  _GEN6972 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6973 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6974 = io_x[8] ? _GEN6973 : _GEN6972;
wire  _GEN6975 = io_x[25] ? _GEN6974 : _GEN6971;
wire  _GEN6976 = io_x[3] ? _GEN6975 : _GEN6968;
wire  _GEN6977 = io_x[5] ? _GEN6976 : _GEN6961;
wire  _GEN6978 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6979 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6980 = io_x[8] ? _GEN6979 : _GEN6978;
wire  _GEN6981 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6982 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6983 = io_x[8] ? _GEN6982 : _GEN6981;
wire  _GEN6984 = io_x[25] ? _GEN6983 : _GEN6980;
wire  _GEN6985 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6986 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6987 = io_x[8] ? _GEN6986 : _GEN6985;
wire  _GEN6988 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6989 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6990 = io_x[8] ? _GEN6989 : _GEN6988;
wire  _GEN6991 = io_x[25] ? _GEN6990 : _GEN6987;
wire  _GEN6992 = io_x[3] ? _GEN6991 : _GEN6984;
wire  _GEN6993 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6994 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6995 = io_x[8] ? _GEN6994 : _GEN6993;
wire  _GEN6996 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN6997 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN6998 = io_x[8] ? _GEN6997 : _GEN6996;
wire  _GEN6999 = io_x[25] ? _GEN6998 : _GEN6995;
wire  _GEN7000 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN7001 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN7002 = io_x[8] ? _GEN7001 : _GEN7000;
wire  _GEN7003 = io_x[4] ? _GEN6523 : _GEN6524;
wire  _GEN7004 = io_x[4] ? _GEN6524 : _GEN6523;
wire  _GEN7005 = io_x[8] ? _GEN7004 : _GEN7003;
wire  _GEN7006 = io_x[25] ? _GEN7005 : _GEN7002;
wire  _GEN7007 = io_x[3] ? _GEN7006 : _GEN6999;
wire  _GEN7008 = io_x[5] ? _GEN7007 : _GEN6992;
wire  _GEN7009 = io_x[7] ? _GEN7008 : _GEN6977;
wire  _GEN7010 = io_x[9] ? _GEN7009 : _GEN6946;
wire  _GEN7011 = io_x[0] ? _GEN7010 : _GEN6886;
wire  _GEN7012 = io_x[12] ? _GEN7011 : _GEN6764;
assign io_y[5] = _GEN7012;
wire  _GEN7013 = 1'b0;
wire  _GEN7014 = 1'b1;
wire  _GEN7015 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7016 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7017 = io_x[22] ? _GEN7016 : _GEN7015;
wire  _GEN7018 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7019 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7020 = io_x[22] ? _GEN7019 : _GEN7018;
wire  _GEN7021 = io_x[28] ? _GEN7020 : _GEN7017;
wire  _GEN7022 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7023 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7024 = io_x[22] ? _GEN7023 : _GEN7022;
wire  _GEN7025 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7026 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7027 = io_x[22] ? _GEN7026 : _GEN7025;
wire  _GEN7028 = io_x[28] ? _GEN7027 : _GEN7024;
wire  _GEN7029 = io_x[17] ? _GEN7028 : _GEN7021;
wire  _GEN7030 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7031 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7032 = io_x[22] ? _GEN7031 : _GEN7030;
wire  _GEN7033 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7034 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7035 = io_x[22] ? _GEN7034 : _GEN7033;
wire  _GEN7036 = io_x[28] ? _GEN7035 : _GEN7032;
wire  _GEN7037 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7038 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7039 = io_x[22] ? _GEN7038 : _GEN7037;
wire  _GEN7040 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7041 = io_x[24] ? _GEN7014 : _GEN7013;
wire  _GEN7042 = io_x[22] ? _GEN7041 : _GEN7040;
wire  _GEN7043 = io_x[28] ? _GEN7042 : _GEN7039;
wire  _GEN7044 = io_x[17] ? _GEN7043 : _GEN7036;
wire  _GEN7045 = io_x[23] ? _GEN7044 : _GEN7029;
assign io_y[4] = _GEN7045;
wire  _GEN7046 = 1'b0;
wire  _GEN7047 = 1'b1;
wire  _GEN7048 = io_x[23] ? _GEN7047 : _GEN7046;
wire  _GEN7049 = io_x[23] ? _GEN7047 : _GEN7046;
wire  _GEN7050 = io_x[16] ? _GEN7049 : _GEN7048;
assign io_y[3] = _GEN7050;
wire  _GEN7051 = 1'b0;
wire  _GEN7052 = 1'b1;
wire  _GEN7053 = io_x[22] ? _GEN7052 : _GEN7051;
assign io_y[2] = _GEN7053;
wire  _GEN7054 = 1'b0;
wire  _GEN7055 = 1'b1;
wire  _GEN7056 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7057 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7058 = io_x[22] ? _GEN7057 : _GEN7056;
wire  _GEN7059 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7060 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7061 = io_x[22] ? _GEN7060 : _GEN7059;
wire  _GEN7062 = io_x[5] ? _GEN7061 : _GEN7058;
wire  _GEN7063 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7064 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7065 = io_x[22] ? _GEN7064 : _GEN7063;
wire  _GEN7066 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7067 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7068 = io_x[22] ? _GEN7067 : _GEN7066;
wire  _GEN7069 = io_x[5] ? _GEN7068 : _GEN7065;
wire  _GEN7070 = io_x[3] ? _GEN7069 : _GEN7062;
wire  _GEN7071 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7072 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7073 = io_x[22] ? _GEN7072 : _GEN7071;
wire  _GEN7074 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7075 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7076 = io_x[22] ? _GEN7075 : _GEN7074;
wire  _GEN7077 = io_x[5] ? _GEN7076 : _GEN7073;
wire  _GEN7078 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7079 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7080 = io_x[22] ? _GEN7079 : _GEN7078;
wire  _GEN7081 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7082 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7083 = io_x[22] ? _GEN7082 : _GEN7081;
wire  _GEN7084 = io_x[5] ? _GEN7083 : _GEN7080;
wire  _GEN7085 = io_x[3] ? _GEN7084 : _GEN7077;
wire  _GEN7086 = io_x[30] ? _GEN7085 : _GEN7070;
wire  _GEN7087 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7088 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7089 = io_x[22] ? _GEN7088 : _GEN7087;
wire  _GEN7090 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7091 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7092 = io_x[22] ? _GEN7091 : _GEN7090;
wire  _GEN7093 = io_x[5] ? _GEN7092 : _GEN7089;
wire  _GEN7094 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7095 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7096 = io_x[22] ? _GEN7095 : _GEN7094;
wire  _GEN7097 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7098 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7099 = io_x[22] ? _GEN7098 : _GEN7097;
wire  _GEN7100 = io_x[5] ? _GEN7099 : _GEN7096;
wire  _GEN7101 = io_x[3] ? _GEN7100 : _GEN7093;
wire  _GEN7102 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7103 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7104 = io_x[22] ? _GEN7103 : _GEN7102;
wire  _GEN7105 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7106 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7107 = io_x[22] ? _GEN7106 : _GEN7105;
wire  _GEN7108 = io_x[5] ? _GEN7107 : _GEN7104;
wire  _GEN7109 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7110 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7111 = io_x[22] ? _GEN7110 : _GEN7109;
wire  _GEN7112 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7113 = io_x[21] ? _GEN7055 : _GEN7054;
wire  _GEN7114 = io_x[22] ? _GEN7113 : _GEN7112;
wire  _GEN7115 = io_x[5] ? _GEN7114 : _GEN7111;
wire  _GEN7116 = io_x[3] ? _GEN7115 : _GEN7108;
wire  _GEN7117 = io_x[30] ? _GEN7116 : _GEN7101;
wire  _GEN7118 = io_x[17] ? _GEN7117 : _GEN7086;
assign io_y[1] = _GEN7118;
wire  _GEN7119 = 1'b0;
wire  _GEN7120 = 1'b1;
wire  _GEN7121 = io_x[20] ? _GEN7120 : _GEN7119;
wire  _GEN7122 = io_x[20] ? _GEN7120 : _GEN7119;
wire  _GEN7123 = io_x[1] ? _GEN7122 : _GEN7121;
wire  _GEN7124 = io_x[20] ? _GEN7120 : _GEN7119;
wire  _GEN7125 = io_x[20] ? _GEN7120 : _GEN7119;
wire  _GEN7126 = io_x[1] ? _GEN7125 : _GEN7124;
wire  _GEN7127 = io_x[22] ? _GEN7126 : _GEN7123;
wire  _GEN7128 = io_x[20] ? _GEN7120 : _GEN7119;
wire  _GEN7129 = io_x[20] ? _GEN7120 : _GEN7119;
wire  _GEN7130 = io_x[1] ? _GEN7129 : _GEN7128;
wire  _GEN7131 = io_x[20] ? _GEN7120 : _GEN7119;
wire  _GEN7132 = io_x[20] ? _GEN7120 : _GEN7119;
wire  _GEN7133 = io_x[1] ? _GEN7132 : _GEN7131;
wire  _GEN7134 = io_x[22] ? _GEN7133 : _GEN7130;
wire  _GEN7135 = io_x[30] ? _GEN7134 : _GEN7127;
assign io_y[0] = _GEN7135;
endmodule
module sim_GShare_train(
    input [31:0] train_pc,
    input  train_taken,
    input [15:0] train_ghr_rdata,
    output  pht_wdata,
    output [8:0] pht_waddr,
    output  ghr_wdata
);
wire [48:0] io_x;
wire [10:0] io_y;
assign io_x = { train_pc, train_taken, train_ghr_rdata };
assign { pht_wdata, pht_waddr, ghr_wdata } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN3 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN4 = io_x[6] ? _GEN3 : _GEN2;
wire  _GEN5 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN6 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN7 = io_x[6] ? _GEN6 : _GEN5;
wire  _GEN8 = io_x[2] ? _GEN7 : _GEN4;
wire  _GEN9 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN10 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN11 = io_x[6] ? _GEN10 : _GEN9;
wire  _GEN12 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN13 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN14 = io_x[6] ? _GEN13 : _GEN12;
wire  _GEN15 = io_x[2] ? _GEN14 : _GEN11;
wire  _GEN16 = io_x[30] ? _GEN15 : _GEN8;
wire  _GEN17 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN18 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN19 = io_x[6] ? _GEN18 : _GEN17;
wire  _GEN20 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN21 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN22 = io_x[6] ? _GEN21 : _GEN20;
wire  _GEN23 = io_x[2] ? _GEN22 : _GEN19;
wire  _GEN24 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN25 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN26 = io_x[6] ? _GEN25 : _GEN24;
wire  _GEN27 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN28 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN29 = io_x[6] ? _GEN28 : _GEN27;
wire  _GEN30 = io_x[2] ? _GEN29 : _GEN26;
wire  _GEN31 = io_x[30] ? _GEN30 : _GEN23;
wire  _GEN32 = io_x[4] ? _GEN31 : _GEN16;
wire  _GEN33 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN34 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN35 = io_x[6] ? _GEN34 : _GEN33;
wire  _GEN36 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN37 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN38 = io_x[6] ? _GEN37 : _GEN36;
wire  _GEN39 = io_x[2] ? _GEN38 : _GEN35;
wire  _GEN40 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN41 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN42 = io_x[6] ? _GEN41 : _GEN40;
wire  _GEN43 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN44 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN45 = io_x[6] ? _GEN44 : _GEN43;
wire  _GEN46 = io_x[2] ? _GEN45 : _GEN42;
wire  _GEN47 = io_x[30] ? _GEN46 : _GEN39;
wire  _GEN48 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN49 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN50 = io_x[6] ? _GEN49 : _GEN48;
wire  _GEN51 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN52 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN53 = io_x[6] ? _GEN52 : _GEN51;
wire  _GEN54 = io_x[2] ? _GEN53 : _GEN50;
wire  _GEN55 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN56 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN57 = io_x[6] ? _GEN56 : _GEN55;
wire  _GEN58 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN59 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN60 = io_x[6] ? _GEN59 : _GEN58;
wire  _GEN61 = io_x[2] ? _GEN60 : _GEN57;
wire  _GEN62 = io_x[30] ? _GEN61 : _GEN54;
wire  _GEN63 = io_x[4] ? _GEN62 : _GEN47;
wire  _GEN64 = io_x[0] ? _GEN63 : _GEN32;
assign io_y[10] = _GEN64;
wire  _GEN65 = 1'b1;
wire  _GEN66 = 1'b1;
wire  _GEN67 = 1'b1;
wire  _GEN68 = 1'b1;
wire  _GEN69 = 1'b0;
wire  _GEN70 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN71 = io_x[11] ? _GEN70 : _GEN67;
wire  _GEN72 = io_x[3] ? _GEN71 : _GEN66;
wire  _GEN73 = io_x[7] ? _GEN72 : _GEN65;
wire  _GEN74 = 1'b0;
wire  _GEN75 = io_x[23] ? _GEN74 : _GEN73;
wire  _GEN76 = 1'b0;
wire  _GEN77 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN78 = 1'b0;
wire  _GEN79 = io_x[3] ? _GEN78 : _GEN77;
wire  _GEN80 = io_x[7] ? _GEN79 : _GEN65;
wire  _GEN81 = 1'b1;
wire  _GEN82 = io_x[23] ? _GEN81 : _GEN80;
wire  _GEN83 = io_x[2] ? _GEN82 : _GEN75;
wire  _GEN84 = 1'b0;
wire  _GEN85 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN86 = io_x[23] ? _GEN85 : _GEN74;
wire  _GEN87 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN88 = io_x[11] ? _GEN76 : _GEN87;
wire  _GEN89 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN90 = io_x[3] ? _GEN89 : _GEN88;
wire  _GEN91 = io_x[7] ? _GEN90 : _GEN65;
wire  _GEN92 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN93 = io_x[3] ? _GEN78 : _GEN92;
wire  _GEN94 = io_x[7] ? _GEN93 : _GEN84;
wire  _GEN95 = io_x[23] ? _GEN94 : _GEN91;
wire  _GEN96 = io_x[2] ? _GEN95 : _GEN86;
wire  _GEN97 = io_x[16] ? _GEN96 : _GEN83;
wire  _GEN98 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN99 = io_x[11] ? _GEN98 : _GEN67;
wire  _GEN100 = io_x[3] ? _GEN66 : _GEN99;
wire  _GEN101 = io_x[7] ? _GEN100 : _GEN65;
wire  _GEN102 = io_x[23] ? _GEN81 : _GEN101;
wire  _GEN103 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN104 = io_x[3] ? _GEN66 : _GEN103;
wire  _GEN105 = io_x[7] ? _GEN104 : _GEN65;
wire  _GEN106 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN107 = io_x[3] ? _GEN66 : _GEN106;
wire  _GEN108 = io_x[7] ? _GEN84 : _GEN107;
wire  _GEN109 = io_x[23] ? _GEN108 : _GEN105;
wire  _GEN110 = io_x[2] ? _GEN109 : _GEN102;
wire  _GEN111 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN112 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN113 = io_x[11] ? _GEN112 : _GEN67;
wire  _GEN114 = io_x[3] ? _GEN113 : _GEN66;
wire  _GEN115 = io_x[7] ? _GEN114 : _GEN65;
wire  _GEN116 = io_x[23] ? _GEN115 : _GEN111;
wire  _GEN117 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN118 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN119 = io_x[11] ? _GEN118 : _GEN76;
wire  _GEN120 = io_x[3] ? _GEN119 : _GEN66;
wire  _GEN121 = io_x[7] ? _GEN120 : _GEN117;
wire  _GEN122 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN123 = io_x[11] ? _GEN122 : _GEN67;
wire  _GEN124 = io_x[3] ? _GEN66 : _GEN123;
wire  _GEN125 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN126 = io_x[3] ? _GEN66 : _GEN125;
wire  _GEN127 = io_x[7] ? _GEN126 : _GEN124;
wire  _GEN128 = io_x[23] ? _GEN127 : _GEN121;
wire  _GEN129 = io_x[2] ? _GEN128 : _GEN116;
wire  _GEN130 = io_x[16] ? _GEN129 : _GEN110;
wire  _GEN131 = io_x[15] ? _GEN130 : _GEN97;
wire  _GEN132 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN133 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN134 = io_x[23] ? _GEN133 : _GEN132;
wire  _GEN135 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN136 = io_x[3] ? _GEN66 : _GEN135;
wire  _GEN137 = io_x[7] ? _GEN136 : _GEN84;
wire  _GEN138 = io_x[23] ? _GEN137 : _GEN74;
wire  _GEN139 = io_x[2] ? _GEN138 : _GEN134;
wire  _GEN140 = 1'b0;
wire  _GEN141 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN142 = io_x[11] ? _GEN141 : _GEN67;
wire  _GEN143 = io_x[3] ? _GEN142 : _GEN66;
wire  _GEN144 = io_x[7] ? _GEN143 : _GEN84;
wire  _GEN145 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN146 = io_x[7] ? _GEN145 : _GEN84;
wire  _GEN147 = io_x[23] ? _GEN146 : _GEN144;
wire  _GEN148 = io_x[2] ? _GEN147 : _GEN140;
wire  _GEN149 = io_x[16] ? _GEN148 : _GEN139;
wire  _GEN150 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN151 = io_x[11] ? _GEN67 : _GEN150;
wire  _GEN152 = io_x[3] ? _GEN151 : _GEN66;
wire  _GEN153 = io_x[7] ? _GEN152 : _GEN65;
wire  _GEN154 = io_x[23] ? _GEN81 : _GEN153;
wire  _GEN155 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN156 = io_x[7] ? _GEN65 : _GEN155;
wire  _GEN157 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN158 = io_x[3] ? _GEN66 : _GEN157;
wire  _GEN159 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN160 = io_x[3] ? _GEN66 : _GEN159;
wire  _GEN161 = io_x[7] ? _GEN160 : _GEN158;
wire  _GEN162 = io_x[23] ? _GEN161 : _GEN156;
wire  _GEN163 = io_x[2] ? _GEN162 : _GEN154;
wire  _GEN164 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN165 = io_x[23] ? _GEN81 : _GEN164;
wire  _GEN166 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN167 = io_x[11] ? _GEN166 : _GEN67;
wire  _GEN168 = io_x[3] ? _GEN78 : _GEN167;
wire  _GEN169 = io_x[7] ? _GEN168 : _GEN65;
wire  _GEN170 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN171 = io_x[3] ? _GEN170 : _GEN66;
wire  _GEN172 = io_x[7] ? _GEN171 : _GEN65;
wire  _GEN173 = io_x[23] ? _GEN172 : _GEN169;
wire  _GEN174 = io_x[2] ? _GEN173 : _GEN165;
wire  _GEN175 = io_x[16] ? _GEN174 : _GEN163;
wire  _GEN176 = io_x[15] ? _GEN175 : _GEN149;
wire  _GEN177 = io_x[12] ? _GEN176 : _GEN131;
wire  _GEN178 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN179 = io_x[23] ? _GEN81 : _GEN74;
wire  _GEN180 = io_x[2] ? _GEN179 : _GEN178;
wire  _GEN181 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN182 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN183 = io_x[3] ? _GEN182 : _GEN66;
wire  _GEN184 = io_x[7] ? _GEN183 : _GEN84;
wire  _GEN185 = io_x[23] ? _GEN184 : _GEN181;
wire  _GEN186 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN187 = io_x[3] ? _GEN186 : _GEN66;
wire  _GEN188 = io_x[7] ? _GEN187 : _GEN65;
wire  _GEN189 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN190 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN191 = io_x[7] ? _GEN190 : _GEN189;
wire  _GEN192 = io_x[23] ? _GEN191 : _GEN188;
wire  _GEN193 = io_x[2] ? _GEN192 : _GEN185;
wire  _GEN194 = io_x[16] ? _GEN193 : _GEN180;
wire  _GEN195 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN196 = io_x[11] ? _GEN195 : _GEN76;
wire  _GEN197 = io_x[3] ? _GEN196 : _GEN66;
wire  _GEN198 = io_x[7] ? _GEN197 : _GEN65;
wire  _GEN199 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN200 = io_x[3] ? _GEN66 : _GEN199;
wire  _GEN201 = io_x[7] ? _GEN84 : _GEN200;
wire  _GEN202 = io_x[23] ? _GEN201 : _GEN198;
wire  _GEN203 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN204 = io_x[3] ? _GEN203 : _GEN66;
wire  _GEN205 = io_x[7] ? _GEN204 : _GEN84;
wire  _GEN206 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN207 = io_x[7] ? _GEN206 : _GEN65;
wire  _GEN208 = io_x[23] ? _GEN207 : _GEN205;
wire  _GEN209 = io_x[2] ? _GEN208 : _GEN202;
wire  _GEN210 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN211 = io_x[11] ? _GEN67 : _GEN210;
wire  _GEN212 = io_x[3] ? _GEN78 : _GEN211;
wire  _GEN213 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN214 = io_x[3] ? _GEN213 : _GEN66;
wire  _GEN215 = io_x[7] ? _GEN214 : _GEN212;
wire  _GEN216 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN217 = io_x[3] ? _GEN216 : _GEN66;
wire  _GEN218 = io_x[7] ? _GEN217 : _GEN65;
wire  _GEN219 = io_x[23] ? _GEN218 : _GEN215;
wire  _GEN220 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN221 = io_x[11] ? _GEN220 : _GEN76;
wire  _GEN222 = io_x[3] ? _GEN221 : _GEN66;
wire  _GEN223 = io_x[7] ? _GEN222 : _GEN65;
wire  _GEN224 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN225 = io_x[3] ? _GEN224 : _GEN66;
wire  _GEN226 = io_x[7] ? _GEN225 : _GEN65;
wire  _GEN227 = io_x[23] ? _GEN226 : _GEN223;
wire  _GEN228 = io_x[2] ? _GEN227 : _GEN219;
wire  _GEN229 = io_x[16] ? _GEN228 : _GEN209;
wire  _GEN230 = io_x[15] ? _GEN229 : _GEN194;
wire  _GEN231 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN232 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN233 = io_x[11] ? _GEN76 : _GEN232;
wire  _GEN234 = io_x[3] ? _GEN233 : _GEN66;
wire  _GEN235 = io_x[7] ? _GEN234 : _GEN231;
wire  _GEN236 = io_x[23] ? _GEN74 : _GEN235;
wire  _GEN237 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN238 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN239 = io_x[3] ? _GEN66 : _GEN238;
wire  _GEN240 = io_x[7] ? _GEN239 : _GEN65;
wire  _GEN241 = io_x[23] ? _GEN240 : _GEN237;
wire  _GEN242 = io_x[2] ? _GEN241 : _GEN236;
wire  _GEN243 = io_x[23] ? _GEN81 : _GEN74;
wire  _GEN244 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN245 = io_x[11] ? _GEN67 : _GEN244;
wire  _GEN246 = io_x[3] ? _GEN245 : _GEN78;
wire  _GEN247 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN248 = io_x[11] ? _GEN247 : _GEN67;
wire  _GEN249 = io_x[3] ? _GEN248 : _GEN66;
wire  _GEN250 = io_x[7] ? _GEN249 : _GEN246;
wire  _GEN251 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN252 = io_x[11] ? _GEN76 : _GEN251;
wire  _GEN253 = io_x[3] ? _GEN252 : _GEN78;
wire  _GEN254 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN255 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN256 = io_x[3] ? _GEN255 : _GEN254;
wire  _GEN257 = io_x[7] ? _GEN256 : _GEN253;
wire  _GEN258 = io_x[23] ? _GEN257 : _GEN250;
wire  _GEN259 = io_x[2] ? _GEN258 : _GEN243;
wire  _GEN260 = io_x[16] ? _GEN259 : _GEN242;
wire  _GEN261 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN262 = io_x[3] ? _GEN261 : _GEN66;
wire  _GEN263 = io_x[7] ? _GEN262 : _GEN84;
wire  _GEN264 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN265 = io_x[11] ? _GEN264 : _GEN67;
wire  _GEN266 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN267 = io_x[3] ? _GEN266 : _GEN265;
wire  _GEN268 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN269 = io_x[11] ? _GEN268 : _GEN67;
wire  _GEN270 = io_x[3] ? _GEN269 : _GEN78;
wire  _GEN271 = io_x[7] ? _GEN270 : _GEN267;
wire  _GEN272 = io_x[23] ? _GEN271 : _GEN263;
wire  _GEN273 = io_x[2] ? _GEN272 : _GEN140;
wire  _GEN274 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN275 = io_x[3] ? _GEN274 : _GEN66;
wire  _GEN276 = io_x[7] ? _GEN65 : _GEN275;
wire  _GEN277 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN278 = io_x[3] ? _GEN277 : _GEN66;
wire  _GEN279 = io_x[7] ? _GEN65 : _GEN278;
wire  _GEN280 = io_x[23] ? _GEN279 : _GEN276;
wire  _GEN281 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN282 = io_x[3] ? _GEN281 : _GEN66;
wire  _GEN283 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN284 = io_x[7] ? _GEN283 : _GEN282;
wire  _GEN285 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN286 = io_x[11] ? _GEN285 : _GEN67;
wire  _GEN287 = io_x[3] ? _GEN286 : _GEN78;
wire  _GEN288 = io_x[7] ? _GEN287 : _GEN84;
wire  _GEN289 = io_x[23] ? _GEN288 : _GEN284;
wire  _GEN290 = io_x[2] ? _GEN289 : _GEN280;
wire  _GEN291 = io_x[16] ? _GEN290 : _GEN273;
wire  _GEN292 = io_x[15] ? _GEN291 : _GEN260;
wire  _GEN293 = io_x[12] ? _GEN292 : _GEN230;
wire  _GEN294 = io_x[10] ? _GEN293 : _GEN177;
wire  _GEN295 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN296 = io_x[11] ? _GEN295 : _GEN67;
wire  _GEN297 = io_x[3] ? _GEN66 : _GEN296;
wire  _GEN298 = io_x[7] ? _GEN297 : _GEN65;
wire  _GEN299 = io_x[23] ? _GEN81 : _GEN298;
wire  _GEN300 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN301 = io_x[11] ? _GEN300 : _GEN67;
wire  _GEN302 = io_x[3] ? _GEN66 : _GEN301;
wire  _GEN303 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN304 = io_x[11] ? _GEN303 : _GEN67;
wire  _GEN305 = io_x[3] ? _GEN78 : _GEN304;
wire  _GEN306 = io_x[7] ? _GEN305 : _GEN302;
wire  _GEN307 = io_x[23] ? _GEN74 : _GEN306;
wire  _GEN308 = io_x[2] ? _GEN307 : _GEN299;
wire  _GEN309 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN310 = io_x[11] ? _GEN309 : _GEN67;
wire  _GEN311 = io_x[3] ? _GEN66 : _GEN310;
wire  _GEN312 = io_x[7] ? _GEN311 : _GEN65;
wire  _GEN313 = io_x[23] ? _GEN74 : _GEN312;
wire  _GEN314 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN315 = io_x[11] ? _GEN67 : _GEN314;
wire  _GEN316 = io_x[3] ? _GEN78 : _GEN315;
wire  _GEN317 = io_x[7] ? _GEN316 : _GEN65;
wire  _GEN318 = io_x[23] ? _GEN317 : _GEN81;
wire  _GEN319 = io_x[2] ? _GEN318 : _GEN313;
wire  _GEN320 = io_x[16] ? _GEN319 : _GEN308;
wire  _GEN321 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN322 = io_x[11] ? _GEN321 : _GEN67;
wire  _GEN323 = io_x[3] ? _GEN66 : _GEN322;
wire  _GEN324 = io_x[7] ? _GEN323 : _GEN65;
wire  _GEN325 = io_x[23] ? _GEN81 : _GEN324;
wire  _GEN326 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN327 = io_x[11] ? _GEN326 : _GEN76;
wire  _GEN328 = io_x[3] ? _GEN66 : _GEN327;
wire  _GEN329 = io_x[7] ? _GEN328 : _GEN84;
wire  _GEN330 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN331 = io_x[7] ? _GEN84 : _GEN330;
wire  _GEN332 = io_x[23] ? _GEN331 : _GEN329;
wire  _GEN333 = io_x[2] ? _GEN332 : _GEN325;
wire  _GEN334 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN335 = io_x[3] ? _GEN66 : _GEN334;
wire  _GEN336 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN337 = io_x[3] ? _GEN66 : _GEN336;
wire  _GEN338 = io_x[7] ? _GEN337 : _GEN335;
wire  _GEN339 = io_x[23] ? _GEN81 : _GEN338;
wire  _GEN340 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN341 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN342 = io_x[3] ? _GEN78 : _GEN341;
wire  _GEN343 = io_x[7] ? _GEN65 : _GEN342;
wire  _GEN344 = io_x[23] ? _GEN343 : _GEN340;
wire  _GEN345 = io_x[2] ? _GEN344 : _GEN339;
wire  _GEN346 = io_x[16] ? _GEN345 : _GEN333;
wire  _GEN347 = io_x[15] ? _GEN346 : _GEN320;
wire  _GEN348 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN349 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN350 = io_x[11] ? _GEN349 : _GEN67;
wire  _GEN351 = io_x[3] ? _GEN350 : _GEN348;
wire  _GEN352 = io_x[7] ? _GEN351 : _GEN65;
wire  _GEN353 = io_x[23] ? _GEN81 : _GEN352;
wire  _GEN354 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN355 = io_x[3] ? _GEN66 : _GEN354;
wire  _GEN356 = io_x[7] ? _GEN65 : _GEN355;
wire  _GEN357 = io_x[23] ? _GEN356 : _GEN81;
wire  _GEN358 = io_x[2] ? _GEN357 : _GEN353;
wire  _GEN359 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN360 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN361 = io_x[7] ? _GEN360 : _GEN65;
wire  _GEN362 = io_x[23] ? _GEN361 : _GEN359;
wire  _GEN363 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN364 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN365 = io_x[11] ? _GEN364 : _GEN76;
wire  _GEN366 = io_x[3] ? _GEN66 : _GEN365;
wire  _GEN367 = io_x[7] ? _GEN65 : _GEN366;
wire  _GEN368 = io_x[23] ? _GEN367 : _GEN363;
wire  _GEN369 = io_x[2] ? _GEN368 : _GEN362;
wire  _GEN370 = io_x[16] ? _GEN369 : _GEN358;
wire  _GEN371 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN372 = io_x[3] ? _GEN78 : _GEN371;
wire  _GEN373 = io_x[7] ? _GEN372 : _GEN65;
wire  _GEN374 = io_x[23] ? _GEN81 : _GEN373;
wire  _GEN375 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN376 = io_x[3] ? _GEN375 : _GEN78;
wire  _GEN377 = io_x[7] ? _GEN376 : _GEN84;
wire  _GEN378 = io_x[23] ? _GEN377 : _GEN74;
wire  _GEN379 = io_x[2] ? _GEN378 : _GEN374;
wire  _GEN380 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN381 = io_x[11] ? _GEN380 : _GEN76;
wire  _GEN382 = io_x[3] ? _GEN381 : _GEN78;
wire  _GEN383 = io_x[7] ? _GEN382 : _GEN65;
wire  _GEN384 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN385 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN386 = io_x[3] ? _GEN66 : _GEN385;
wire  _GEN387 = io_x[7] ? _GEN386 : _GEN384;
wire  _GEN388 = io_x[23] ? _GEN387 : _GEN383;
wire  _GEN389 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN390 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN391 = io_x[11] ? _GEN390 : _GEN389;
wire  _GEN392 = io_x[3] ? _GEN391 : _GEN78;
wire  _GEN393 = io_x[7] ? _GEN392 : _GEN65;
wire  _GEN394 = io_x[23] ? _GEN393 : _GEN74;
wire  _GEN395 = io_x[2] ? _GEN394 : _GEN388;
wire  _GEN396 = io_x[16] ? _GEN395 : _GEN379;
wire  _GEN397 = io_x[15] ? _GEN396 : _GEN370;
wire  _GEN398 = io_x[12] ? _GEN397 : _GEN347;
wire  _GEN399 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN400 = io_x[3] ? _GEN66 : _GEN399;
wire  _GEN401 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN402 = io_x[11] ? _GEN76 : _GEN401;
wire  _GEN403 = io_x[3] ? _GEN66 : _GEN402;
wire  _GEN404 = io_x[7] ? _GEN403 : _GEN400;
wire  _GEN405 = io_x[23] ? _GEN74 : _GEN404;
wire  _GEN406 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN407 = io_x[11] ? _GEN406 : _GEN67;
wire  _GEN408 = io_x[3] ? _GEN66 : _GEN407;
wire  _GEN409 = io_x[7] ? _GEN408 : _GEN84;
wire  _GEN410 = io_x[23] ? _GEN81 : _GEN409;
wire  _GEN411 = io_x[2] ? _GEN410 : _GEN405;
wire  _GEN412 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN413 = io_x[11] ? _GEN412 : _GEN67;
wire  _GEN414 = io_x[3] ? _GEN413 : _GEN66;
wire  _GEN415 = io_x[7] ? _GEN414 : _GEN65;
wire  _GEN416 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN417 = io_x[11] ? _GEN67 : _GEN416;
wire  _GEN418 = io_x[3] ? _GEN66 : _GEN417;
wire  _GEN419 = io_x[7] ? _GEN418 : _GEN65;
wire  _GEN420 = io_x[23] ? _GEN419 : _GEN415;
wire  _GEN421 = io_x[2] ? _GEN420 : _GEN140;
wire  _GEN422 = io_x[16] ? _GEN421 : _GEN411;
wire  _GEN423 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN424 = io_x[3] ? _GEN423 : _GEN66;
wire  _GEN425 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN426 = io_x[11] ? _GEN425 : _GEN67;
wire  _GEN427 = io_x[3] ? _GEN78 : _GEN426;
wire  _GEN428 = io_x[7] ? _GEN427 : _GEN424;
wire  _GEN429 = io_x[23] ? _GEN74 : _GEN428;
wire  _GEN430 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN431 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN432 = io_x[11] ? _GEN431 : _GEN76;
wire  _GEN433 = io_x[3] ? _GEN66 : _GEN432;
wire  _GEN434 = io_x[7] ? _GEN433 : _GEN430;
wire  _GEN435 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN436 = io_x[7] ? _GEN435 : _GEN65;
wire  _GEN437 = io_x[23] ? _GEN436 : _GEN434;
wire  _GEN438 = io_x[2] ? _GEN437 : _GEN429;
wire  _GEN439 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN440 = io_x[11] ? _GEN439 : _GEN76;
wire  _GEN441 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN442 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN443 = io_x[11] ? _GEN442 : _GEN441;
wire  _GEN444 = io_x[3] ? _GEN443 : _GEN440;
wire  _GEN445 = io_x[7] ? _GEN444 : _GEN65;
wire  _GEN446 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN447 = io_x[11] ? _GEN446 : _GEN67;
wire  _GEN448 = io_x[3] ? _GEN447 : _GEN66;
wire  _GEN449 = io_x[7] ? _GEN448 : _GEN65;
wire  _GEN450 = io_x[23] ? _GEN449 : _GEN445;
wire  _GEN451 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN452 = io_x[11] ? _GEN451 : _GEN67;
wire  _GEN453 = io_x[3] ? _GEN452 : _GEN78;
wire  _GEN454 = io_x[7] ? _GEN453 : _GEN65;
wire  _GEN455 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN456 = io_x[11] ? _GEN67 : _GEN455;
wire  _GEN457 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN458 = io_x[11] ? _GEN76 : _GEN457;
wire  _GEN459 = io_x[3] ? _GEN458 : _GEN456;
wire  _GEN460 = io_x[7] ? _GEN84 : _GEN459;
wire  _GEN461 = io_x[23] ? _GEN460 : _GEN454;
wire  _GEN462 = io_x[2] ? _GEN461 : _GEN450;
wire  _GEN463 = io_x[16] ? _GEN462 : _GEN438;
wire  _GEN464 = io_x[15] ? _GEN463 : _GEN422;
wire  _GEN465 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN466 = io_x[7] ? _GEN465 : _GEN65;
wire  _GEN467 = io_x[23] ? _GEN81 : _GEN466;
wire  _GEN468 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN469 = io_x[11] ? _GEN76 : _GEN468;
wire  _GEN470 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN471 = io_x[11] ? _GEN470 : _GEN67;
wire  _GEN472 = io_x[3] ? _GEN471 : _GEN469;
wire  _GEN473 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN474 = io_x[7] ? _GEN473 : _GEN472;
wire  _GEN475 = io_x[23] ? _GEN74 : _GEN474;
wire  _GEN476 = io_x[2] ? _GEN475 : _GEN467;
wire  _GEN477 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN478 = io_x[3] ? _GEN66 : _GEN477;
wire  _GEN479 = io_x[7] ? _GEN478 : _GEN65;
wire  _GEN480 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN481 = io_x[11] ? _GEN480 : _GEN76;
wire  _GEN482 = io_x[3] ? _GEN66 : _GEN481;
wire  _GEN483 = io_x[7] ? _GEN482 : _GEN84;
wire  _GEN484 = io_x[23] ? _GEN483 : _GEN479;
wire  _GEN485 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN486 = io_x[7] ? _GEN84 : _GEN485;
wire  _GEN487 = io_x[23] ? _GEN486 : _GEN81;
wire  _GEN488 = io_x[2] ? _GEN487 : _GEN484;
wire  _GEN489 = io_x[16] ? _GEN488 : _GEN476;
wire  _GEN490 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN491 = io_x[11] ? _GEN490 : _GEN67;
wire  _GEN492 = io_x[3] ? _GEN66 : _GEN491;
wire  _GEN493 = io_x[7] ? _GEN492 : _GEN65;
wire  _GEN494 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN495 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN496 = io_x[3] ? _GEN495 : _GEN494;
wire  _GEN497 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN498 = io_x[11] ? _GEN497 : _GEN67;
wire  _GEN499 = io_x[3] ? _GEN66 : _GEN498;
wire  _GEN500 = io_x[7] ? _GEN499 : _GEN496;
wire  _GEN501 = io_x[23] ? _GEN500 : _GEN493;
wire  _GEN502 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN503 = io_x[11] ? _GEN502 : _GEN67;
wire  _GEN504 = io_x[3] ? _GEN66 : _GEN503;
wire  _GEN505 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN506 = io_x[11] ? _GEN76 : _GEN505;
wire  _GEN507 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN508 = io_x[11] ? _GEN507 : _GEN67;
wire  _GEN509 = io_x[3] ? _GEN508 : _GEN506;
wire  _GEN510 = io_x[7] ? _GEN509 : _GEN504;
wire  _GEN511 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN512 = io_x[11] ? _GEN511 : _GEN67;
wire  _GEN513 = io_x[3] ? _GEN512 : _GEN78;
wire  _GEN514 = io_x[7] ? _GEN65 : _GEN513;
wire  _GEN515 = io_x[23] ? _GEN514 : _GEN510;
wire  _GEN516 = io_x[2] ? _GEN515 : _GEN501;
wire  _GEN517 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN518 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN519 = io_x[11] ? _GEN76 : _GEN518;
wire  _GEN520 = io_x[3] ? _GEN519 : _GEN517;
wire  _GEN521 = io_x[7] ? _GEN520 : _GEN84;
wire  _GEN522 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN523 = io_x[11] ? _GEN522 : _GEN76;
wire  _GEN524 = io_x[3] ? _GEN523 : _GEN78;
wire  _GEN525 = io_x[7] ? _GEN524 : _GEN65;
wire  _GEN526 = io_x[23] ? _GEN525 : _GEN521;
wire  _GEN527 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN528 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN529 = io_x[11] ? _GEN528 : _GEN67;
wire  _GEN530 = io_x[3] ? _GEN529 : _GEN527;
wire  _GEN531 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN532 = io_x[11] ? _GEN531 : _GEN67;
wire  _GEN533 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN534 = io_x[11] ? _GEN533 : _GEN67;
wire  _GEN535 = io_x[3] ? _GEN534 : _GEN532;
wire  _GEN536 = io_x[7] ? _GEN535 : _GEN530;
wire  _GEN537 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN538 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN539 = io_x[11] ? _GEN538 : _GEN76;
wire  _GEN540 = io_x[3] ? _GEN539 : _GEN66;
wire  _GEN541 = io_x[7] ? _GEN540 : _GEN537;
wire  _GEN542 = io_x[23] ? _GEN541 : _GEN536;
wire  _GEN543 = io_x[2] ? _GEN542 : _GEN526;
wire  _GEN544 = io_x[16] ? _GEN543 : _GEN516;
wire  _GEN545 = io_x[15] ? _GEN544 : _GEN489;
wire  _GEN546 = io_x[12] ? _GEN545 : _GEN464;
wire  _GEN547 = io_x[10] ? _GEN546 : _GEN398;
wire  _GEN548 = io_x[4] ? _GEN547 : _GEN294;
wire  _GEN549 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN550 = io_x[3] ? _GEN549 : _GEN66;
wire  _GEN551 = io_x[7] ? _GEN550 : _GEN84;
wire  _GEN552 = io_x[23] ? _GEN551 : _GEN81;
wire  _GEN553 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN554 = io_x[7] ? _GEN553 : _GEN65;
wire  _GEN555 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN556 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN557 = io_x[3] ? _GEN556 : _GEN555;
wire  _GEN558 = io_x[7] ? _GEN557 : _GEN84;
wire  _GEN559 = io_x[23] ? _GEN558 : _GEN554;
wire  _GEN560 = io_x[2] ? _GEN559 : _GEN552;
wire  _GEN561 = io_x[23] ? _GEN81 : _GEN74;
wire  _GEN562 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN563 = io_x[11] ? _GEN562 : _GEN67;
wire  _GEN564 = io_x[3] ? _GEN66 : _GEN563;
wire  _GEN565 = io_x[7] ? _GEN564 : _GEN65;
wire  _GEN566 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN567 = io_x[11] ? _GEN566 : _GEN67;
wire  _GEN568 = io_x[3] ? _GEN567 : _GEN66;
wire  _GEN569 = io_x[7] ? _GEN65 : _GEN568;
wire  _GEN570 = io_x[23] ? _GEN569 : _GEN565;
wire  _GEN571 = io_x[2] ? _GEN570 : _GEN561;
wire  _GEN572 = io_x[16] ? _GEN571 : _GEN560;
wire  _GEN573 = 1'b1;
wire  _GEN574 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN575 = io_x[23] ? _GEN81 : _GEN574;
wire  _GEN576 = io_x[2] ? _GEN575 : _GEN573;
wire  _GEN577 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN578 = io_x[11] ? _GEN577 : _GEN67;
wire  _GEN579 = io_x[3] ? _GEN578 : _GEN66;
wire  _GEN580 = io_x[7] ? _GEN579 : _GEN65;
wire  _GEN581 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN582 = io_x[23] ? _GEN581 : _GEN580;
wire  _GEN583 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN584 = io_x[11] ? _GEN583 : _GEN67;
wire  _GEN585 = io_x[3] ? _GEN78 : _GEN584;
wire  _GEN586 = io_x[7] ? _GEN585 : _GEN65;
wire  _GEN587 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN588 = io_x[11] ? _GEN587 : _GEN67;
wire  _GEN589 = io_x[3] ? _GEN588 : _GEN66;
wire  _GEN590 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN591 = io_x[3] ? _GEN590 : _GEN66;
wire  _GEN592 = io_x[7] ? _GEN591 : _GEN589;
wire  _GEN593 = io_x[23] ? _GEN592 : _GEN586;
wire  _GEN594 = io_x[2] ? _GEN593 : _GEN582;
wire  _GEN595 = io_x[16] ? _GEN594 : _GEN576;
wire  _GEN596 = io_x[15] ? _GEN595 : _GEN572;
wire  _GEN597 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN598 = io_x[3] ? _GEN597 : _GEN66;
wire  _GEN599 = io_x[7] ? _GEN84 : _GEN598;
wire  _GEN600 = io_x[23] ? _GEN599 : _GEN81;
wire  _GEN601 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN602 = io_x[11] ? _GEN601 : _GEN67;
wire  _GEN603 = io_x[3] ? _GEN78 : _GEN602;
wire  _GEN604 = io_x[7] ? _GEN603 : _GEN65;
wire  _GEN605 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN606 = io_x[3] ? _GEN605 : _GEN78;
wire  _GEN607 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN608 = io_x[3] ? _GEN78 : _GEN607;
wire  _GEN609 = io_x[7] ? _GEN608 : _GEN606;
wire  _GEN610 = io_x[23] ? _GEN609 : _GEN604;
wire  _GEN611 = io_x[2] ? _GEN610 : _GEN600;
wire  _GEN612 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN613 = io_x[11] ? _GEN612 : _GEN67;
wire  _GEN614 = io_x[3] ? _GEN613 : _GEN66;
wire  _GEN615 = io_x[7] ? _GEN614 : _GEN65;
wire  _GEN616 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN617 = io_x[7] ? _GEN65 : _GEN616;
wire  _GEN618 = io_x[23] ? _GEN617 : _GEN615;
wire  _GEN619 = io_x[2] ? _GEN618 : _GEN140;
wire  _GEN620 = io_x[16] ? _GEN619 : _GEN611;
wire  _GEN621 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN622 = io_x[11] ? _GEN67 : _GEN621;
wire  _GEN623 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN624 = io_x[3] ? _GEN623 : _GEN622;
wire  _GEN625 = io_x[7] ? _GEN624 : _GEN65;
wire  _GEN626 = io_x[23] ? _GEN74 : _GEN625;
wire  _GEN627 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN628 = io_x[7] ? _GEN65 : _GEN627;
wire  _GEN629 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN630 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN631 = io_x[3] ? _GEN66 : _GEN630;
wire  _GEN632 = io_x[7] ? _GEN631 : _GEN629;
wire  _GEN633 = io_x[23] ? _GEN632 : _GEN628;
wire  _GEN634 = io_x[2] ? _GEN633 : _GEN626;
wire  _GEN635 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN636 = io_x[7] ? _GEN65 : _GEN635;
wire  _GEN637 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN638 = io_x[11] ? _GEN67 : _GEN637;
wire  _GEN639 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN640 = io_x[3] ? _GEN639 : _GEN638;
wire  _GEN641 = io_x[7] ? _GEN65 : _GEN640;
wire  _GEN642 = io_x[23] ? _GEN641 : _GEN636;
wire  _GEN643 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN644 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN645 = io_x[11] ? _GEN644 : _GEN67;
wire  _GEN646 = io_x[3] ? _GEN78 : _GEN645;
wire  _GEN647 = io_x[7] ? _GEN646 : _GEN643;
wire  _GEN648 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN649 = io_x[11] ? _GEN67 : _GEN648;
wire  _GEN650 = io_x[3] ? _GEN78 : _GEN649;
wire  _GEN651 = io_x[7] ? _GEN84 : _GEN650;
wire  _GEN652 = io_x[23] ? _GEN651 : _GEN647;
wire  _GEN653 = io_x[2] ? _GEN652 : _GEN642;
wire  _GEN654 = io_x[16] ? _GEN653 : _GEN634;
wire  _GEN655 = io_x[15] ? _GEN654 : _GEN620;
wire  _GEN656 = io_x[12] ? _GEN655 : _GEN596;
wire  _GEN657 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN658 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN659 = io_x[23] ? _GEN658 : _GEN657;
wire  _GEN660 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN661 = io_x[2] ? _GEN660 : _GEN659;
wire  _GEN662 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN663 = io_x[23] ? _GEN81 : _GEN662;
wire  _GEN664 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN665 = io_x[7] ? _GEN65 : _GEN664;
wire  _GEN666 = io_x[23] ? _GEN665 : _GEN74;
wire  _GEN667 = io_x[2] ? _GEN666 : _GEN663;
wire  _GEN668 = io_x[16] ? _GEN667 : _GEN661;
wire  _GEN669 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN670 = io_x[3] ? _GEN669 : _GEN78;
wire  _GEN671 = io_x[7] ? _GEN65 : _GEN670;
wire  _GEN672 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN673 = io_x[3] ? _GEN672 : _GEN66;
wire  _GEN674 = io_x[7] ? _GEN673 : _GEN65;
wire  _GEN675 = io_x[23] ? _GEN674 : _GEN671;
wire  _GEN676 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN677 = io_x[23] ? _GEN74 : _GEN676;
wire  _GEN678 = io_x[2] ? _GEN677 : _GEN675;
wire  _GEN679 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN680 = io_x[11] ? _GEN67 : _GEN679;
wire  _GEN681 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN682 = io_x[3] ? _GEN681 : _GEN680;
wire  _GEN683 = io_x[7] ? _GEN84 : _GEN682;
wire  _GEN684 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN685 = io_x[3] ? _GEN684 : _GEN78;
wire  _GEN686 = io_x[7] ? _GEN685 : _GEN84;
wire  _GEN687 = io_x[23] ? _GEN686 : _GEN683;
wire  _GEN688 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN689 = io_x[3] ? _GEN66 : _GEN688;
wire  _GEN690 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN691 = io_x[3] ? _GEN690 : _GEN66;
wire  _GEN692 = io_x[7] ? _GEN691 : _GEN689;
wire  _GEN693 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN694 = io_x[3] ? _GEN66 : _GEN693;
wire  _GEN695 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN696 = io_x[3] ? _GEN695 : _GEN66;
wire  _GEN697 = io_x[7] ? _GEN696 : _GEN694;
wire  _GEN698 = io_x[23] ? _GEN697 : _GEN692;
wire  _GEN699 = io_x[2] ? _GEN698 : _GEN687;
wire  _GEN700 = io_x[16] ? _GEN699 : _GEN678;
wire  _GEN701 = io_x[15] ? _GEN700 : _GEN668;
wire  _GEN702 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN703 = io_x[3] ? _GEN702 : _GEN66;
wire  _GEN704 = io_x[7] ? _GEN703 : _GEN84;
wire  _GEN705 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN706 = io_x[23] ? _GEN705 : _GEN704;
wire  _GEN707 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN708 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN709 = io_x[11] ? _GEN708 : _GEN67;
wire  _GEN710 = io_x[3] ? _GEN709 : _GEN707;
wire  _GEN711 = io_x[7] ? _GEN710 : _GEN84;
wire  _GEN712 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN713 = io_x[3] ? _GEN78 : _GEN712;
wire  _GEN714 = io_x[7] ? _GEN65 : _GEN713;
wire  _GEN715 = io_x[23] ? _GEN714 : _GEN711;
wire  _GEN716 = io_x[2] ? _GEN715 : _GEN706;
wire  _GEN717 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN718 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN719 = io_x[11] ? _GEN718 : _GEN67;
wire  _GEN720 = io_x[3] ? _GEN66 : _GEN719;
wire  _GEN721 = io_x[7] ? _GEN720 : _GEN65;
wire  _GEN722 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN723 = io_x[3] ? _GEN66 : _GEN722;
wire  _GEN724 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN725 = io_x[3] ? _GEN724 : _GEN66;
wire  _GEN726 = io_x[7] ? _GEN725 : _GEN723;
wire  _GEN727 = io_x[23] ? _GEN726 : _GEN721;
wire  _GEN728 = io_x[2] ? _GEN727 : _GEN717;
wire  _GEN729 = io_x[16] ? _GEN728 : _GEN716;
wire  _GEN730 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN731 = io_x[3] ? _GEN730 : _GEN78;
wire  _GEN732 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN733 = io_x[11] ? _GEN732 : _GEN76;
wire  _GEN734 = io_x[3] ? _GEN733 : _GEN66;
wire  _GEN735 = io_x[7] ? _GEN734 : _GEN731;
wire  _GEN736 = io_x[23] ? _GEN81 : _GEN735;
wire  _GEN737 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN738 = io_x[11] ? _GEN76 : _GEN737;
wire  _GEN739 = io_x[3] ? _GEN66 : _GEN738;
wire  _GEN740 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN741 = io_x[11] ? _GEN740 : _GEN67;
wire  _GEN742 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN743 = io_x[11] ? _GEN742 : _GEN76;
wire  _GEN744 = io_x[3] ? _GEN743 : _GEN741;
wire  _GEN745 = io_x[7] ? _GEN744 : _GEN739;
wire  _GEN746 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN747 = io_x[11] ? _GEN746 : _GEN67;
wire  _GEN748 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN749 = io_x[11] ? _GEN748 : _GEN76;
wire  _GEN750 = io_x[3] ? _GEN749 : _GEN747;
wire  _GEN751 = io_x[7] ? _GEN750 : _GEN84;
wire  _GEN752 = io_x[23] ? _GEN751 : _GEN745;
wire  _GEN753 = io_x[2] ? _GEN752 : _GEN736;
wire  _GEN754 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN755 = io_x[11] ? _GEN67 : _GEN754;
wire  _GEN756 = io_x[3] ? _GEN755 : _GEN66;
wire  _GEN757 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN758 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN759 = io_x[3] ? _GEN758 : _GEN757;
wire  _GEN760 = io_x[7] ? _GEN759 : _GEN756;
wire  _GEN761 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN762 = io_x[7] ? _GEN761 : _GEN84;
wire  _GEN763 = io_x[23] ? _GEN762 : _GEN760;
wire  _GEN764 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN765 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN766 = io_x[11] ? _GEN765 : _GEN67;
wire  _GEN767 = io_x[3] ? _GEN766 : _GEN764;
wire  _GEN768 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN769 = io_x[11] ? _GEN768 : _GEN67;
wire  _GEN770 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN771 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN772 = io_x[11] ? _GEN771 : _GEN770;
wire  _GEN773 = io_x[3] ? _GEN772 : _GEN769;
wire  _GEN774 = io_x[7] ? _GEN773 : _GEN767;
wire  _GEN775 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN776 = io_x[11] ? _GEN775 : _GEN67;
wire  _GEN777 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN778 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN779 = io_x[11] ? _GEN778 : _GEN777;
wire  _GEN780 = io_x[3] ? _GEN779 : _GEN776;
wire  _GEN781 = io_x[7] ? _GEN780 : _GEN65;
wire  _GEN782 = io_x[23] ? _GEN781 : _GEN774;
wire  _GEN783 = io_x[2] ? _GEN782 : _GEN763;
wire  _GEN784 = io_x[16] ? _GEN783 : _GEN753;
wire  _GEN785 = io_x[15] ? _GEN784 : _GEN729;
wire  _GEN786 = io_x[12] ? _GEN785 : _GEN701;
wire  _GEN787 = io_x[10] ? _GEN786 : _GEN656;
wire  _GEN788 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN789 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN790 = io_x[7] ? _GEN65 : _GEN789;
wire  _GEN791 = io_x[23] ? _GEN790 : _GEN788;
wire  _GEN792 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN793 = io_x[11] ? _GEN792 : _GEN67;
wire  _GEN794 = io_x[3] ? _GEN66 : _GEN793;
wire  _GEN795 = io_x[7] ? _GEN65 : _GEN794;
wire  _GEN796 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN797 = io_x[7] ? _GEN796 : _GEN65;
wire  _GEN798 = io_x[23] ? _GEN797 : _GEN795;
wire  _GEN799 = io_x[2] ? _GEN798 : _GEN791;
wire  _GEN800 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN801 = io_x[11] ? _GEN800 : _GEN67;
wire  _GEN802 = io_x[3] ? _GEN801 : _GEN66;
wire  _GEN803 = io_x[7] ? _GEN802 : _GEN84;
wire  _GEN804 = io_x[23] ? _GEN81 : _GEN803;
wire  _GEN805 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN806 = io_x[3] ? _GEN66 : _GEN805;
wire  _GEN807 = io_x[7] ? _GEN65 : _GEN806;
wire  _GEN808 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN809 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN810 = io_x[11] ? _GEN809 : _GEN67;
wire  _GEN811 = io_x[3] ? _GEN810 : _GEN66;
wire  _GEN812 = io_x[7] ? _GEN811 : _GEN808;
wire  _GEN813 = io_x[23] ? _GEN812 : _GEN807;
wire  _GEN814 = io_x[2] ? _GEN813 : _GEN804;
wire  _GEN815 = io_x[16] ? _GEN814 : _GEN799;
wire  _GEN816 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN817 = io_x[11] ? _GEN816 : _GEN67;
wire  _GEN818 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN819 = io_x[11] ? _GEN818 : _GEN67;
wire  _GEN820 = io_x[3] ? _GEN819 : _GEN817;
wire  _GEN821 = io_x[7] ? _GEN820 : _GEN65;
wire  _GEN822 = io_x[23] ? _GEN74 : _GEN821;
wire  _GEN823 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN824 = io_x[11] ? _GEN823 : _GEN67;
wire  _GEN825 = io_x[3] ? _GEN66 : _GEN824;
wire  _GEN826 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN827 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN828 = io_x[11] ? _GEN827 : _GEN67;
wire  _GEN829 = io_x[3] ? _GEN828 : _GEN826;
wire  _GEN830 = io_x[7] ? _GEN829 : _GEN825;
wire  _GEN831 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN832 = io_x[7] ? _GEN831 : _GEN65;
wire  _GEN833 = io_x[23] ? _GEN832 : _GEN830;
wire  _GEN834 = io_x[2] ? _GEN833 : _GEN822;
wire  _GEN835 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN836 = io_x[11] ? _GEN835 : _GEN67;
wire  _GEN837 = io_x[3] ? _GEN66 : _GEN836;
wire  _GEN838 = io_x[7] ? _GEN837 : _GEN65;
wire  _GEN839 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN840 = io_x[11] ? _GEN839 : _GEN67;
wire  _GEN841 = io_x[3] ? _GEN840 : _GEN78;
wire  _GEN842 = io_x[7] ? _GEN841 : _GEN84;
wire  _GEN843 = io_x[23] ? _GEN842 : _GEN838;
wire  _GEN844 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN845 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN846 = io_x[11] ? _GEN845 : _GEN67;
wire  _GEN847 = io_x[3] ? _GEN846 : _GEN66;
wire  _GEN848 = io_x[7] ? _GEN847 : _GEN844;
wire  _GEN849 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN850 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN851 = io_x[11] ? _GEN850 : _GEN67;
wire  _GEN852 = io_x[3] ? _GEN851 : _GEN849;
wire  _GEN853 = io_x[7] ? _GEN852 : _GEN65;
wire  _GEN854 = io_x[23] ? _GEN853 : _GEN848;
wire  _GEN855 = io_x[2] ? _GEN854 : _GEN843;
wire  _GEN856 = io_x[16] ? _GEN855 : _GEN834;
wire  _GEN857 = io_x[15] ? _GEN856 : _GEN815;
wire  _GEN858 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN859 = io_x[11] ? _GEN858 : _GEN67;
wire  _GEN860 = io_x[3] ? _GEN859 : _GEN78;
wire  _GEN861 = io_x[7] ? _GEN860 : _GEN65;
wire  _GEN862 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN863 = io_x[3] ? _GEN862 : _GEN66;
wire  _GEN864 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN865 = io_x[7] ? _GEN864 : _GEN863;
wire  _GEN866 = io_x[23] ? _GEN865 : _GEN861;
wire  _GEN867 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN868 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN869 = io_x[11] ? _GEN868 : _GEN67;
wire  _GEN870 = io_x[3] ? _GEN869 : _GEN66;
wire  _GEN871 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN872 = io_x[11] ? _GEN67 : _GEN871;
wire  _GEN873 = io_x[3] ? _GEN872 : _GEN78;
wire  _GEN874 = io_x[7] ? _GEN873 : _GEN870;
wire  _GEN875 = io_x[23] ? _GEN874 : _GEN867;
wire  _GEN876 = io_x[2] ? _GEN875 : _GEN866;
wire  _GEN877 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN878 = io_x[23] ? _GEN81 : _GEN877;
wire  _GEN879 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN880 = io_x[11] ? _GEN879 : _GEN67;
wire  _GEN881 = io_x[3] ? _GEN880 : _GEN66;
wire  _GEN882 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN883 = io_x[11] ? _GEN882 : _GEN67;
wire  _GEN884 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN885 = io_x[11] ? _GEN884 : _GEN67;
wire  _GEN886 = io_x[3] ? _GEN885 : _GEN883;
wire  _GEN887 = io_x[7] ? _GEN886 : _GEN881;
wire  _GEN888 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN889 = io_x[3] ? _GEN888 : _GEN66;
wire  _GEN890 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN891 = io_x[11] ? _GEN890 : _GEN67;
wire  _GEN892 = io_x[3] ? _GEN66 : _GEN891;
wire  _GEN893 = io_x[7] ? _GEN892 : _GEN889;
wire  _GEN894 = io_x[23] ? _GEN893 : _GEN887;
wire  _GEN895 = io_x[2] ? _GEN894 : _GEN878;
wire  _GEN896 = io_x[16] ? _GEN895 : _GEN876;
wire  _GEN897 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN898 = io_x[3] ? _GEN897 : _GEN66;
wire  _GEN899 = io_x[7] ? _GEN84 : _GEN898;
wire  _GEN900 = io_x[23] ? _GEN899 : _GEN81;
wire  _GEN901 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN902 = io_x[11] ? _GEN76 : _GEN901;
wire  _GEN903 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN904 = io_x[11] ? _GEN76 : _GEN903;
wire  _GEN905 = io_x[3] ? _GEN904 : _GEN902;
wire  _GEN906 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN907 = io_x[11] ? _GEN906 : _GEN67;
wire  _GEN908 = io_x[3] ? _GEN907 : _GEN66;
wire  _GEN909 = io_x[7] ? _GEN908 : _GEN905;
wire  _GEN910 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN911 = io_x[11] ? _GEN910 : _GEN67;
wire  _GEN912 = io_x[3] ? _GEN911 : _GEN78;
wire  _GEN913 = io_x[7] ? _GEN65 : _GEN912;
wire  _GEN914 = io_x[23] ? _GEN913 : _GEN909;
wire  _GEN915 = io_x[2] ? _GEN914 : _GEN900;
wire  _GEN916 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN917 = io_x[11] ? _GEN67 : _GEN916;
wire  _GEN918 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN919 = io_x[11] ? _GEN67 : _GEN918;
wire  _GEN920 = io_x[3] ? _GEN919 : _GEN917;
wire  _GEN921 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN922 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN923 = io_x[11] ? _GEN922 : _GEN921;
wire  _GEN924 = io_x[3] ? _GEN923 : _GEN66;
wire  _GEN925 = io_x[7] ? _GEN924 : _GEN920;
wire  _GEN926 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN927 = io_x[3] ? _GEN926 : _GEN66;
wire  _GEN928 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN929 = io_x[3] ? _GEN928 : _GEN78;
wire  _GEN930 = io_x[7] ? _GEN929 : _GEN927;
wire  _GEN931 = io_x[23] ? _GEN930 : _GEN925;
wire  _GEN932 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN933 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN934 = io_x[3] ? _GEN933 : _GEN932;
wire  _GEN935 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN936 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN937 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN938 = io_x[11] ? _GEN937 : _GEN936;
wire  _GEN939 = io_x[3] ? _GEN938 : _GEN935;
wire  _GEN940 = io_x[7] ? _GEN939 : _GEN934;
wire  _GEN941 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN942 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN943 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN944 = io_x[11] ? _GEN943 : _GEN942;
wire  _GEN945 = io_x[3] ? _GEN944 : _GEN941;
wire  _GEN946 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN947 = io_x[11] ? _GEN946 : _GEN67;
wire  _GEN948 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN949 = io_x[11] ? _GEN948 : _GEN67;
wire  _GEN950 = io_x[3] ? _GEN949 : _GEN947;
wire  _GEN951 = io_x[7] ? _GEN950 : _GEN945;
wire  _GEN952 = io_x[23] ? _GEN951 : _GEN940;
wire  _GEN953 = io_x[2] ? _GEN952 : _GEN931;
wire  _GEN954 = io_x[16] ? _GEN953 : _GEN915;
wire  _GEN955 = io_x[15] ? _GEN954 : _GEN896;
wire  _GEN956 = io_x[12] ? _GEN955 : _GEN857;
wire  _GEN957 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN958 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN959 = io_x[11] ? _GEN76 : _GEN958;
wire  _GEN960 = io_x[3] ? _GEN66 : _GEN959;
wire  _GEN961 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN962 = io_x[11] ? _GEN76 : _GEN961;
wire  _GEN963 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN964 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN965 = io_x[11] ? _GEN964 : _GEN963;
wire  _GEN966 = io_x[3] ? _GEN965 : _GEN962;
wire  _GEN967 = io_x[7] ? _GEN966 : _GEN960;
wire  _GEN968 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN969 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN970 = io_x[11] ? _GEN969 : _GEN67;
wire  _GEN971 = io_x[3] ? _GEN970 : _GEN968;
wire  _GEN972 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN973 = io_x[3] ? _GEN66 : _GEN972;
wire  _GEN974 = io_x[7] ? _GEN973 : _GEN971;
wire  _GEN975 = io_x[23] ? _GEN974 : _GEN967;
wire  _GEN976 = io_x[2] ? _GEN975 : _GEN957;
wire  _GEN977 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN978 = io_x[3] ? _GEN977 : _GEN78;
wire  _GEN979 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN980 = io_x[11] ? _GEN979 : _GEN67;
wire  _GEN981 = io_x[3] ? _GEN980 : _GEN66;
wire  _GEN982 = io_x[7] ? _GEN981 : _GEN978;
wire  _GEN983 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN984 = io_x[11] ? _GEN76 : _GEN983;
wire  _GEN985 = io_x[3] ? _GEN984 : _GEN66;
wire  _GEN986 = io_x[7] ? _GEN65 : _GEN985;
wire  _GEN987 = io_x[23] ? _GEN986 : _GEN982;
wire  _GEN988 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN989 = io_x[11] ? _GEN988 : _GEN67;
wire  _GEN990 = io_x[3] ? _GEN78 : _GEN989;
wire  _GEN991 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN992 = io_x[11] ? _GEN76 : _GEN991;
wire  _GEN993 = io_x[3] ? _GEN66 : _GEN992;
wire  _GEN994 = io_x[7] ? _GEN993 : _GEN990;
wire  _GEN995 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN996 = io_x[3] ? _GEN995 : _GEN66;
wire  _GEN997 = io_x[7] ? _GEN996 : _GEN84;
wire  _GEN998 = io_x[23] ? _GEN997 : _GEN994;
wire  _GEN999 = io_x[2] ? _GEN998 : _GEN987;
wire  _GEN1000 = io_x[16] ? _GEN999 : _GEN976;
wire  _GEN1001 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1002 = io_x[11] ? _GEN76 : _GEN1001;
wire  _GEN1003 = io_x[3] ? _GEN1002 : _GEN66;
wire  _GEN1004 = io_x[7] ? _GEN84 : _GEN1003;
wire  _GEN1005 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1006 = io_x[7] ? _GEN65 : _GEN1005;
wire  _GEN1007 = io_x[23] ? _GEN1006 : _GEN1004;
wire  _GEN1008 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1009 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1010 = io_x[11] ? _GEN1009 : _GEN1008;
wire  _GEN1011 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1012 = io_x[11] ? _GEN1011 : _GEN67;
wire  _GEN1013 = io_x[3] ? _GEN1012 : _GEN1010;
wire  _GEN1014 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1015 = io_x[7] ? _GEN1014 : _GEN1013;
wire  _GEN1016 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1017 = io_x[11] ? _GEN1016 : _GEN67;
wire  _GEN1018 = io_x[3] ? _GEN1017 : _GEN66;
wire  _GEN1019 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1020 = io_x[11] ? _GEN1019 : _GEN76;
wire  _GEN1021 = io_x[3] ? _GEN1020 : _GEN66;
wire  _GEN1022 = io_x[7] ? _GEN1021 : _GEN1018;
wire  _GEN1023 = io_x[23] ? _GEN1022 : _GEN1015;
wire  _GEN1024 = io_x[2] ? _GEN1023 : _GEN1007;
wire  _GEN1025 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1026 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1027 = io_x[3] ? _GEN1026 : _GEN1025;
wire  _GEN1028 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1029 = io_x[3] ? _GEN1028 : _GEN78;
wire  _GEN1030 = io_x[7] ? _GEN1029 : _GEN1027;
wire  _GEN1031 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1032 = io_x[11] ? _GEN67 : _GEN1031;
wire  _GEN1033 = io_x[3] ? _GEN1032 : _GEN66;
wire  _GEN1034 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1035 = io_x[11] ? _GEN1034 : _GEN67;
wire  _GEN1036 = io_x[3] ? _GEN1035 : _GEN66;
wire  _GEN1037 = io_x[7] ? _GEN1036 : _GEN1033;
wire  _GEN1038 = io_x[23] ? _GEN1037 : _GEN1030;
wire  _GEN1039 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1040 = io_x[11] ? _GEN1039 : _GEN67;
wire  _GEN1041 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1042 = io_x[11] ? _GEN1041 : _GEN67;
wire  _GEN1043 = io_x[3] ? _GEN1042 : _GEN1040;
wire  _GEN1044 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1045 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1046 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1047 = io_x[11] ? _GEN1046 : _GEN1045;
wire  _GEN1048 = io_x[3] ? _GEN1047 : _GEN1044;
wire  _GEN1049 = io_x[7] ? _GEN1048 : _GEN1043;
wire  _GEN1050 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1051 = io_x[11] ? _GEN1050 : _GEN67;
wire  _GEN1052 = io_x[3] ? _GEN1051 : _GEN66;
wire  _GEN1053 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1054 = io_x[11] ? _GEN1053 : _GEN67;
wire  _GEN1055 = io_x[3] ? _GEN1054 : _GEN66;
wire  _GEN1056 = io_x[7] ? _GEN1055 : _GEN1052;
wire  _GEN1057 = io_x[23] ? _GEN1056 : _GEN1049;
wire  _GEN1058 = io_x[2] ? _GEN1057 : _GEN1038;
wire  _GEN1059 = io_x[16] ? _GEN1058 : _GEN1024;
wire  _GEN1060 = io_x[15] ? _GEN1059 : _GEN1000;
wire  _GEN1061 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1062 = io_x[11] ? _GEN1061 : _GEN67;
wire  _GEN1063 = io_x[3] ? _GEN1062 : _GEN78;
wire  _GEN1064 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1065 = io_x[3] ? _GEN1064 : _GEN66;
wire  _GEN1066 = io_x[7] ? _GEN1065 : _GEN1063;
wire  _GEN1067 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1068 = io_x[3] ? _GEN66 : _GEN1067;
wire  _GEN1069 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1070 = io_x[7] ? _GEN1069 : _GEN1068;
wire  _GEN1071 = io_x[23] ? _GEN1070 : _GEN1066;
wire  _GEN1072 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1073 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1074 = io_x[11] ? _GEN1073 : _GEN1072;
wire  _GEN1075 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1076 = io_x[3] ? _GEN1075 : _GEN1074;
wire  _GEN1077 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1078 = io_x[11] ? _GEN1077 : _GEN67;
wire  _GEN1079 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1080 = io_x[11] ? _GEN1079 : _GEN76;
wire  _GEN1081 = io_x[3] ? _GEN1080 : _GEN1078;
wire  _GEN1082 = io_x[7] ? _GEN1081 : _GEN1076;
wire  _GEN1083 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1084 = io_x[11] ? _GEN1083 : _GEN67;
wire  _GEN1085 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1086 = io_x[3] ? _GEN1085 : _GEN1084;
wire  _GEN1087 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1088 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1089 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1090 = io_x[11] ? _GEN1089 : _GEN1088;
wire  _GEN1091 = io_x[3] ? _GEN1090 : _GEN1087;
wire  _GEN1092 = io_x[7] ? _GEN1091 : _GEN1086;
wire  _GEN1093 = io_x[23] ? _GEN1092 : _GEN1082;
wire  _GEN1094 = io_x[2] ? _GEN1093 : _GEN1071;
wire  _GEN1095 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1096 = io_x[23] ? _GEN81 : _GEN1095;
wire  _GEN1097 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1098 = io_x[11] ? _GEN67 : _GEN1097;
wire  _GEN1099 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1100 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1101 = io_x[11] ? _GEN1100 : _GEN1099;
wire  _GEN1102 = io_x[3] ? _GEN1101 : _GEN1098;
wire  _GEN1103 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1104 = io_x[11] ? _GEN1103 : _GEN67;
wire  _GEN1105 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1106 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1107 = io_x[11] ? _GEN1106 : _GEN1105;
wire  _GEN1108 = io_x[3] ? _GEN1107 : _GEN1104;
wire  _GEN1109 = io_x[7] ? _GEN1108 : _GEN1102;
wire  _GEN1110 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1111 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1112 = io_x[11] ? _GEN1111 : _GEN1110;
wire  _GEN1113 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1114 = io_x[3] ? _GEN1113 : _GEN1112;
wire  _GEN1115 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1116 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1117 = io_x[11] ? _GEN1116 : _GEN1115;
wire  _GEN1118 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1119 = io_x[11] ? _GEN1118 : _GEN76;
wire  _GEN1120 = io_x[3] ? _GEN1119 : _GEN1117;
wire  _GEN1121 = io_x[7] ? _GEN1120 : _GEN1114;
wire  _GEN1122 = io_x[23] ? _GEN1121 : _GEN1109;
wire  _GEN1123 = io_x[2] ? _GEN1122 : _GEN1096;
wire  _GEN1124 = io_x[16] ? _GEN1123 : _GEN1094;
wire  _GEN1125 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1126 = io_x[3] ? _GEN1125 : _GEN66;
wire  _GEN1127 = io_x[7] ? _GEN1126 : _GEN65;
wire  _GEN1128 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1129 = io_x[3] ? _GEN1128 : _GEN78;
wire  _GEN1130 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1131 = io_x[11] ? _GEN1130 : _GEN76;
wire  _GEN1132 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1133 = io_x[11] ? _GEN1132 : _GEN67;
wire  _GEN1134 = io_x[3] ? _GEN1133 : _GEN1131;
wire  _GEN1135 = io_x[7] ? _GEN1134 : _GEN1129;
wire  _GEN1136 = io_x[23] ? _GEN1135 : _GEN1127;
wire  _GEN1137 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1138 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1139 = io_x[11] ? _GEN1138 : _GEN1137;
wire  _GEN1140 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1141 = io_x[11] ? _GEN1140 : _GEN76;
wire  _GEN1142 = io_x[3] ? _GEN1141 : _GEN1139;
wire  _GEN1143 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1144 = io_x[11] ? _GEN67 : _GEN1143;
wire  _GEN1145 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1146 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1147 = io_x[11] ? _GEN1146 : _GEN1145;
wire  _GEN1148 = io_x[3] ? _GEN1147 : _GEN1144;
wire  _GEN1149 = io_x[7] ? _GEN1148 : _GEN1142;
wire  _GEN1150 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1151 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1152 = io_x[11] ? _GEN1151 : _GEN67;
wire  _GEN1153 = io_x[3] ? _GEN1152 : _GEN1150;
wire  _GEN1154 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1155 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1156 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1157 = io_x[11] ? _GEN1156 : _GEN1155;
wire  _GEN1158 = io_x[3] ? _GEN1157 : _GEN1154;
wire  _GEN1159 = io_x[7] ? _GEN1158 : _GEN1153;
wire  _GEN1160 = io_x[23] ? _GEN1159 : _GEN1149;
wire  _GEN1161 = io_x[2] ? _GEN1160 : _GEN1136;
wire  _GEN1162 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1163 = io_x[11] ? _GEN1162 : _GEN67;
wire  _GEN1164 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1165 = io_x[11] ? _GEN1164 : _GEN67;
wire  _GEN1166 = io_x[3] ? _GEN1165 : _GEN1163;
wire  _GEN1167 = io_x[7] ? _GEN1166 : _GEN65;
wire  _GEN1168 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1169 = io_x[11] ? _GEN1168 : _GEN76;
wire  _GEN1170 = io_x[3] ? _GEN1169 : _GEN66;
wire  _GEN1171 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1172 = io_x[11] ? _GEN1171 : _GEN67;
wire  _GEN1173 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1174 = io_x[11] ? _GEN1173 : _GEN67;
wire  _GEN1175 = io_x[3] ? _GEN1174 : _GEN1172;
wire  _GEN1176 = io_x[7] ? _GEN1175 : _GEN1170;
wire  _GEN1177 = io_x[23] ? _GEN1176 : _GEN1167;
wire  _GEN1178 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1179 = io_x[11] ? _GEN76 : _GEN1178;
wire  _GEN1180 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1181 = io_x[11] ? _GEN1180 : _GEN76;
wire  _GEN1182 = io_x[3] ? _GEN1181 : _GEN1179;
wire  _GEN1183 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1184 = io_x[11] ? _GEN1183 : _GEN76;
wire  _GEN1185 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1186 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1187 = io_x[11] ? _GEN1186 : _GEN1185;
wire  _GEN1188 = io_x[3] ? _GEN1187 : _GEN1184;
wire  _GEN1189 = io_x[7] ? _GEN1188 : _GEN1182;
wire  _GEN1190 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1191 = io_x[11] ? _GEN1190 : _GEN76;
wire  _GEN1192 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1193 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1194 = io_x[11] ? _GEN1193 : _GEN1192;
wire  _GEN1195 = io_x[3] ? _GEN1194 : _GEN1191;
wire  _GEN1196 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1197 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1198 = io_x[11] ? _GEN1197 : _GEN1196;
wire  _GEN1199 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1200 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1201 = io_x[11] ? _GEN1200 : _GEN1199;
wire  _GEN1202 = io_x[3] ? _GEN1201 : _GEN1198;
wire  _GEN1203 = io_x[7] ? _GEN1202 : _GEN1195;
wire  _GEN1204 = io_x[23] ? _GEN1203 : _GEN1189;
wire  _GEN1205 = io_x[2] ? _GEN1204 : _GEN1177;
wire  _GEN1206 = io_x[16] ? _GEN1205 : _GEN1161;
wire  _GEN1207 = io_x[15] ? _GEN1206 : _GEN1124;
wire  _GEN1208 = io_x[12] ? _GEN1207 : _GEN1060;
wire  _GEN1209 = io_x[10] ? _GEN1208 : _GEN956;
wire  _GEN1210 = io_x[4] ? _GEN1209 : _GEN787;
wire  _GEN1211 = io_x[8] ? _GEN1210 : _GEN548;
wire  _GEN1212 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN1213 = io_x[2] ? _GEN573 : _GEN1212;
wire  _GEN1214 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1215 = io_x[11] ? _GEN1214 : _GEN67;
wire  _GEN1216 = io_x[3] ? _GEN1215 : _GEN66;
wire  _GEN1217 = io_x[7] ? _GEN1216 : _GEN65;
wire  _GEN1218 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1219 = io_x[11] ? _GEN1218 : _GEN67;
wire  _GEN1220 = io_x[3] ? _GEN1219 : _GEN66;
wire  _GEN1221 = io_x[7] ? _GEN1220 : _GEN65;
wire  _GEN1222 = io_x[23] ? _GEN1221 : _GEN1217;
wire  _GEN1223 = io_x[2] ? _GEN573 : _GEN1222;
wire  _GEN1224 = io_x[16] ? _GEN1223 : _GEN1213;
wire  _GEN1225 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1226 = io_x[3] ? _GEN1225 : _GEN66;
wire  _GEN1227 = io_x[7] ? _GEN65 : _GEN1226;
wire  _GEN1228 = io_x[23] ? _GEN81 : _GEN1227;
wire  _GEN1229 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1230 = io_x[7] ? _GEN1229 : _GEN65;
wire  _GEN1231 = io_x[23] ? _GEN1230 : _GEN74;
wire  _GEN1232 = io_x[2] ? _GEN1231 : _GEN1228;
wire  _GEN1233 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1234 = io_x[23] ? _GEN1233 : _GEN81;
wire  _GEN1235 = io_x[2] ? _GEN573 : _GEN1234;
wire  _GEN1236 = io_x[16] ? _GEN1235 : _GEN1232;
wire  _GEN1237 = io_x[15] ? _GEN1236 : _GEN1224;
wire  _GEN1238 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN1239 = io_x[2] ? _GEN1238 : _GEN140;
wire  _GEN1240 = 1'b1;
wire  _GEN1241 = io_x[16] ? _GEN1240 : _GEN1239;
wire  _GEN1242 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1243 = io_x[3] ? _GEN1242 : _GEN66;
wire  _GEN1244 = io_x[7] ? _GEN84 : _GEN1243;
wire  _GEN1245 = io_x[23] ? _GEN81 : _GEN1244;
wire  _GEN1246 = io_x[2] ? _GEN140 : _GEN1245;
wire  _GEN1247 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1248 = io_x[7] ? _GEN65 : _GEN1247;
wire  _GEN1249 = io_x[23] ? _GEN1248 : _GEN81;
wire  _GEN1250 = io_x[2] ? _GEN1249 : _GEN573;
wire  _GEN1251 = io_x[16] ? _GEN1250 : _GEN1246;
wire  _GEN1252 = io_x[15] ? _GEN1251 : _GEN1241;
wire  _GEN1253 = io_x[12] ? _GEN1252 : _GEN1237;
wire  _GEN1254 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1255 = io_x[3] ? _GEN1254 : _GEN66;
wire  _GEN1256 = io_x[7] ? _GEN1255 : _GEN84;
wire  _GEN1257 = io_x[23] ? _GEN81 : _GEN1256;
wire  _GEN1258 = io_x[2] ? _GEN1257 : _GEN573;
wire  _GEN1259 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN1260 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1261 = io_x[11] ? _GEN1260 : _GEN76;
wire  _GEN1262 = io_x[3] ? _GEN1261 : _GEN66;
wire  _GEN1263 = io_x[7] ? _GEN1262 : _GEN65;
wire  _GEN1264 = io_x[23] ? _GEN81 : _GEN1263;
wire  _GEN1265 = io_x[2] ? _GEN1264 : _GEN1259;
wire  _GEN1266 = io_x[16] ? _GEN1265 : _GEN1258;
wire  _GEN1267 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1268 = io_x[23] ? _GEN1267 : _GEN81;
wire  _GEN1269 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1270 = io_x[3] ? _GEN66 : _GEN1269;
wire  _GEN1271 = io_x[7] ? _GEN84 : _GEN1270;
wire  _GEN1272 = io_x[23] ? _GEN81 : _GEN1271;
wire  _GEN1273 = io_x[2] ? _GEN1272 : _GEN1268;
wire  _GEN1274 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1275 = io_x[11] ? _GEN1274 : _GEN67;
wire  _GEN1276 = io_x[3] ? _GEN1275 : _GEN66;
wire  _GEN1277 = io_x[7] ? _GEN1276 : _GEN65;
wire  _GEN1278 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1279 = io_x[3] ? _GEN78 : _GEN1278;
wire  _GEN1280 = io_x[7] ? _GEN1279 : _GEN65;
wire  _GEN1281 = io_x[23] ? _GEN1280 : _GEN1277;
wire  _GEN1282 = io_x[2] ? _GEN1281 : _GEN573;
wire  _GEN1283 = io_x[16] ? _GEN1282 : _GEN1273;
wire  _GEN1284 = io_x[15] ? _GEN1283 : _GEN1266;
wire  _GEN1285 = io_x[23] ? _GEN81 : _GEN74;
wire  _GEN1286 = io_x[2] ? _GEN1285 : _GEN140;
wire  _GEN1287 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1288 = io_x[11] ? _GEN67 : _GEN1287;
wire  _GEN1289 = io_x[3] ? _GEN1288 : _GEN66;
wire  _GEN1290 = io_x[7] ? _GEN1289 : _GEN65;
wire  _GEN1291 = io_x[23] ? _GEN1290 : _GEN81;
wire  _GEN1292 = io_x[2] ? _GEN1291 : _GEN573;
wire  _GEN1293 = io_x[16] ? _GEN1292 : _GEN1286;
wire  _GEN1294 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1295 = io_x[3] ? _GEN1294 : _GEN66;
wire  _GEN1296 = io_x[7] ? _GEN1295 : _GEN65;
wire  _GEN1297 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1298 = io_x[3] ? _GEN78 : _GEN1297;
wire  _GEN1299 = io_x[7] ? _GEN1298 : _GEN65;
wire  _GEN1300 = io_x[23] ? _GEN1299 : _GEN1296;
wire  _GEN1301 = io_x[2] ? _GEN1300 : _GEN573;
wire  _GEN1302 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1303 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1304 = io_x[11] ? _GEN67 : _GEN1303;
wire  _GEN1305 = io_x[3] ? _GEN1304 : _GEN66;
wire  _GEN1306 = io_x[7] ? _GEN1305 : _GEN1302;
wire  _GEN1307 = io_x[23] ? _GEN1306 : _GEN81;
wire  _GEN1308 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1309 = io_x[3] ? _GEN1308 : _GEN66;
wire  _GEN1310 = io_x[7] ? _GEN1309 : _GEN65;
wire  _GEN1311 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1312 = io_x[11] ? _GEN1311 : _GEN76;
wire  _GEN1313 = io_x[3] ? _GEN1312 : _GEN66;
wire  _GEN1314 = io_x[7] ? _GEN1313 : _GEN65;
wire  _GEN1315 = io_x[23] ? _GEN1314 : _GEN1310;
wire  _GEN1316 = io_x[2] ? _GEN1315 : _GEN1307;
wire  _GEN1317 = io_x[16] ? _GEN1316 : _GEN1301;
wire  _GEN1318 = io_x[15] ? _GEN1317 : _GEN1293;
wire  _GEN1319 = io_x[12] ? _GEN1318 : _GEN1284;
wire  _GEN1320 = io_x[10] ? _GEN1319 : _GEN1253;
wire  _GEN1321 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1322 = io_x[3] ? _GEN1321 : _GEN66;
wire  _GEN1323 = io_x[7] ? _GEN1322 : _GEN65;
wire  _GEN1324 = io_x[23] ? _GEN81 : _GEN1323;
wire  _GEN1325 = io_x[2] ? _GEN140 : _GEN1324;
wire  _GEN1326 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1327 = io_x[3] ? _GEN1326 : _GEN66;
wire  _GEN1328 = io_x[7] ? _GEN1327 : _GEN65;
wire  _GEN1329 = io_x[23] ? _GEN81 : _GEN1328;
wire  _GEN1330 = io_x[2] ? _GEN1329 : _GEN573;
wire  _GEN1331 = io_x[16] ? _GEN1330 : _GEN1325;
wire  _GEN1332 = 1'b0;
wire  _GEN1333 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1334 = io_x[3] ? _GEN1333 : _GEN66;
wire  _GEN1335 = io_x[7] ? _GEN1334 : _GEN65;
wire  _GEN1336 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1337 = io_x[11] ? _GEN1336 : _GEN67;
wire  _GEN1338 = io_x[3] ? _GEN1337 : _GEN66;
wire  _GEN1339 = io_x[7] ? _GEN1338 : _GEN65;
wire  _GEN1340 = io_x[23] ? _GEN1339 : _GEN1335;
wire  _GEN1341 = io_x[2] ? _GEN1340 : _GEN573;
wire  _GEN1342 = io_x[16] ? _GEN1341 : _GEN1332;
wire  _GEN1343 = io_x[15] ? _GEN1342 : _GEN1331;
wire  _GEN1344 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1345 = io_x[7] ? _GEN1344 : _GEN65;
wire  _GEN1346 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1347 = io_x[3] ? _GEN78 : _GEN1346;
wire  _GEN1348 = io_x[7] ? _GEN1347 : _GEN65;
wire  _GEN1349 = io_x[23] ? _GEN1348 : _GEN1345;
wire  _GEN1350 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN1351 = io_x[2] ? _GEN1350 : _GEN1349;
wire  _GEN1352 = io_x[16] ? _GEN1351 : _GEN1240;
wire  _GEN1353 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1354 = io_x[23] ? _GEN81 : _GEN1353;
wire  _GEN1355 = io_x[23] ? _GEN81 : _GEN74;
wire  _GEN1356 = io_x[2] ? _GEN1355 : _GEN1354;
wire  _GEN1357 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1358 = io_x[7] ? _GEN1357 : _GEN65;
wire  _GEN1359 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1360 = io_x[11] ? _GEN1359 : _GEN76;
wire  _GEN1361 = io_x[3] ? _GEN66 : _GEN1360;
wire  _GEN1362 = io_x[7] ? _GEN1361 : _GEN65;
wire  _GEN1363 = io_x[23] ? _GEN1362 : _GEN1358;
wire  _GEN1364 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1365 = io_x[3] ? _GEN1364 : _GEN66;
wire  _GEN1366 = io_x[7] ? _GEN1365 : _GEN84;
wire  _GEN1367 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1368 = io_x[11] ? _GEN76 : _GEN1367;
wire  _GEN1369 = io_x[3] ? _GEN1368 : _GEN66;
wire  _GEN1370 = io_x[7] ? _GEN1369 : _GEN84;
wire  _GEN1371 = io_x[23] ? _GEN1370 : _GEN1366;
wire  _GEN1372 = io_x[2] ? _GEN1371 : _GEN1363;
wire  _GEN1373 = io_x[16] ? _GEN1372 : _GEN1356;
wire  _GEN1374 = io_x[15] ? _GEN1373 : _GEN1352;
wire  _GEN1375 = io_x[12] ? _GEN1374 : _GEN1343;
wire  _GEN1376 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1377 = io_x[3] ? _GEN66 : _GEN1376;
wire  _GEN1378 = io_x[7] ? _GEN1377 : _GEN84;
wire  _GEN1379 = io_x[23] ? _GEN74 : _GEN1378;
wire  _GEN1380 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1381 = io_x[23] ? _GEN81 : _GEN1380;
wire  _GEN1382 = io_x[2] ? _GEN1381 : _GEN1379;
wire  _GEN1383 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1384 = io_x[23] ? _GEN1383 : _GEN81;
wire  _GEN1385 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1386 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1387 = io_x[3] ? _GEN1386 : _GEN66;
wire  _GEN1388 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1389 = io_x[11] ? _GEN1388 : _GEN67;
wire  _GEN1390 = io_x[3] ? _GEN1389 : _GEN66;
wire  _GEN1391 = io_x[7] ? _GEN1390 : _GEN1387;
wire  _GEN1392 = io_x[23] ? _GEN1391 : _GEN1385;
wire  _GEN1393 = io_x[2] ? _GEN1392 : _GEN1384;
wire  _GEN1394 = io_x[16] ? _GEN1393 : _GEN1382;
wire  _GEN1395 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1396 = io_x[23] ? _GEN81 : _GEN1395;
wire  _GEN1397 = io_x[2] ? _GEN573 : _GEN1396;
wire  _GEN1398 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1399 = io_x[3] ? _GEN66 : _GEN1398;
wire  _GEN1400 = io_x[7] ? _GEN1399 : _GEN65;
wire  _GEN1401 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1402 = io_x[23] ? _GEN1401 : _GEN1400;
wire  _GEN1403 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1404 = io_x[11] ? _GEN1403 : _GEN67;
wire  _GEN1405 = io_x[3] ? _GEN1404 : _GEN66;
wire  _GEN1406 = io_x[7] ? _GEN1405 : _GEN65;
wire  _GEN1407 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1408 = io_x[11] ? _GEN1407 : _GEN67;
wire  _GEN1409 = io_x[3] ? _GEN1408 : _GEN66;
wire  _GEN1410 = io_x[7] ? _GEN1409 : _GEN65;
wire  _GEN1411 = io_x[23] ? _GEN1410 : _GEN1406;
wire  _GEN1412 = io_x[2] ? _GEN1411 : _GEN1402;
wire  _GEN1413 = io_x[16] ? _GEN1412 : _GEN1397;
wire  _GEN1414 = io_x[15] ? _GEN1413 : _GEN1394;
wire  _GEN1415 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1416 = io_x[7] ? _GEN1415 : _GEN65;
wire  _GEN1417 = io_x[23] ? _GEN81 : _GEN1416;
wire  _GEN1418 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1419 = io_x[23] ? _GEN81 : _GEN1418;
wire  _GEN1420 = io_x[2] ? _GEN1419 : _GEN1417;
wire  _GEN1421 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1422 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1423 = io_x[7] ? _GEN84 : _GEN1422;
wire  _GEN1424 = io_x[23] ? _GEN1423 : _GEN1421;
wire  _GEN1425 = io_x[2] ? _GEN1424 : _GEN140;
wire  _GEN1426 = io_x[16] ? _GEN1425 : _GEN1420;
wire  _GEN1427 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1428 = io_x[7] ? _GEN1427 : _GEN65;
wire  _GEN1429 = io_x[23] ? _GEN74 : _GEN1428;
wire  _GEN1430 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1431 = io_x[23] ? _GEN1430 : _GEN81;
wire  _GEN1432 = io_x[2] ? _GEN1431 : _GEN1429;
wire  _GEN1433 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1434 = io_x[7] ? _GEN1433 : _GEN65;
wire  _GEN1435 = io_x[23] ? _GEN1434 : _GEN81;
wire  _GEN1436 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1437 = io_x[3] ? _GEN1436 : _GEN78;
wire  _GEN1438 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1439 = io_x[11] ? _GEN1438 : _GEN67;
wire  _GEN1440 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1441 = io_x[11] ? _GEN1440 : _GEN67;
wire  _GEN1442 = io_x[3] ? _GEN1441 : _GEN1439;
wire  _GEN1443 = io_x[7] ? _GEN1442 : _GEN1437;
wire  _GEN1444 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1445 = io_x[11] ? _GEN1444 : _GEN67;
wire  _GEN1446 = io_x[3] ? _GEN1445 : _GEN78;
wire  _GEN1447 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1448 = io_x[11] ? _GEN1447 : _GEN67;
wire  _GEN1449 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1450 = io_x[11] ? _GEN1449 : _GEN67;
wire  _GEN1451 = io_x[3] ? _GEN1450 : _GEN1448;
wire  _GEN1452 = io_x[7] ? _GEN1451 : _GEN1446;
wire  _GEN1453 = io_x[23] ? _GEN1452 : _GEN1443;
wire  _GEN1454 = io_x[2] ? _GEN1453 : _GEN1435;
wire  _GEN1455 = io_x[16] ? _GEN1454 : _GEN1432;
wire  _GEN1456 = io_x[15] ? _GEN1455 : _GEN1426;
wire  _GEN1457 = io_x[12] ? _GEN1456 : _GEN1414;
wire  _GEN1458 = io_x[10] ? _GEN1457 : _GEN1375;
wire  _GEN1459 = io_x[4] ? _GEN1458 : _GEN1320;
wire  _GEN1460 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1461 = io_x[23] ? _GEN1460 : _GEN74;
wire  _GEN1462 = io_x[2] ? _GEN1461 : _GEN140;
wire  _GEN1463 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1464 = io_x[7] ? _GEN65 : _GEN1463;
wire  _GEN1465 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1466 = io_x[7] ? _GEN65 : _GEN1465;
wire  _GEN1467 = io_x[23] ? _GEN1466 : _GEN1464;
wire  _GEN1468 = io_x[2] ? _GEN1467 : _GEN140;
wire  _GEN1469 = io_x[16] ? _GEN1468 : _GEN1462;
wire  _GEN1470 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN1471 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1472 = io_x[23] ? _GEN1471 : _GEN81;
wire  _GEN1473 = io_x[2] ? _GEN1472 : _GEN1470;
wire  _GEN1474 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1475 = io_x[3] ? _GEN78 : _GEN1474;
wire  _GEN1476 = io_x[7] ? _GEN65 : _GEN1475;
wire  _GEN1477 = io_x[23] ? _GEN1476 : _GEN81;
wire  _GEN1478 = io_x[2] ? _GEN1477 : _GEN140;
wire  _GEN1479 = io_x[16] ? _GEN1478 : _GEN1473;
wire  _GEN1480 = io_x[15] ? _GEN1479 : _GEN1469;
wire  _GEN1481 = io_x[23] ? _GEN81 : _GEN74;
wire  _GEN1482 = io_x[2] ? _GEN1481 : _GEN573;
wire  _GEN1483 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1484 = io_x[7] ? _GEN84 : _GEN1483;
wire  _GEN1485 = io_x[23] ? _GEN1484 : _GEN81;
wire  _GEN1486 = io_x[2] ? _GEN1485 : _GEN573;
wire  _GEN1487 = io_x[16] ? _GEN1486 : _GEN1482;
wire  _GEN1488 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN1489 = io_x[2] ? _GEN1488 : _GEN573;
wire  _GEN1490 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1491 = io_x[3] ? _GEN1490 : _GEN78;
wire  _GEN1492 = io_x[7] ? _GEN84 : _GEN1491;
wire  _GEN1493 = io_x[23] ? _GEN1492 : _GEN81;
wire  _GEN1494 = io_x[2] ? _GEN1493 : _GEN140;
wire  _GEN1495 = io_x[16] ? _GEN1494 : _GEN1489;
wire  _GEN1496 = io_x[15] ? _GEN1495 : _GEN1487;
wire  _GEN1497 = io_x[12] ? _GEN1496 : _GEN1480;
wire  _GEN1498 = io_x[23] ? _GEN81 : _GEN74;
wire  _GEN1499 = io_x[2] ? _GEN1498 : _GEN140;
wire  _GEN1500 = io_x[16] ? _GEN1332 : _GEN1499;
wire  _GEN1501 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1502 = io_x[3] ? _GEN1501 : _GEN66;
wire  _GEN1503 = io_x[7] ? _GEN1502 : _GEN65;
wire  _GEN1504 = io_x[23] ? _GEN81 : _GEN1503;
wire  _GEN1505 = io_x[2] ? _GEN1504 : _GEN140;
wire  _GEN1506 = io_x[16] ? _GEN1505 : _GEN1240;
wire  _GEN1507 = io_x[15] ? _GEN1506 : _GEN1500;
wire  _GEN1508 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1509 = io_x[3] ? _GEN66 : _GEN1508;
wire  _GEN1510 = io_x[7] ? _GEN65 : _GEN1509;
wire  _GEN1511 = io_x[23] ? _GEN81 : _GEN1510;
wire  _GEN1512 = io_x[2] ? _GEN1511 : _GEN573;
wire  _GEN1513 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1514 = io_x[11] ? _GEN1513 : _GEN67;
wire  _GEN1515 = io_x[3] ? _GEN1514 : _GEN66;
wire  _GEN1516 = io_x[7] ? _GEN1515 : _GEN84;
wire  _GEN1517 = io_x[23] ? _GEN81 : _GEN1516;
wire  _GEN1518 = io_x[2] ? _GEN1517 : _GEN573;
wire  _GEN1519 = io_x[16] ? _GEN1518 : _GEN1512;
wire  _GEN1520 = io_x[23] ? _GEN81 : _GEN74;
wire  _GEN1521 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1522 = io_x[7] ? _GEN1521 : _GEN65;
wire  _GEN1523 = io_x[23] ? _GEN1522 : _GEN74;
wire  _GEN1524 = io_x[2] ? _GEN1523 : _GEN1520;
wire  _GEN1525 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1526 = io_x[7] ? _GEN1525 : _GEN65;
wire  _GEN1527 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1528 = io_x[11] ? _GEN1527 : _GEN67;
wire  _GEN1529 = io_x[3] ? _GEN1528 : _GEN78;
wire  _GEN1530 = io_x[7] ? _GEN1529 : _GEN84;
wire  _GEN1531 = io_x[23] ? _GEN1530 : _GEN1526;
wire  _GEN1532 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1533 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1534 = io_x[11] ? _GEN1533 : _GEN67;
wire  _GEN1535 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1536 = io_x[11] ? _GEN1535 : _GEN67;
wire  _GEN1537 = io_x[3] ? _GEN1536 : _GEN1534;
wire  _GEN1538 = io_x[7] ? _GEN1537 : _GEN1532;
wire  _GEN1539 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1540 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1541 = io_x[11] ? _GEN1540 : _GEN67;
wire  _GEN1542 = io_x[3] ? _GEN78 : _GEN1541;
wire  _GEN1543 = io_x[7] ? _GEN1542 : _GEN1539;
wire  _GEN1544 = io_x[23] ? _GEN1543 : _GEN1538;
wire  _GEN1545 = io_x[2] ? _GEN1544 : _GEN1531;
wire  _GEN1546 = io_x[16] ? _GEN1545 : _GEN1524;
wire  _GEN1547 = io_x[15] ? _GEN1546 : _GEN1519;
wire  _GEN1548 = io_x[12] ? _GEN1547 : _GEN1507;
wire  _GEN1549 = io_x[10] ? _GEN1548 : _GEN1497;
wire  _GEN1550 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1551 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1552 = io_x[23] ? _GEN1551 : _GEN1550;
wire  _GEN1553 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN1554 = io_x[2] ? _GEN1553 : _GEN1552;
wire  _GEN1555 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1556 = io_x[23] ? _GEN81 : _GEN1555;
wire  _GEN1557 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN1558 = io_x[2] ? _GEN1557 : _GEN1556;
wire  _GEN1559 = io_x[16] ? _GEN1558 : _GEN1554;
wire  _GEN1560 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1561 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1562 = io_x[23] ? _GEN1561 : _GEN1560;
wire  _GEN1563 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1564 = io_x[23] ? _GEN1563 : _GEN74;
wire  _GEN1565 = io_x[2] ? _GEN1564 : _GEN1562;
wire  _GEN1566 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1567 = io_x[23] ? _GEN81 : _GEN1566;
wire  _GEN1568 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1569 = io_x[11] ? _GEN1568 : _GEN76;
wire  _GEN1570 = io_x[3] ? _GEN1569 : _GEN66;
wire  _GEN1571 = io_x[7] ? _GEN1570 : _GEN65;
wire  _GEN1572 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1573 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1574 = io_x[11] ? _GEN1573 : _GEN1572;
wire  _GEN1575 = io_x[3] ? _GEN1574 : _GEN66;
wire  _GEN1576 = io_x[7] ? _GEN1575 : _GEN65;
wire  _GEN1577 = io_x[23] ? _GEN1576 : _GEN1571;
wire  _GEN1578 = io_x[2] ? _GEN1577 : _GEN1567;
wire  _GEN1579 = io_x[16] ? _GEN1578 : _GEN1565;
wire  _GEN1580 = io_x[15] ? _GEN1579 : _GEN1559;
wire  _GEN1581 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1582 = io_x[3] ? _GEN66 : _GEN1581;
wire  _GEN1583 = io_x[7] ? _GEN84 : _GEN1582;
wire  _GEN1584 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1585 = io_x[23] ? _GEN1584 : _GEN1583;
wire  _GEN1586 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1587 = io_x[7] ? _GEN1586 : _GEN84;
wire  _GEN1588 = io_x[23] ? _GEN81 : _GEN1587;
wire  _GEN1589 = io_x[2] ? _GEN1588 : _GEN1585;
wire  _GEN1590 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1591 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1592 = io_x[11] ? _GEN67 : _GEN1591;
wire  _GEN1593 = io_x[3] ? _GEN78 : _GEN1592;
wire  _GEN1594 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1595 = io_x[11] ? _GEN1594 : _GEN67;
wire  _GEN1596 = io_x[3] ? _GEN1595 : _GEN78;
wire  _GEN1597 = io_x[7] ? _GEN1596 : _GEN1593;
wire  _GEN1598 = io_x[23] ? _GEN1597 : _GEN1590;
wire  _GEN1599 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1600 = io_x[11] ? _GEN1599 : _GEN67;
wire  _GEN1601 = io_x[3] ? _GEN66 : _GEN1600;
wire  _GEN1602 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1603 = io_x[3] ? _GEN1602 : _GEN66;
wire  _GEN1604 = io_x[7] ? _GEN1603 : _GEN1601;
wire  _GEN1605 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1606 = io_x[3] ? _GEN1605 : _GEN66;
wire  _GEN1607 = io_x[7] ? _GEN1606 : _GEN65;
wire  _GEN1608 = io_x[23] ? _GEN1607 : _GEN1604;
wire  _GEN1609 = io_x[2] ? _GEN1608 : _GEN1598;
wire  _GEN1610 = io_x[16] ? _GEN1609 : _GEN1589;
wire  _GEN1611 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1612 = io_x[7] ? _GEN1611 : _GEN84;
wire  _GEN1613 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1614 = io_x[23] ? _GEN1613 : _GEN1612;
wire  _GEN1615 = io_x[23] ? _GEN81 : _GEN74;
wire  _GEN1616 = io_x[2] ? _GEN1615 : _GEN1614;
wire  _GEN1617 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1618 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1619 = io_x[11] ? _GEN1618 : _GEN67;
wire  _GEN1620 = io_x[3] ? _GEN1619 : _GEN66;
wire  _GEN1621 = io_x[7] ? _GEN1620 : _GEN84;
wire  _GEN1622 = io_x[23] ? _GEN1621 : _GEN1617;
wire  _GEN1623 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1624 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1625 = io_x[11] ? _GEN1624 : _GEN1623;
wire  _GEN1626 = io_x[3] ? _GEN1625 : _GEN66;
wire  _GEN1627 = io_x[7] ? _GEN1626 : _GEN84;
wire  _GEN1628 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1629 = io_x[11] ? _GEN1628 : _GEN67;
wire  _GEN1630 = io_x[3] ? _GEN1629 : _GEN66;
wire  _GEN1631 = io_x[7] ? _GEN1630 : _GEN65;
wire  _GEN1632 = io_x[23] ? _GEN1631 : _GEN1627;
wire  _GEN1633 = io_x[2] ? _GEN1632 : _GEN1622;
wire  _GEN1634 = io_x[16] ? _GEN1633 : _GEN1616;
wire  _GEN1635 = io_x[15] ? _GEN1634 : _GEN1610;
wire  _GEN1636 = io_x[12] ? _GEN1635 : _GEN1580;
wire  _GEN1637 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1638 = io_x[11] ? _GEN1637 : _GEN67;
wire  _GEN1639 = io_x[3] ? _GEN1638 : _GEN66;
wire  _GEN1640 = io_x[7] ? _GEN1639 : _GEN65;
wire  _GEN1641 = io_x[23] ? _GEN74 : _GEN1640;
wire  _GEN1642 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1643 = io_x[7] ? _GEN65 : _GEN1642;
wire  _GEN1644 = io_x[23] ? _GEN1643 : _GEN81;
wire  _GEN1645 = io_x[2] ? _GEN1644 : _GEN1641;
wire  _GEN1646 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1647 = io_x[3] ? _GEN1646 : _GEN66;
wire  _GEN1648 = io_x[7] ? _GEN1647 : _GEN84;
wire  _GEN1649 = io_x[23] ? _GEN1648 : _GEN81;
wire  _GEN1650 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1651 = io_x[11] ? _GEN1650 : _GEN67;
wire  _GEN1652 = io_x[3] ? _GEN1651 : _GEN66;
wire  _GEN1653 = io_x[7] ? _GEN1652 : _GEN84;
wire  _GEN1654 = io_x[23] ? _GEN81 : _GEN1653;
wire  _GEN1655 = io_x[2] ? _GEN1654 : _GEN1649;
wire  _GEN1656 = io_x[16] ? _GEN1655 : _GEN1645;
wire  _GEN1657 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1658 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1659 = io_x[23] ? _GEN1658 : _GEN1657;
wire  _GEN1660 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1661 = io_x[3] ? _GEN1660 : _GEN66;
wire  _GEN1662 = io_x[7] ? _GEN1661 : _GEN65;
wire  _GEN1663 = io_x[23] ? _GEN1662 : _GEN74;
wire  _GEN1664 = io_x[2] ? _GEN1663 : _GEN1659;
wire  _GEN1665 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1666 = io_x[7] ? _GEN65 : _GEN1665;
wire  _GEN1667 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1668 = io_x[11] ? _GEN1667 : _GEN67;
wire  _GEN1669 = io_x[3] ? _GEN1668 : _GEN66;
wire  _GEN1670 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1671 = io_x[11] ? _GEN1670 : _GEN67;
wire  _GEN1672 = io_x[3] ? _GEN1671 : _GEN66;
wire  _GEN1673 = io_x[7] ? _GEN1672 : _GEN1669;
wire  _GEN1674 = io_x[23] ? _GEN1673 : _GEN1666;
wire  _GEN1675 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1676 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1677 = io_x[11] ? _GEN1676 : _GEN1675;
wire  _GEN1678 = io_x[3] ? _GEN1677 : _GEN66;
wire  _GEN1679 = io_x[7] ? _GEN1678 : _GEN84;
wire  _GEN1680 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1681 = io_x[11] ? _GEN1680 : _GEN67;
wire  _GEN1682 = io_x[3] ? _GEN1681 : _GEN78;
wire  _GEN1683 = io_x[7] ? _GEN1682 : _GEN84;
wire  _GEN1684 = io_x[23] ? _GEN1683 : _GEN1679;
wire  _GEN1685 = io_x[2] ? _GEN1684 : _GEN1674;
wire  _GEN1686 = io_x[16] ? _GEN1685 : _GEN1664;
wire  _GEN1687 = io_x[15] ? _GEN1686 : _GEN1656;
wire  _GEN1688 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1689 = io_x[3] ? _GEN66 : _GEN1688;
wire  _GEN1690 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1691 = io_x[3] ? _GEN66 : _GEN1690;
wire  _GEN1692 = io_x[7] ? _GEN1691 : _GEN1689;
wire  _GEN1693 = io_x[23] ? _GEN81 : _GEN1692;
wire  _GEN1694 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1695 = io_x[11] ? _GEN67 : _GEN1694;
wire  _GEN1696 = io_x[3] ? _GEN1695 : _GEN78;
wire  _GEN1697 = io_x[7] ? _GEN1696 : _GEN65;
wire  _GEN1698 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1699 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1700 = io_x[11] ? _GEN1699 : _GEN1698;
wire  _GEN1701 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1702 = io_x[11] ? _GEN1701 : _GEN76;
wire  _GEN1703 = io_x[3] ? _GEN1702 : _GEN1700;
wire  _GEN1704 = io_x[7] ? _GEN1703 : _GEN65;
wire  _GEN1705 = io_x[23] ? _GEN1704 : _GEN1697;
wire  _GEN1706 = io_x[2] ? _GEN1705 : _GEN1693;
wire  _GEN1707 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1708 = io_x[3] ? _GEN78 : _GEN1707;
wire  _GEN1709 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1710 = io_x[11] ? _GEN76 : _GEN1709;
wire  _GEN1711 = io_x[3] ? _GEN1710 : _GEN66;
wire  _GEN1712 = io_x[7] ? _GEN1711 : _GEN1708;
wire  _GEN1713 = io_x[23] ? _GEN1712 : _GEN74;
wire  _GEN1714 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1715 = io_x[11] ? _GEN67 : _GEN1714;
wire  _GEN1716 = io_x[3] ? _GEN1715 : _GEN66;
wire  _GEN1717 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1718 = io_x[11] ? _GEN76 : _GEN1717;
wire  _GEN1719 = io_x[3] ? _GEN1718 : _GEN66;
wire  _GEN1720 = io_x[7] ? _GEN1719 : _GEN1716;
wire  _GEN1721 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1722 = io_x[11] ? _GEN67 : _GEN1721;
wire  _GEN1723 = io_x[3] ? _GEN1722 : _GEN66;
wire  _GEN1724 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1725 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1726 = io_x[11] ? _GEN1725 : _GEN1724;
wire  _GEN1727 = io_x[3] ? _GEN1726 : _GEN78;
wire  _GEN1728 = io_x[7] ? _GEN1727 : _GEN1723;
wire  _GEN1729 = io_x[23] ? _GEN1728 : _GEN1720;
wire  _GEN1730 = io_x[2] ? _GEN1729 : _GEN1713;
wire  _GEN1731 = io_x[16] ? _GEN1730 : _GEN1706;
wire  _GEN1732 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1733 = io_x[3] ? _GEN66 : _GEN1732;
wire  _GEN1734 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1735 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1736 = io_x[11] ? _GEN1735 : _GEN67;
wire  _GEN1737 = io_x[3] ? _GEN1736 : _GEN1734;
wire  _GEN1738 = io_x[7] ? _GEN1737 : _GEN1733;
wire  _GEN1739 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1740 = io_x[3] ? _GEN1739 : _GEN78;
wire  _GEN1741 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1742 = io_x[11] ? _GEN1741 : _GEN67;
wire  _GEN1743 = io_x[3] ? _GEN1742 : _GEN66;
wire  _GEN1744 = io_x[7] ? _GEN1743 : _GEN1740;
wire  _GEN1745 = io_x[23] ? _GEN1744 : _GEN1738;
wire  _GEN1746 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1747 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1748 = io_x[11] ? _GEN1747 : _GEN1746;
wire  _GEN1749 = io_x[3] ? _GEN1748 : _GEN66;
wire  _GEN1750 = io_x[7] ? _GEN1749 : _GEN65;
wire  _GEN1751 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1752 = io_x[11] ? _GEN76 : _GEN1751;
wire  _GEN1753 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1754 = io_x[11] ? _GEN1753 : _GEN67;
wire  _GEN1755 = io_x[3] ? _GEN1754 : _GEN1752;
wire  _GEN1756 = io_x[7] ? _GEN1755 : _GEN84;
wire  _GEN1757 = io_x[23] ? _GEN1756 : _GEN1750;
wire  _GEN1758 = io_x[2] ? _GEN1757 : _GEN1745;
wire  _GEN1759 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1760 = io_x[3] ? _GEN78 : _GEN1759;
wire  _GEN1761 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1762 = io_x[11] ? _GEN1761 : _GEN67;
wire  _GEN1763 = io_x[3] ? _GEN1762 : _GEN78;
wire  _GEN1764 = io_x[7] ? _GEN1763 : _GEN1760;
wire  _GEN1765 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1766 = io_x[3] ? _GEN1765 : _GEN66;
wire  _GEN1767 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1768 = io_x[11] ? _GEN1767 : _GEN67;
wire  _GEN1769 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1770 = io_x[11] ? _GEN1769 : _GEN67;
wire  _GEN1771 = io_x[3] ? _GEN1770 : _GEN1768;
wire  _GEN1772 = io_x[7] ? _GEN1771 : _GEN1766;
wire  _GEN1773 = io_x[23] ? _GEN1772 : _GEN1764;
wire  _GEN1774 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1775 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1776 = io_x[11] ? _GEN1775 : _GEN1774;
wire  _GEN1777 = io_x[3] ? _GEN1776 : _GEN78;
wire  _GEN1778 = io_x[7] ? _GEN1777 : _GEN84;
wire  _GEN1779 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1780 = io_x[11] ? _GEN1779 : _GEN67;
wire  _GEN1781 = io_x[3] ? _GEN1780 : _GEN78;
wire  _GEN1782 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1783 = io_x[11] ? _GEN1782 : _GEN67;
wire  _GEN1784 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1785 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1786 = io_x[11] ? _GEN1785 : _GEN1784;
wire  _GEN1787 = io_x[3] ? _GEN1786 : _GEN1783;
wire  _GEN1788 = io_x[7] ? _GEN1787 : _GEN1781;
wire  _GEN1789 = io_x[23] ? _GEN1788 : _GEN1778;
wire  _GEN1790 = io_x[2] ? _GEN1789 : _GEN1773;
wire  _GEN1791 = io_x[16] ? _GEN1790 : _GEN1758;
wire  _GEN1792 = io_x[15] ? _GEN1791 : _GEN1731;
wire  _GEN1793 = io_x[12] ? _GEN1792 : _GEN1687;
wire  _GEN1794 = io_x[10] ? _GEN1793 : _GEN1636;
wire  _GEN1795 = io_x[4] ? _GEN1794 : _GEN1549;
wire  _GEN1796 = io_x[8] ? _GEN1795 : _GEN1459;
wire  _GEN1797 = io_x[28] ? _GEN1796 : _GEN1211;
wire  _GEN1798 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1799 = io_x[23] ? _GEN1798 : _GEN74;
wire  _GEN1800 = io_x[2] ? _GEN573 : _GEN1799;
wire  _GEN1801 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1802 = io_x[11] ? _GEN1801 : _GEN76;
wire  _GEN1803 = io_x[3] ? _GEN1802 : _GEN78;
wire  _GEN1804 = io_x[7] ? _GEN1803 : _GEN65;
wire  _GEN1805 = io_x[23] ? _GEN81 : _GEN1804;
wire  _GEN1806 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1807 = io_x[11] ? _GEN1806 : _GEN76;
wire  _GEN1808 = io_x[3] ? _GEN1807 : _GEN66;
wire  _GEN1809 = io_x[7] ? _GEN1808 : _GEN65;
wire  _GEN1810 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1811 = io_x[23] ? _GEN1810 : _GEN1809;
wire  _GEN1812 = io_x[2] ? _GEN1811 : _GEN1805;
wire  _GEN1813 = io_x[16] ? _GEN1812 : _GEN1800;
wire  _GEN1814 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1815 = io_x[11] ? _GEN1814 : _GEN67;
wire  _GEN1816 = io_x[3] ? _GEN1815 : _GEN66;
wire  _GEN1817 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1818 = io_x[3] ? _GEN1817 : _GEN66;
wire  _GEN1819 = io_x[7] ? _GEN1818 : _GEN1816;
wire  _GEN1820 = io_x[23] ? _GEN74 : _GEN1819;
wire  _GEN1821 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1822 = io_x[23] ? _GEN1821 : _GEN74;
wire  _GEN1823 = io_x[2] ? _GEN1822 : _GEN1820;
wire  _GEN1824 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1825 = io_x[11] ? _GEN1824 : _GEN67;
wire  _GEN1826 = io_x[3] ? _GEN1825 : _GEN66;
wire  _GEN1827 = io_x[7] ? _GEN1826 : _GEN65;
wire  _GEN1828 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1829 = io_x[11] ? _GEN1828 : _GEN76;
wire  _GEN1830 = io_x[3] ? _GEN1829 : _GEN66;
wire  _GEN1831 = io_x[7] ? _GEN1830 : _GEN84;
wire  _GEN1832 = io_x[23] ? _GEN1831 : _GEN1827;
wire  _GEN1833 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1834 = io_x[11] ? _GEN1833 : _GEN67;
wire  _GEN1835 = io_x[3] ? _GEN1834 : _GEN66;
wire  _GEN1836 = io_x[7] ? _GEN1835 : _GEN84;
wire  _GEN1837 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1838 = io_x[11] ? _GEN1837 : _GEN67;
wire  _GEN1839 = io_x[3] ? _GEN1838 : _GEN66;
wire  _GEN1840 = io_x[7] ? _GEN1839 : _GEN65;
wire  _GEN1841 = io_x[23] ? _GEN1840 : _GEN1836;
wire  _GEN1842 = io_x[2] ? _GEN1841 : _GEN1832;
wire  _GEN1843 = io_x[16] ? _GEN1842 : _GEN1823;
wire  _GEN1844 = io_x[15] ? _GEN1843 : _GEN1813;
wire  _GEN1845 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN1846 = io_x[2] ? _GEN573 : _GEN1845;
wire  _GEN1847 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1848 = io_x[3] ? _GEN1847 : _GEN66;
wire  _GEN1849 = io_x[7] ? _GEN84 : _GEN1848;
wire  _GEN1850 = io_x[23] ? _GEN81 : _GEN1849;
wire  _GEN1851 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1852 = io_x[3] ? _GEN1851 : _GEN66;
wire  _GEN1853 = io_x[7] ? _GEN84 : _GEN1852;
wire  _GEN1854 = io_x[23] ? _GEN74 : _GEN1853;
wire  _GEN1855 = io_x[2] ? _GEN1854 : _GEN1850;
wire  _GEN1856 = io_x[16] ? _GEN1855 : _GEN1846;
wire  _GEN1857 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1858 = io_x[3] ? _GEN1857 : _GEN66;
wire  _GEN1859 = io_x[7] ? _GEN1858 : _GEN84;
wire  _GEN1860 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1861 = io_x[3] ? _GEN1860 : _GEN66;
wire  _GEN1862 = io_x[7] ? _GEN65 : _GEN1861;
wire  _GEN1863 = io_x[23] ? _GEN1862 : _GEN1859;
wire  _GEN1864 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1865 = io_x[3] ? _GEN1864 : _GEN66;
wire  _GEN1866 = io_x[7] ? _GEN1865 : _GEN84;
wire  _GEN1867 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN1868 = io_x[23] ? _GEN1867 : _GEN1866;
wire  _GEN1869 = io_x[2] ? _GEN1868 : _GEN1863;
wire  _GEN1870 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1871 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1872 = io_x[11] ? _GEN1871 : _GEN67;
wire  _GEN1873 = io_x[3] ? _GEN1872 : _GEN66;
wire  _GEN1874 = io_x[7] ? _GEN1873 : _GEN1870;
wire  _GEN1875 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1876 = io_x[11] ? _GEN76 : _GEN1875;
wire  _GEN1877 = io_x[3] ? _GEN1876 : _GEN66;
wire  _GEN1878 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1879 = io_x[3] ? _GEN1878 : _GEN66;
wire  _GEN1880 = io_x[7] ? _GEN1879 : _GEN1877;
wire  _GEN1881 = io_x[23] ? _GEN1880 : _GEN1874;
wire  _GEN1882 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1883 = io_x[11] ? _GEN1882 : _GEN67;
wire  _GEN1884 = io_x[3] ? _GEN1883 : _GEN78;
wire  _GEN1885 = io_x[7] ? _GEN1884 : _GEN65;
wire  _GEN1886 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1887 = io_x[11] ? _GEN76 : _GEN1886;
wire  _GEN1888 = io_x[3] ? _GEN1887 : _GEN66;
wire  _GEN1889 = io_x[7] ? _GEN65 : _GEN1888;
wire  _GEN1890 = io_x[23] ? _GEN1889 : _GEN1885;
wire  _GEN1891 = io_x[2] ? _GEN1890 : _GEN1881;
wire  _GEN1892 = io_x[16] ? _GEN1891 : _GEN1869;
wire  _GEN1893 = io_x[15] ? _GEN1892 : _GEN1856;
wire  _GEN1894 = io_x[12] ? _GEN1893 : _GEN1844;
wire  _GEN1895 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN1896 = io_x[2] ? _GEN140 : _GEN1895;
wire  _GEN1897 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1898 = io_x[11] ? _GEN1897 : _GEN67;
wire  _GEN1899 = io_x[3] ? _GEN1898 : _GEN66;
wire  _GEN1900 = io_x[7] ? _GEN1899 : _GEN65;
wire  _GEN1901 = io_x[23] ? _GEN74 : _GEN1900;
wire  _GEN1902 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1903 = io_x[7] ? _GEN1902 : _GEN65;
wire  _GEN1904 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN1905 = io_x[7] ? _GEN1904 : _GEN84;
wire  _GEN1906 = io_x[23] ? _GEN1905 : _GEN1903;
wire  _GEN1907 = io_x[2] ? _GEN1906 : _GEN1901;
wire  _GEN1908 = io_x[16] ? _GEN1907 : _GEN1896;
wire  _GEN1909 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1910 = io_x[3] ? _GEN1909 : _GEN66;
wire  _GEN1911 = io_x[7] ? _GEN1910 : _GEN84;
wire  _GEN1912 = io_x[23] ? _GEN81 : _GEN1911;
wire  _GEN1913 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1914 = io_x[11] ? _GEN1913 : _GEN67;
wire  _GEN1915 = io_x[3] ? _GEN1914 : _GEN66;
wire  _GEN1916 = io_x[7] ? _GEN1915 : _GEN65;
wire  _GEN1917 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1918 = io_x[3] ? _GEN1917 : _GEN66;
wire  _GEN1919 = io_x[7] ? _GEN1918 : _GEN84;
wire  _GEN1920 = io_x[23] ? _GEN1919 : _GEN1916;
wire  _GEN1921 = io_x[2] ? _GEN1920 : _GEN1912;
wire  _GEN1922 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1923 = io_x[11] ? _GEN1922 : _GEN67;
wire  _GEN1924 = io_x[3] ? _GEN1923 : _GEN66;
wire  _GEN1925 = io_x[7] ? _GEN1924 : _GEN65;
wire  _GEN1926 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1927 = io_x[3] ? _GEN66 : _GEN1926;
wire  _GEN1928 = io_x[7] ? _GEN65 : _GEN1927;
wire  _GEN1929 = io_x[23] ? _GEN1928 : _GEN1925;
wire  _GEN1930 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1931 = io_x[11] ? _GEN1930 : _GEN76;
wire  _GEN1932 = io_x[3] ? _GEN1931 : _GEN66;
wire  _GEN1933 = io_x[7] ? _GEN1932 : _GEN84;
wire  _GEN1934 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1935 = io_x[11] ? _GEN1934 : _GEN76;
wire  _GEN1936 = io_x[3] ? _GEN1935 : _GEN66;
wire  _GEN1937 = io_x[7] ? _GEN1936 : _GEN65;
wire  _GEN1938 = io_x[23] ? _GEN1937 : _GEN1933;
wire  _GEN1939 = io_x[2] ? _GEN1938 : _GEN1929;
wire  _GEN1940 = io_x[16] ? _GEN1939 : _GEN1921;
wire  _GEN1941 = io_x[15] ? _GEN1940 : _GEN1908;
wire  _GEN1942 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1943 = io_x[7] ? _GEN65 : _GEN1942;
wire  _GEN1944 = io_x[23] ? _GEN74 : _GEN1943;
wire  _GEN1945 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1946 = io_x[11] ? _GEN67 : _GEN1945;
wire  _GEN1947 = io_x[3] ? _GEN1946 : _GEN66;
wire  _GEN1948 = io_x[7] ? _GEN1947 : _GEN84;
wire  _GEN1949 = io_x[23] ? _GEN1948 : _GEN74;
wire  _GEN1950 = io_x[2] ? _GEN1949 : _GEN1944;
wire  _GEN1951 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1952 = io_x[11] ? _GEN67 : _GEN1951;
wire  _GEN1953 = io_x[3] ? _GEN1952 : _GEN66;
wire  _GEN1954 = io_x[7] ? _GEN1953 : _GEN65;
wire  _GEN1955 = io_x[23] ? _GEN81 : _GEN1954;
wire  _GEN1956 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1957 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1958 = io_x[11] ? _GEN1957 : _GEN1956;
wire  _GEN1959 = io_x[3] ? _GEN1958 : _GEN66;
wire  _GEN1960 = io_x[7] ? _GEN1959 : _GEN65;
wire  _GEN1961 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN1962 = io_x[11] ? _GEN67 : _GEN1961;
wire  _GEN1963 = io_x[3] ? _GEN1962 : _GEN66;
wire  _GEN1964 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1965 = io_x[7] ? _GEN1964 : _GEN1963;
wire  _GEN1966 = io_x[23] ? _GEN1965 : _GEN1960;
wire  _GEN1967 = io_x[2] ? _GEN1966 : _GEN1955;
wire  _GEN1968 = io_x[16] ? _GEN1967 : _GEN1950;
wire  _GEN1969 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1970 = io_x[3] ? _GEN1969 : _GEN66;
wire  _GEN1971 = io_x[7] ? _GEN1970 : _GEN65;
wire  _GEN1972 = io_x[23] ? _GEN74 : _GEN1971;
wire  _GEN1973 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1974 = io_x[3] ? _GEN1973 : _GEN66;
wire  _GEN1975 = io_x[7] ? _GEN1974 : _GEN65;
wire  _GEN1976 = io_x[23] ? _GEN1975 : _GEN74;
wire  _GEN1977 = io_x[2] ? _GEN1976 : _GEN1972;
wire  _GEN1978 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN1979 = io_x[3] ? _GEN1978 : _GEN66;
wire  _GEN1980 = io_x[7] ? _GEN1979 : _GEN65;
wire  _GEN1981 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN1982 = io_x[23] ? _GEN1981 : _GEN1980;
wire  _GEN1983 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1984 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN1985 = io_x[11] ? _GEN1984 : _GEN76;
wire  _GEN1986 = io_x[3] ? _GEN1985 : _GEN66;
wire  _GEN1987 = io_x[7] ? _GEN1986 : _GEN1983;
wire  _GEN1988 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN1989 = io_x[3] ? _GEN78 : _GEN1988;
wire  _GEN1990 = io_x[7] ? _GEN1989 : _GEN65;
wire  _GEN1991 = io_x[23] ? _GEN1990 : _GEN1987;
wire  _GEN1992 = io_x[2] ? _GEN1991 : _GEN1982;
wire  _GEN1993 = io_x[16] ? _GEN1992 : _GEN1977;
wire  _GEN1994 = io_x[15] ? _GEN1993 : _GEN1968;
wire  _GEN1995 = io_x[12] ? _GEN1994 : _GEN1941;
wire  _GEN1996 = io_x[10] ? _GEN1995 : _GEN1894;
wire  _GEN1997 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN1998 = io_x[7] ? _GEN1997 : _GEN84;
wire  _GEN1999 = io_x[23] ? _GEN74 : _GEN1998;
wire  _GEN2000 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN2001 = io_x[7] ? _GEN2000 : _GEN65;
wire  _GEN2002 = io_x[23] ? _GEN2001 : _GEN74;
wire  _GEN2003 = io_x[2] ? _GEN2002 : _GEN1999;
wire  _GEN2004 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2005 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2006 = io_x[3] ? _GEN2005 : _GEN66;
wire  _GEN2007 = io_x[7] ? _GEN2006 : _GEN84;
wire  _GEN2008 = io_x[23] ? _GEN2007 : _GEN2004;
wire  _GEN2009 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2010 = io_x[11] ? _GEN2009 : _GEN76;
wire  _GEN2011 = io_x[3] ? _GEN2010 : _GEN78;
wire  _GEN2012 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2013 = io_x[11] ? _GEN67 : _GEN2012;
wire  _GEN2014 = io_x[3] ? _GEN78 : _GEN2013;
wire  _GEN2015 = io_x[7] ? _GEN2014 : _GEN2011;
wire  _GEN2016 = io_x[23] ? _GEN2015 : _GEN81;
wire  _GEN2017 = io_x[2] ? _GEN2016 : _GEN2008;
wire  _GEN2018 = io_x[16] ? _GEN2017 : _GEN2003;
wire  _GEN2019 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN2020 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2021 = io_x[7] ? _GEN2020 : _GEN65;
wire  _GEN2022 = io_x[23] ? _GEN2021 : _GEN2019;
wire  _GEN2023 = io_x[2] ? _GEN140 : _GEN2022;
wire  _GEN2024 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2025 = io_x[11] ? _GEN2024 : _GEN67;
wire  _GEN2026 = io_x[3] ? _GEN2025 : _GEN66;
wire  _GEN2027 = io_x[7] ? _GEN2026 : _GEN65;
wire  _GEN2028 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN2029 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2030 = io_x[11] ? _GEN2029 : _GEN67;
wire  _GEN2031 = io_x[3] ? _GEN66 : _GEN2030;
wire  _GEN2032 = io_x[7] ? _GEN2031 : _GEN2028;
wire  _GEN2033 = io_x[23] ? _GEN2032 : _GEN2027;
wire  _GEN2034 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2035 = io_x[3] ? _GEN2034 : _GEN66;
wire  _GEN2036 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2037 = io_x[11] ? _GEN2036 : _GEN67;
wire  _GEN2038 = io_x[3] ? _GEN2037 : _GEN78;
wire  _GEN2039 = io_x[7] ? _GEN2038 : _GEN2035;
wire  _GEN2040 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2041 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2042 = io_x[11] ? _GEN2041 : _GEN67;
wire  _GEN2043 = io_x[3] ? _GEN2042 : _GEN78;
wire  _GEN2044 = io_x[7] ? _GEN2043 : _GEN2040;
wire  _GEN2045 = io_x[23] ? _GEN2044 : _GEN2039;
wire  _GEN2046 = io_x[2] ? _GEN2045 : _GEN2033;
wire  _GEN2047 = io_x[16] ? _GEN2046 : _GEN2023;
wire  _GEN2048 = io_x[15] ? _GEN2047 : _GEN2018;
wire  _GEN2049 = io_x[2] ? _GEN573 : _GEN140;
wire  _GEN2050 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN2051 = io_x[7] ? _GEN2050 : _GEN65;
wire  _GEN2052 = io_x[23] ? _GEN2051 : _GEN81;
wire  _GEN2053 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2054 = io_x[11] ? _GEN2053 : _GEN67;
wire  _GEN2055 = io_x[3] ? _GEN2054 : _GEN66;
wire  _GEN2056 = io_x[7] ? _GEN2055 : _GEN65;
wire  _GEN2057 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2058 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2059 = io_x[11] ? _GEN2058 : _GEN2057;
wire  _GEN2060 = io_x[3] ? _GEN2059 : _GEN66;
wire  _GEN2061 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2062 = io_x[11] ? _GEN2061 : _GEN76;
wire  _GEN2063 = io_x[3] ? _GEN2062 : _GEN66;
wire  _GEN2064 = io_x[7] ? _GEN2063 : _GEN2060;
wire  _GEN2065 = io_x[23] ? _GEN2064 : _GEN2056;
wire  _GEN2066 = io_x[2] ? _GEN2065 : _GEN2052;
wire  _GEN2067 = io_x[16] ? _GEN2066 : _GEN2049;
wire  _GEN2068 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2069 = io_x[3] ? _GEN78 : _GEN2068;
wire  _GEN2070 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2071 = io_x[11] ? _GEN2070 : _GEN67;
wire  _GEN2072 = io_x[3] ? _GEN66 : _GEN2071;
wire  _GEN2073 = io_x[7] ? _GEN2072 : _GEN2069;
wire  _GEN2074 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2075 = io_x[7] ? _GEN2074 : _GEN65;
wire  _GEN2076 = io_x[23] ? _GEN2075 : _GEN2073;
wire  _GEN2077 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2078 = io_x[23] ? _GEN81 : _GEN2077;
wire  _GEN2079 = io_x[2] ? _GEN2078 : _GEN2076;
wire  _GEN2080 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2081 = io_x[3] ? _GEN2080 : _GEN66;
wire  _GEN2082 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN2083 = io_x[7] ? _GEN2082 : _GEN2081;
wire  _GEN2084 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2085 = io_x[3] ? _GEN66 : _GEN2084;
wire  _GEN2086 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2087 = io_x[3] ? _GEN2086 : _GEN78;
wire  _GEN2088 = io_x[7] ? _GEN2087 : _GEN2085;
wire  _GEN2089 = io_x[23] ? _GEN2088 : _GEN2083;
wire  _GEN2090 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2091 = io_x[3] ? _GEN2090 : _GEN66;
wire  _GEN2092 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2093 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2094 = io_x[11] ? _GEN76 : _GEN2093;
wire  _GEN2095 = io_x[3] ? _GEN2094 : _GEN2092;
wire  _GEN2096 = io_x[7] ? _GEN2095 : _GEN2091;
wire  _GEN2097 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2098 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2099 = io_x[11] ? _GEN76 : _GEN2098;
wire  _GEN2100 = io_x[3] ? _GEN2099 : _GEN2097;
wire  _GEN2101 = io_x[7] ? _GEN2100 : _GEN84;
wire  _GEN2102 = io_x[23] ? _GEN2101 : _GEN2096;
wire  _GEN2103 = io_x[2] ? _GEN2102 : _GEN2089;
wire  _GEN2104 = io_x[16] ? _GEN2103 : _GEN2079;
wire  _GEN2105 = io_x[15] ? _GEN2104 : _GEN2067;
wire  _GEN2106 = io_x[12] ? _GEN2105 : _GEN2048;
wire  _GEN2107 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2108 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2109 = io_x[11] ? _GEN2108 : _GEN2107;
wire  _GEN2110 = io_x[3] ? _GEN66 : _GEN2109;
wire  _GEN2111 = io_x[7] ? _GEN2110 : _GEN84;
wire  _GEN2112 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN2113 = io_x[23] ? _GEN2112 : _GEN2111;
wire  _GEN2114 = io_x[2] ? _GEN140 : _GEN2113;
wire  _GEN2115 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2116 = io_x[11] ? _GEN76 : _GEN2115;
wire  _GEN2117 = io_x[3] ? _GEN2116 : _GEN78;
wire  _GEN2118 = io_x[7] ? _GEN65 : _GEN2117;
wire  _GEN2119 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2120 = io_x[3] ? _GEN66 : _GEN2119;
wire  _GEN2121 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2122 = io_x[7] ? _GEN2121 : _GEN2120;
wire  _GEN2123 = io_x[23] ? _GEN2122 : _GEN2118;
wire  _GEN2124 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2125 = io_x[11] ? _GEN2124 : _GEN67;
wire  _GEN2126 = io_x[3] ? _GEN2125 : _GEN78;
wire  _GEN2127 = io_x[7] ? _GEN2126 : _GEN65;
wire  _GEN2128 = io_x[23] ? _GEN2127 : _GEN74;
wire  _GEN2129 = io_x[2] ? _GEN2128 : _GEN2123;
wire  _GEN2130 = io_x[16] ? _GEN2129 : _GEN2114;
wire  _GEN2131 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2132 = io_x[23] ? _GEN2131 : _GEN81;
wire  _GEN2133 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2134 = io_x[23] ? _GEN81 : _GEN2133;
wire  _GEN2135 = io_x[2] ? _GEN2134 : _GEN2132;
wire  _GEN2136 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2137 = io_x[3] ? _GEN66 : _GEN2136;
wire  _GEN2138 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2139 = io_x[3] ? _GEN2138 : _GEN66;
wire  _GEN2140 = io_x[7] ? _GEN2139 : _GEN2137;
wire  _GEN2141 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2142 = io_x[3] ? _GEN66 : _GEN2141;
wire  _GEN2143 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2144 = io_x[3] ? _GEN2143 : _GEN66;
wire  _GEN2145 = io_x[7] ? _GEN2144 : _GEN2142;
wire  _GEN2146 = io_x[23] ? _GEN2145 : _GEN2140;
wire  _GEN2147 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2148 = io_x[11] ? _GEN2147 : _GEN67;
wire  _GEN2149 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2150 = io_x[11] ? _GEN2149 : _GEN67;
wire  _GEN2151 = io_x[3] ? _GEN2150 : _GEN2148;
wire  _GEN2152 = io_x[7] ? _GEN2151 : _GEN65;
wire  _GEN2153 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2154 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2155 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2156 = io_x[11] ? _GEN2155 : _GEN2154;
wire  _GEN2157 = io_x[3] ? _GEN2156 : _GEN2153;
wire  _GEN2158 = io_x[7] ? _GEN2157 : _GEN65;
wire  _GEN2159 = io_x[23] ? _GEN2158 : _GEN2152;
wire  _GEN2160 = io_x[2] ? _GEN2159 : _GEN2146;
wire  _GEN2161 = io_x[16] ? _GEN2160 : _GEN2135;
wire  _GEN2162 = io_x[15] ? _GEN2161 : _GEN2130;
wire  _GEN2163 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2164 = io_x[11] ? _GEN2163 : _GEN76;
wire  _GEN2165 = io_x[3] ? _GEN78 : _GEN2164;
wire  _GEN2166 = io_x[7] ? _GEN2165 : _GEN65;
wire  _GEN2167 = io_x[23] ? _GEN81 : _GEN2166;
wire  _GEN2168 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2169 = io_x[7] ? _GEN2168 : _GEN65;
wire  _GEN2170 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2171 = io_x[11] ? _GEN67 : _GEN2170;
wire  _GEN2172 = io_x[3] ? _GEN66 : _GEN2171;
wire  _GEN2173 = io_x[7] ? _GEN65 : _GEN2172;
wire  _GEN2174 = io_x[23] ? _GEN2173 : _GEN2169;
wire  _GEN2175 = io_x[2] ? _GEN2174 : _GEN2167;
wire  _GEN2176 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2177 = io_x[3] ? _GEN2176 : _GEN66;
wire  _GEN2178 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2179 = io_x[11] ? _GEN67 : _GEN2178;
wire  _GEN2180 = io_x[3] ? _GEN2179 : _GEN66;
wire  _GEN2181 = io_x[7] ? _GEN2180 : _GEN2177;
wire  _GEN2182 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2183 = io_x[23] ? _GEN2182 : _GEN2181;
wire  _GEN2184 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2185 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2186 = io_x[3] ? _GEN2185 : _GEN2184;
wire  _GEN2187 = io_x[7] ? _GEN2186 : _GEN65;
wire  _GEN2188 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2189 = io_x[3] ? _GEN2188 : _GEN78;
wire  _GEN2190 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2191 = io_x[7] ? _GEN2190 : _GEN2189;
wire  _GEN2192 = io_x[23] ? _GEN2191 : _GEN2187;
wire  _GEN2193 = io_x[2] ? _GEN2192 : _GEN2183;
wire  _GEN2194 = io_x[16] ? _GEN2193 : _GEN2175;
wire  _GEN2195 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2196 = io_x[3] ? _GEN2195 : _GEN78;
wire  _GEN2197 = io_x[7] ? _GEN2196 : _GEN84;
wire  _GEN2198 = io_x[23] ? _GEN74 : _GEN2197;
wire  _GEN2199 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2200 = io_x[11] ? _GEN2199 : _GEN67;
wire  _GEN2201 = io_x[3] ? _GEN2200 : _GEN66;
wire  _GEN2202 = io_x[7] ? _GEN2201 : _GEN84;
wire  _GEN2203 = io_x[23] ? _GEN81 : _GEN2202;
wire  _GEN2204 = io_x[2] ? _GEN2203 : _GEN2198;
wire  _GEN2205 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2206 = io_x[11] ? _GEN2205 : _GEN67;
wire  _GEN2207 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2208 = io_x[3] ? _GEN2207 : _GEN2206;
wire  _GEN2209 = io_x[7] ? _GEN2208 : _GEN65;
wire  _GEN2210 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2211 = io_x[7] ? _GEN84 : _GEN2210;
wire  _GEN2212 = io_x[23] ? _GEN2211 : _GEN2209;
wire  _GEN2213 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2214 = io_x[11] ? _GEN2213 : _GEN67;
wire  _GEN2215 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2216 = io_x[11] ? _GEN2215 : _GEN76;
wire  _GEN2217 = io_x[3] ? _GEN2216 : _GEN2214;
wire  _GEN2218 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2219 = io_x[11] ? _GEN2218 : _GEN67;
wire  _GEN2220 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2221 = io_x[3] ? _GEN2220 : _GEN2219;
wire  _GEN2222 = io_x[7] ? _GEN2221 : _GEN2217;
wire  _GEN2223 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2224 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2225 = io_x[11] ? _GEN2224 : _GEN76;
wire  _GEN2226 = io_x[3] ? _GEN2225 : _GEN2223;
wire  _GEN2227 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2228 = io_x[11] ? _GEN67 : _GEN2227;
wire  _GEN2229 = io_x[3] ? _GEN78 : _GEN2228;
wire  _GEN2230 = io_x[7] ? _GEN2229 : _GEN2226;
wire  _GEN2231 = io_x[23] ? _GEN2230 : _GEN2222;
wire  _GEN2232 = io_x[2] ? _GEN2231 : _GEN2212;
wire  _GEN2233 = io_x[16] ? _GEN2232 : _GEN2204;
wire  _GEN2234 = io_x[15] ? _GEN2233 : _GEN2194;
wire  _GEN2235 = io_x[12] ? _GEN2234 : _GEN2162;
wire  _GEN2236 = io_x[10] ? _GEN2235 : _GEN2106;
wire  _GEN2237 = io_x[4] ? _GEN2236 : _GEN1996;
wire  _GEN2238 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN2239 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2240 = io_x[11] ? _GEN2239 : _GEN67;
wire  _GEN2241 = io_x[3] ? _GEN2240 : _GEN66;
wire  _GEN2242 = io_x[7] ? _GEN2241 : _GEN65;
wire  _GEN2243 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2244 = io_x[23] ? _GEN2243 : _GEN2242;
wire  _GEN2245 = io_x[2] ? _GEN2244 : _GEN2238;
wire  _GEN2246 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2247 = io_x[11] ? _GEN2246 : _GEN67;
wire  _GEN2248 = io_x[3] ? _GEN2247 : _GEN66;
wire  _GEN2249 = io_x[7] ? _GEN2248 : _GEN65;
wire  _GEN2250 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN2251 = io_x[23] ? _GEN2250 : _GEN2249;
wire  _GEN2252 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2253 = io_x[23] ? _GEN81 : _GEN2252;
wire  _GEN2254 = io_x[2] ? _GEN2253 : _GEN2251;
wire  _GEN2255 = io_x[16] ? _GEN2254 : _GEN2245;
wire  _GEN2256 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2257 = io_x[3] ? _GEN78 : _GEN2256;
wire  _GEN2258 = io_x[7] ? _GEN2257 : _GEN84;
wire  _GEN2259 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2260 = io_x[23] ? _GEN2259 : _GEN2258;
wire  _GEN2261 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2262 = io_x[11] ? _GEN2261 : _GEN67;
wire  _GEN2263 = io_x[3] ? _GEN2262 : _GEN66;
wire  _GEN2264 = io_x[7] ? _GEN65 : _GEN2263;
wire  _GEN2265 = io_x[23] ? _GEN2264 : _GEN74;
wire  _GEN2266 = io_x[2] ? _GEN2265 : _GEN2260;
wire  _GEN2267 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2268 = io_x[11] ? _GEN2267 : _GEN67;
wire  _GEN2269 = io_x[3] ? _GEN2268 : _GEN66;
wire  _GEN2270 = io_x[7] ? _GEN2269 : _GEN84;
wire  _GEN2271 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2272 = io_x[23] ? _GEN2271 : _GEN2270;
wire  _GEN2273 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2274 = io_x[11] ? _GEN2273 : _GEN67;
wire  _GEN2275 = io_x[3] ? _GEN66 : _GEN2274;
wire  _GEN2276 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2277 = io_x[11] ? _GEN2276 : _GEN67;
wire  _GEN2278 = io_x[3] ? _GEN2277 : _GEN78;
wire  _GEN2279 = io_x[7] ? _GEN2278 : _GEN2275;
wire  _GEN2280 = io_x[23] ? _GEN81 : _GEN2279;
wire  _GEN2281 = io_x[2] ? _GEN2280 : _GEN2272;
wire  _GEN2282 = io_x[16] ? _GEN2281 : _GEN2266;
wire  _GEN2283 = io_x[15] ? _GEN2282 : _GEN2255;
wire  _GEN2284 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN2285 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN2286 = io_x[23] ? _GEN2285 : _GEN2284;
wire  _GEN2287 = io_x[2] ? _GEN573 : _GEN2286;
wire  _GEN2288 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2289 = io_x[3] ? _GEN78 : _GEN2288;
wire  _GEN2290 = io_x[7] ? _GEN84 : _GEN2289;
wire  _GEN2291 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2292 = io_x[11] ? _GEN2291 : _GEN67;
wire  _GEN2293 = io_x[3] ? _GEN2292 : _GEN66;
wire  _GEN2294 = io_x[7] ? _GEN2293 : _GEN65;
wire  _GEN2295 = io_x[23] ? _GEN2294 : _GEN2290;
wire  _GEN2296 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2297 = io_x[11] ? _GEN2296 : _GEN67;
wire  _GEN2298 = io_x[3] ? _GEN2297 : _GEN66;
wire  _GEN2299 = io_x[7] ? _GEN2298 : _GEN65;
wire  _GEN2300 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2301 = io_x[7] ? _GEN2300 : _GEN65;
wire  _GEN2302 = io_x[23] ? _GEN2301 : _GEN2299;
wire  _GEN2303 = io_x[2] ? _GEN2302 : _GEN2295;
wire  _GEN2304 = io_x[16] ? _GEN2303 : _GEN2287;
wire  _GEN2305 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2306 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2307 = io_x[3] ? _GEN2306 : _GEN66;
wire  _GEN2308 = io_x[7] ? _GEN2307 : _GEN2305;
wire  _GEN2309 = io_x[23] ? _GEN81 : _GEN2308;
wire  _GEN2310 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2311 = io_x[11] ? _GEN67 : _GEN2310;
wire  _GEN2312 = io_x[3] ? _GEN2311 : _GEN66;
wire  _GEN2313 = io_x[7] ? _GEN2312 : _GEN65;
wire  _GEN2314 = io_x[23] ? _GEN2313 : _GEN74;
wire  _GEN2315 = io_x[2] ? _GEN2314 : _GEN2309;
wire  _GEN2316 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2317 = io_x[11] ? _GEN2316 : _GEN67;
wire  _GEN2318 = io_x[3] ? _GEN2317 : _GEN78;
wire  _GEN2319 = io_x[7] ? _GEN2318 : _GEN65;
wire  _GEN2320 = io_x[23] ? _GEN81 : _GEN2319;
wire  _GEN2321 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2322 = io_x[3] ? _GEN66 : _GEN2321;
wire  _GEN2323 = io_x[7] ? _GEN84 : _GEN2322;
wire  _GEN2324 = io_x[23] ? _GEN81 : _GEN2323;
wire  _GEN2325 = io_x[2] ? _GEN2324 : _GEN2320;
wire  _GEN2326 = io_x[16] ? _GEN2325 : _GEN2315;
wire  _GEN2327 = io_x[15] ? _GEN2326 : _GEN2304;
wire  _GEN2328 = io_x[12] ? _GEN2327 : _GEN2283;
wire  _GEN2329 = io_x[23] ? _GEN81 : _GEN74;
wire  _GEN2330 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2331 = io_x[3] ? _GEN66 : _GEN2330;
wire  _GEN2332 = io_x[7] ? _GEN65 : _GEN2331;
wire  _GEN2333 = io_x[23] ? _GEN2332 : _GEN81;
wire  _GEN2334 = io_x[2] ? _GEN2333 : _GEN2329;
wire  _GEN2335 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2336 = io_x[3] ? _GEN2335 : _GEN66;
wire  _GEN2337 = io_x[7] ? _GEN84 : _GEN2336;
wire  _GEN2338 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2339 = io_x[11] ? _GEN2338 : _GEN67;
wire  _GEN2340 = io_x[3] ? _GEN2339 : _GEN66;
wire  _GEN2341 = io_x[7] ? _GEN65 : _GEN2340;
wire  _GEN2342 = io_x[23] ? _GEN2341 : _GEN2337;
wire  _GEN2343 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2344 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2345 = io_x[11] ? _GEN67 : _GEN2344;
wire  _GEN2346 = io_x[3] ? _GEN2345 : _GEN78;
wire  _GEN2347 = io_x[7] ? _GEN65 : _GEN2346;
wire  _GEN2348 = io_x[23] ? _GEN2347 : _GEN2343;
wire  _GEN2349 = io_x[2] ? _GEN2348 : _GEN2342;
wire  _GEN2350 = io_x[16] ? _GEN2349 : _GEN2334;
wire  _GEN2351 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2352 = io_x[11] ? _GEN67 : _GEN2351;
wire  _GEN2353 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2354 = io_x[11] ? _GEN2353 : _GEN67;
wire  _GEN2355 = io_x[3] ? _GEN2354 : _GEN2352;
wire  _GEN2356 = io_x[7] ? _GEN84 : _GEN2355;
wire  _GEN2357 = io_x[23] ? _GEN74 : _GEN2356;
wire  _GEN2358 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2359 = io_x[11] ? _GEN67 : _GEN2358;
wire  _GEN2360 = io_x[3] ? _GEN66 : _GEN2359;
wire  _GEN2361 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2362 = io_x[11] ? _GEN76 : _GEN2361;
wire  _GEN2363 = io_x[3] ? _GEN2362 : _GEN78;
wire  _GEN2364 = io_x[7] ? _GEN2363 : _GEN2360;
wire  _GEN2365 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2366 = io_x[7] ? _GEN2365 : _GEN65;
wire  _GEN2367 = io_x[23] ? _GEN2366 : _GEN2364;
wire  _GEN2368 = io_x[2] ? _GEN2367 : _GEN2357;
wire  _GEN2369 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2370 = io_x[11] ? _GEN2369 : _GEN67;
wire  _GEN2371 = io_x[3] ? _GEN2370 : _GEN66;
wire  _GEN2372 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2373 = io_x[3] ? _GEN2372 : _GEN66;
wire  _GEN2374 = io_x[7] ? _GEN2373 : _GEN2371;
wire  _GEN2375 = io_x[23] ? _GEN74 : _GEN2374;
wire  _GEN2376 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2377 = io_x[11] ? _GEN2376 : _GEN67;
wire  _GEN2378 = io_x[3] ? _GEN2377 : _GEN66;
wire  _GEN2379 = io_x[7] ? _GEN2378 : _GEN84;
wire  _GEN2380 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2381 = io_x[11] ? _GEN2380 : _GEN67;
wire  _GEN2382 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2383 = io_x[3] ? _GEN2382 : _GEN2381;
wire  _GEN2384 = io_x[7] ? _GEN2383 : _GEN65;
wire  _GEN2385 = io_x[23] ? _GEN2384 : _GEN2379;
wire  _GEN2386 = io_x[2] ? _GEN2385 : _GEN2375;
wire  _GEN2387 = io_x[16] ? _GEN2386 : _GEN2368;
wire  _GEN2388 = io_x[15] ? _GEN2387 : _GEN2350;
wire  _GEN2389 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2390 = io_x[11] ? _GEN2389 : _GEN67;
wire  _GEN2391 = io_x[3] ? _GEN2390 : _GEN66;
wire  _GEN2392 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2393 = io_x[11] ? _GEN2392 : _GEN67;
wire  _GEN2394 = io_x[3] ? _GEN66 : _GEN2393;
wire  _GEN2395 = io_x[7] ? _GEN2394 : _GEN2391;
wire  _GEN2396 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2397 = io_x[23] ? _GEN2396 : _GEN2395;
wire  _GEN2398 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2399 = io_x[11] ? _GEN67 : _GEN2398;
wire  _GEN2400 = io_x[3] ? _GEN2399 : _GEN66;
wire  _GEN2401 = io_x[7] ? _GEN2400 : _GEN84;
wire  _GEN2402 = io_x[23] ? _GEN81 : _GEN2401;
wire  _GEN2403 = io_x[2] ? _GEN2402 : _GEN2397;
wire  _GEN2404 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2405 = io_x[11] ? _GEN67 : _GEN2404;
wire  _GEN2406 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2407 = io_x[11] ? _GEN76 : _GEN2406;
wire  _GEN2408 = io_x[3] ? _GEN2407 : _GEN2405;
wire  _GEN2409 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2410 = io_x[11] ? _GEN67 : _GEN2409;
wire  _GEN2411 = io_x[3] ? _GEN2410 : _GEN66;
wire  _GEN2412 = io_x[7] ? _GEN2411 : _GEN2408;
wire  _GEN2413 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN2414 = io_x[7] ? _GEN65 : _GEN2413;
wire  _GEN2415 = io_x[23] ? _GEN2414 : _GEN2412;
wire  _GEN2416 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2417 = io_x[3] ? _GEN66 : _GEN2416;
wire  _GEN2418 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2419 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2420 = io_x[11] ? _GEN2419 : _GEN67;
wire  _GEN2421 = io_x[3] ? _GEN2420 : _GEN2418;
wire  _GEN2422 = io_x[7] ? _GEN2421 : _GEN2417;
wire  _GEN2423 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2424 = io_x[11] ? _GEN2423 : _GEN67;
wire  _GEN2425 = io_x[3] ? _GEN2424 : _GEN78;
wire  _GEN2426 = io_x[7] ? _GEN2425 : _GEN65;
wire  _GEN2427 = io_x[23] ? _GEN2426 : _GEN2422;
wire  _GEN2428 = io_x[2] ? _GEN2427 : _GEN2415;
wire  _GEN2429 = io_x[16] ? _GEN2428 : _GEN2403;
wire  _GEN2430 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2431 = io_x[11] ? _GEN2430 : _GEN67;
wire  _GEN2432 = io_x[3] ? _GEN66 : _GEN2431;
wire  _GEN2433 = io_x[7] ? _GEN2432 : _GEN65;
wire  _GEN2434 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN2435 = io_x[23] ? _GEN2434 : _GEN2433;
wire  _GEN2436 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2437 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2438 = io_x[11] ? _GEN2437 : _GEN2436;
wire  _GEN2439 = io_x[3] ? _GEN2438 : _GEN66;
wire  _GEN2440 = io_x[7] ? _GEN2439 : _GEN84;
wire  _GEN2441 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2442 = io_x[11] ? _GEN2441 : _GEN67;
wire  _GEN2443 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2444 = io_x[11] ? _GEN2443 : _GEN76;
wire  _GEN2445 = io_x[3] ? _GEN2444 : _GEN2442;
wire  _GEN2446 = io_x[7] ? _GEN2445 : _GEN84;
wire  _GEN2447 = io_x[23] ? _GEN2446 : _GEN2440;
wire  _GEN2448 = io_x[2] ? _GEN2447 : _GEN2435;
wire  _GEN2449 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2450 = io_x[11] ? _GEN67 : _GEN2449;
wire  _GEN2451 = io_x[3] ? _GEN2450 : _GEN78;
wire  _GEN2452 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2453 = io_x[11] ? _GEN76 : _GEN2452;
wire  _GEN2454 = io_x[3] ? _GEN2453 : _GEN66;
wire  _GEN2455 = io_x[7] ? _GEN2454 : _GEN2451;
wire  _GEN2456 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2457 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2458 = io_x[11] ? _GEN2457 : _GEN76;
wire  _GEN2459 = io_x[3] ? _GEN2458 : _GEN78;
wire  _GEN2460 = io_x[7] ? _GEN2459 : _GEN2456;
wire  _GEN2461 = io_x[23] ? _GEN2460 : _GEN2455;
wire  _GEN2462 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2463 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2464 = io_x[11] ? _GEN2463 : _GEN2462;
wire  _GEN2465 = io_x[3] ? _GEN2464 : _GEN66;
wire  _GEN2466 = io_x[7] ? _GEN2465 : _GEN65;
wire  _GEN2467 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2468 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2469 = io_x[3] ? _GEN78 : _GEN2468;
wire  _GEN2470 = io_x[7] ? _GEN2469 : _GEN2467;
wire  _GEN2471 = io_x[23] ? _GEN2470 : _GEN2466;
wire  _GEN2472 = io_x[2] ? _GEN2471 : _GEN2461;
wire  _GEN2473 = io_x[16] ? _GEN2472 : _GEN2448;
wire  _GEN2474 = io_x[15] ? _GEN2473 : _GEN2429;
wire  _GEN2475 = io_x[12] ? _GEN2474 : _GEN2388;
wire  _GEN2476 = io_x[10] ? _GEN2475 : _GEN2328;
wire  _GEN2477 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2478 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2479 = io_x[3] ? _GEN2478 : _GEN66;
wire  _GEN2480 = io_x[7] ? _GEN84 : _GEN2479;
wire  _GEN2481 = io_x[23] ? _GEN2480 : _GEN2477;
wire  _GEN2482 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2483 = io_x[7] ? _GEN65 : _GEN2482;
wire  _GEN2484 = io_x[23] ? _GEN2483 : _GEN81;
wire  _GEN2485 = io_x[2] ? _GEN2484 : _GEN2481;
wire  _GEN2486 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2487 = io_x[3] ? _GEN2486 : _GEN66;
wire  _GEN2488 = io_x[7] ? _GEN2487 : _GEN65;
wire  _GEN2489 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2490 = io_x[11] ? _GEN2489 : _GEN76;
wire  _GEN2491 = io_x[3] ? _GEN2490 : _GEN66;
wire  _GEN2492 = io_x[7] ? _GEN84 : _GEN2491;
wire  _GEN2493 = io_x[23] ? _GEN2492 : _GEN2488;
wire  _GEN2494 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2495 = io_x[3] ? _GEN66 : _GEN2494;
wire  _GEN2496 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2497 = io_x[11] ? _GEN2496 : _GEN76;
wire  _GEN2498 = io_x[3] ? _GEN2497 : _GEN66;
wire  _GEN2499 = io_x[7] ? _GEN2498 : _GEN2495;
wire  _GEN2500 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2501 = io_x[11] ? _GEN2500 : _GEN76;
wire  _GEN2502 = io_x[3] ? _GEN2501 : _GEN78;
wire  _GEN2503 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2504 = io_x[11] ? _GEN2503 : _GEN67;
wire  _GEN2505 = io_x[3] ? _GEN66 : _GEN2504;
wire  _GEN2506 = io_x[7] ? _GEN2505 : _GEN2502;
wire  _GEN2507 = io_x[23] ? _GEN2506 : _GEN2499;
wire  _GEN2508 = io_x[2] ? _GEN2507 : _GEN2493;
wire  _GEN2509 = io_x[16] ? _GEN2508 : _GEN2485;
wire  _GEN2510 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN2511 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2512 = io_x[7] ? _GEN2511 : _GEN65;
wire  _GEN2513 = io_x[23] ? _GEN2512 : _GEN2510;
wire  _GEN2514 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2515 = io_x[3] ? _GEN66 : _GEN2514;
wire  _GEN2516 = io_x[7] ? _GEN84 : _GEN2515;
wire  _GEN2517 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN2518 = io_x[7] ? _GEN84 : _GEN2517;
wire  _GEN2519 = io_x[23] ? _GEN2518 : _GEN2516;
wire  _GEN2520 = io_x[2] ? _GEN2519 : _GEN2513;
wire  _GEN2521 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2522 = io_x[11] ? _GEN2521 : _GEN67;
wire  _GEN2523 = io_x[3] ? _GEN2522 : _GEN66;
wire  _GEN2524 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN2525 = io_x[7] ? _GEN2524 : _GEN2523;
wire  _GEN2526 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2527 = io_x[3] ? _GEN2526 : _GEN66;
wire  _GEN2528 = io_x[7] ? _GEN65 : _GEN2527;
wire  _GEN2529 = io_x[23] ? _GEN2528 : _GEN2525;
wire  _GEN2530 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN2531 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2532 = io_x[11] ? _GEN2531 : _GEN67;
wire  _GEN2533 = io_x[3] ? _GEN2532 : _GEN78;
wire  _GEN2534 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2535 = io_x[11] ? _GEN2534 : _GEN67;
wire  _GEN2536 = io_x[3] ? _GEN2535 : _GEN78;
wire  _GEN2537 = io_x[7] ? _GEN2536 : _GEN2533;
wire  _GEN2538 = io_x[23] ? _GEN2537 : _GEN2530;
wire  _GEN2539 = io_x[2] ? _GEN2538 : _GEN2529;
wire  _GEN2540 = io_x[16] ? _GEN2539 : _GEN2520;
wire  _GEN2541 = io_x[15] ? _GEN2540 : _GEN2509;
wire  _GEN2542 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2543 = io_x[7] ? _GEN2542 : _GEN65;
wire  _GEN2544 = io_x[23] ? _GEN74 : _GEN2543;
wire  _GEN2545 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2546 = io_x[11] ? _GEN2545 : _GEN67;
wire  _GEN2547 = io_x[3] ? _GEN2546 : _GEN66;
wire  _GEN2548 = io_x[7] ? _GEN2547 : _GEN84;
wire  _GEN2549 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2550 = io_x[7] ? _GEN2549 : _GEN84;
wire  _GEN2551 = io_x[23] ? _GEN2550 : _GEN2548;
wire  _GEN2552 = io_x[2] ? _GEN2551 : _GEN2544;
wire  _GEN2553 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2554 = io_x[11] ? _GEN2553 : _GEN76;
wire  _GEN2555 = io_x[3] ? _GEN2554 : _GEN66;
wire  _GEN2556 = io_x[7] ? _GEN2555 : _GEN65;
wire  _GEN2557 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN2558 = io_x[23] ? _GEN2557 : _GEN2556;
wire  _GEN2559 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2560 = io_x[11] ? _GEN2559 : _GEN67;
wire  _GEN2561 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2562 = io_x[11] ? _GEN2561 : _GEN67;
wire  _GEN2563 = io_x[3] ? _GEN2562 : _GEN2560;
wire  _GEN2564 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2565 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2566 = io_x[11] ? _GEN2565 : _GEN2564;
wire  _GEN2567 = io_x[3] ? _GEN2566 : _GEN66;
wire  _GEN2568 = io_x[7] ? _GEN2567 : _GEN2563;
wire  _GEN2569 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2570 = io_x[11] ? _GEN2569 : _GEN67;
wire  _GEN2571 = io_x[3] ? _GEN2570 : _GEN66;
wire  _GEN2572 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2573 = io_x[11] ? _GEN67 : _GEN2572;
wire  _GEN2574 = io_x[3] ? _GEN2573 : _GEN66;
wire  _GEN2575 = io_x[7] ? _GEN2574 : _GEN2571;
wire  _GEN2576 = io_x[23] ? _GEN2575 : _GEN2568;
wire  _GEN2577 = io_x[2] ? _GEN2576 : _GEN2558;
wire  _GEN2578 = io_x[16] ? _GEN2577 : _GEN2552;
wire  _GEN2579 = io_x[23] ? _GEN81 : _GEN74;
wire  _GEN2580 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2581 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2582 = io_x[11] ? _GEN2581 : _GEN2580;
wire  _GEN2583 = io_x[3] ? _GEN2582 : _GEN66;
wire  _GEN2584 = io_x[7] ? _GEN2583 : _GEN2515;
wire  _GEN2585 = io_x[23] ? _GEN74 : _GEN2584;
wire  _GEN2586 = io_x[2] ? _GEN2585 : _GEN2579;
wire  _GEN2587 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2588 = io_x[3] ? _GEN2587 : _GEN78;
wire  _GEN2589 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2590 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2591 = io_x[11] ? _GEN2590 : _GEN67;
wire  _GEN2592 = io_x[3] ? _GEN2591 : _GEN2589;
wire  _GEN2593 = io_x[7] ? _GEN2592 : _GEN2588;
wire  _GEN2594 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2595 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2596 = io_x[11] ? _GEN2595 : _GEN2594;
wire  _GEN2597 = io_x[3] ? _GEN2596 : _GEN66;
wire  _GEN2598 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2599 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2600 = io_x[11] ? _GEN2599 : _GEN2598;
wire  _GEN2601 = io_x[3] ? _GEN2600 : _GEN66;
wire  _GEN2602 = io_x[7] ? _GEN2601 : _GEN2597;
wire  _GEN2603 = io_x[23] ? _GEN2602 : _GEN2593;
wire  _GEN2604 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2605 = io_x[11] ? _GEN2604 : _GEN67;
wire  _GEN2606 = io_x[3] ? _GEN2605 : _GEN66;
wire  _GEN2607 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2608 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2609 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2610 = io_x[11] ? _GEN2609 : _GEN2608;
wire  _GEN2611 = io_x[3] ? _GEN2610 : _GEN2607;
wire  _GEN2612 = io_x[7] ? _GEN2611 : _GEN2606;
wire  _GEN2613 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2614 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2615 = io_x[11] ? _GEN2614 : _GEN2613;
wire  _GEN2616 = io_x[3] ? _GEN2615 : _GEN66;
wire  _GEN2617 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2618 = io_x[11] ? _GEN2617 : _GEN76;
wire  _GEN2619 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2620 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2621 = io_x[11] ? _GEN2620 : _GEN2619;
wire  _GEN2622 = io_x[3] ? _GEN2621 : _GEN2618;
wire  _GEN2623 = io_x[7] ? _GEN2622 : _GEN2616;
wire  _GEN2624 = io_x[23] ? _GEN2623 : _GEN2612;
wire  _GEN2625 = io_x[2] ? _GEN2624 : _GEN2603;
wire  _GEN2626 = io_x[16] ? _GEN2625 : _GEN2586;
wire  _GEN2627 = io_x[15] ? _GEN2626 : _GEN2578;
wire  _GEN2628 = io_x[12] ? _GEN2627 : _GEN2541;
wire  _GEN2629 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN2630 = io_x[23] ? _GEN81 : _GEN2629;
wire  _GEN2631 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2632 = io_x[3] ? _GEN2631 : _GEN66;
wire  _GEN2633 = io_x[7] ? _GEN2632 : _GEN65;
wire  _GEN2634 = io_x[23] ? _GEN74 : _GEN2633;
wire  _GEN2635 = io_x[2] ? _GEN2634 : _GEN2630;
wire  _GEN2636 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2637 = io_x[3] ? _GEN2636 : _GEN66;
wire  _GEN2638 = io_x[7] ? _GEN2637 : _GEN65;
wire  _GEN2639 = io_x[23] ? _GEN81 : _GEN2638;
wire  _GEN2640 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2641 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2642 = io_x[11] ? _GEN2641 : _GEN2640;
wire  _GEN2643 = io_x[3] ? _GEN2642 : _GEN66;
wire  _GEN2644 = io_x[7] ? _GEN2643 : _GEN84;
wire  _GEN2645 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2646 = io_x[11] ? _GEN2645 : _GEN76;
wire  _GEN2647 = io_x[3] ? _GEN2646 : _GEN66;
wire  _GEN2648 = io_x[7] ? _GEN2647 : _GEN84;
wire  _GEN2649 = io_x[23] ? _GEN2648 : _GEN2644;
wire  _GEN2650 = io_x[2] ? _GEN2649 : _GEN2639;
wire  _GEN2651 = io_x[16] ? _GEN2650 : _GEN2635;
wire  _GEN2652 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2653 = io_x[11] ? _GEN2652 : _GEN67;
wire  _GEN2654 = io_x[3] ? _GEN78 : _GEN2653;
wire  _GEN2655 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2656 = io_x[3] ? _GEN2655 : _GEN66;
wire  _GEN2657 = io_x[7] ? _GEN2656 : _GEN2654;
wire  _GEN2658 = io_x[23] ? _GEN74 : _GEN2657;
wire  _GEN2659 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN2660 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2661 = io_x[11] ? _GEN2660 : _GEN67;
wire  _GEN2662 = io_x[3] ? _GEN2661 : _GEN66;
wire  _GEN2663 = io_x[7] ? _GEN2662 : _GEN2659;
wire  _GEN2664 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2665 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2666 = io_x[3] ? _GEN2665 : _GEN2664;
wire  _GEN2667 = io_x[7] ? _GEN2666 : _GEN84;
wire  _GEN2668 = io_x[23] ? _GEN2667 : _GEN2663;
wire  _GEN2669 = io_x[2] ? _GEN2668 : _GEN2658;
wire  _GEN2670 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2671 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2672 = io_x[11] ? _GEN2671 : _GEN2670;
wire  _GEN2673 = io_x[3] ? _GEN2672 : _GEN66;
wire  _GEN2674 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2675 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2676 = io_x[11] ? _GEN2675 : _GEN67;
wire  _GEN2677 = io_x[3] ? _GEN2676 : _GEN2674;
wire  _GEN2678 = io_x[7] ? _GEN2677 : _GEN2673;
wire  _GEN2679 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2680 = io_x[11] ? _GEN2679 : _GEN76;
wire  _GEN2681 = io_x[3] ? _GEN2680 : _GEN66;
wire  _GEN2682 = io_x[7] ? _GEN65 : _GEN2681;
wire  _GEN2683 = io_x[23] ? _GEN2682 : _GEN2678;
wire  _GEN2684 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2685 = io_x[11] ? _GEN2684 : _GEN67;
wire  _GEN2686 = io_x[3] ? _GEN2685 : _GEN66;
wire  _GEN2687 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2688 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2689 = io_x[11] ? _GEN2688 : _GEN2687;
wire  _GEN2690 = io_x[3] ? _GEN2689 : _GEN66;
wire  _GEN2691 = io_x[7] ? _GEN2690 : _GEN2686;
wire  _GEN2692 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2693 = io_x[11] ? _GEN2692 : _GEN76;
wire  _GEN2694 = io_x[3] ? _GEN66 : _GEN2693;
wire  _GEN2695 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2696 = io_x[11] ? _GEN2695 : _GEN67;
wire  _GEN2697 = io_x[3] ? _GEN2696 : _GEN66;
wire  _GEN2698 = io_x[7] ? _GEN2697 : _GEN2694;
wire  _GEN2699 = io_x[23] ? _GEN2698 : _GEN2691;
wire  _GEN2700 = io_x[2] ? _GEN2699 : _GEN2683;
wire  _GEN2701 = io_x[16] ? _GEN2700 : _GEN2669;
wire  _GEN2702 = io_x[15] ? _GEN2701 : _GEN2651;
wire  _GEN2703 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2704 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2705 = io_x[3] ? _GEN66 : _GEN2704;
wire  _GEN2706 = io_x[7] ? _GEN2705 : _GEN2703;
wire  _GEN2707 = io_x[23] ? _GEN74 : _GEN2706;
wire  _GEN2708 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2709 = io_x[11] ? _GEN76 : _GEN2708;
wire  _GEN2710 = io_x[3] ? _GEN78 : _GEN2709;
wire  _GEN2711 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2712 = io_x[11] ? _GEN2711 : _GEN76;
wire  _GEN2713 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2714 = io_x[3] ? _GEN2713 : _GEN2712;
wire  _GEN2715 = io_x[7] ? _GEN2714 : _GEN2710;
wire  _GEN2716 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2717 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2718 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2719 = io_x[11] ? _GEN2718 : _GEN2717;
wire  _GEN2720 = io_x[3] ? _GEN2719 : _GEN2716;
wire  _GEN2721 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2722 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2723 = io_x[11] ? _GEN2722 : _GEN2721;
wire  _GEN2724 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2725 = io_x[11] ? _GEN67 : _GEN2724;
wire  _GEN2726 = io_x[3] ? _GEN2725 : _GEN2723;
wire  _GEN2727 = io_x[7] ? _GEN2726 : _GEN2720;
wire  _GEN2728 = io_x[23] ? _GEN2727 : _GEN2715;
wire  _GEN2729 = io_x[2] ? _GEN2728 : _GEN2707;
wire  _GEN2730 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2731 = io_x[11] ? _GEN67 : _GEN2730;
wire  _GEN2732 = io_x[3] ? _GEN2731 : _GEN78;
wire  _GEN2733 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2734 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2735 = io_x[11] ? _GEN2734 : _GEN2733;
wire  _GEN2736 = io_x[3] ? _GEN2735 : _GEN66;
wire  _GEN2737 = io_x[7] ? _GEN2736 : _GEN2732;
wire  _GEN2738 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2739 = io_x[11] ? _GEN67 : _GEN2738;
wire  _GEN2740 = io_x[3] ? _GEN2739 : _GEN78;
wire  _GEN2741 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2742 = io_x[7] ? _GEN2741 : _GEN2740;
wire  _GEN2743 = io_x[23] ? _GEN2742 : _GEN2737;
wire  _GEN2744 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2745 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2746 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2747 = io_x[11] ? _GEN2746 : _GEN2745;
wire  _GEN2748 = io_x[3] ? _GEN2747 : _GEN2744;
wire  _GEN2749 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2750 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2751 = io_x[11] ? _GEN2750 : _GEN2749;
wire  _GEN2752 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2753 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2754 = io_x[11] ? _GEN2753 : _GEN2752;
wire  _GEN2755 = io_x[3] ? _GEN2754 : _GEN2751;
wire  _GEN2756 = io_x[7] ? _GEN2755 : _GEN2748;
wire  _GEN2757 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2758 = io_x[11] ? _GEN67 : _GEN2757;
wire  _GEN2759 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2760 = io_x[11] ? _GEN2759 : _GEN76;
wire  _GEN2761 = io_x[3] ? _GEN2760 : _GEN2758;
wire  _GEN2762 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2763 = io_x[11] ? _GEN76 : _GEN2762;
wire  _GEN2764 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2765 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2766 = io_x[11] ? _GEN2765 : _GEN2764;
wire  _GEN2767 = io_x[3] ? _GEN2766 : _GEN2763;
wire  _GEN2768 = io_x[7] ? _GEN2767 : _GEN2761;
wire  _GEN2769 = io_x[23] ? _GEN2768 : _GEN2756;
wire  _GEN2770 = io_x[2] ? _GEN2769 : _GEN2743;
wire  _GEN2771 = io_x[16] ? _GEN2770 : _GEN2729;
wire  _GEN2772 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN2773 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2774 = io_x[11] ? _GEN2773 : _GEN76;
wire  _GEN2775 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2776 = io_x[11] ? _GEN2775 : _GEN67;
wire  _GEN2777 = io_x[3] ? _GEN2776 : _GEN2774;
wire  _GEN2778 = io_x[7] ? _GEN2777 : _GEN2772;
wire  _GEN2779 = io_x[23] ? _GEN74 : _GEN2778;
wire  _GEN2780 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2781 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2782 = io_x[11] ? _GEN2781 : _GEN67;
wire  _GEN2783 = io_x[3] ? _GEN2782 : _GEN66;
wire  _GEN2784 = io_x[7] ? _GEN2783 : _GEN2780;
wire  _GEN2785 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2786 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2787 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2788 = io_x[11] ? _GEN2787 : _GEN2786;
wire  _GEN2789 = io_x[3] ? _GEN2788 : _GEN2785;
wire  _GEN2790 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2791 = io_x[11] ? _GEN76 : _GEN2790;
wire  _GEN2792 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2793 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2794 = io_x[11] ? _GEN2793 : _GEN2792;
wire  _GEN2795 = io_x[3] ? _GEN2794 : _GEN2791;
wire  _GEN2796 = io_x[7] ? _GEN2795 : _GEN2789;
wire  _GEN2797 = io_x[23] ? _GEN2796 : _GEN2784;
wire  _GEN2798 = io_x[2] ? _GEN2797 : _GEN2779;
wire  _GEN2799 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2800 = io_x[11] ? _GEN2799 : _GEN67;
wire  _GEN2801 = io_x[3] ? _GEN2800 : _GEN66;
wire  _GEN2802 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2803 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2804 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2805 = io_x[11] ? _GEN2804 : _GEN2803;
wire  _GEN2806 = io_x[3] ? _GEN2805 : _GEN2802;
wire  _GEN2807 = io_x[7] ? _GEN2806 : _GEN2801;
wire  _GEN2808 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2809 = io_x[3] ? _GEN2808 : _GEN66;
wire  _GEN2810 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2811 = io_x[11] ? _GEN2810 : _GEN67;
wire  _GEN2812 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2813 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2814 = io_x[11] ? _GEN2813 : _GEN2812;
wire  _GEN2815 = io_x[3] ? _GEN2814 : _GEN2811;
wire  _GEN2816 = io_x[7] ? _GEN2815 : _GEN2809;
wire  _GEN2817 = io_x[23] ? _GEN2816 : _GEN2807;
wire  _GEN2818 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2819 = io_x[3] ? _GEN66 : _GEN2818;
wire  _GEN2820 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2821 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2822 = io_x[11] ? _GEN2821 : _GEN2820;
wire  _GEN2823 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2824 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2825 = io_x[11] ? _GEN2824 : _GEN2823;
wire  _GEN2826 = io_x[3] ? _GEN2825 : _GEN2822;
wire  _GEN2827 = io_x[7] ? _GEN2826 : _GEN2819;
wire  _GEN2828 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2829 = io_x[11] ? _GEN76 : _GEN2828;
wire  _GEN2830 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2831 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2832 = io_x[11] ? _GEN2831 : _GEN2830;
wire  _GEN2833 = io_x[3] ? _GEN2832 : _GEN2829;
wire  _GEN2834 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2835 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2836 = io_x[11] ? _GEN2835 : _GEN2834;
wire  _GEN2837 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2838 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2839 = io_x[11] ? _GEN2838 : _GEN2837;
wire  _GEN2840 = io_x[3] ? _GEN2839 : _GEN2836;
wire  _GEN2841 = io_x[7] ? _GEN2840 : _GEN2833;
wire  _GEN2842 = io_x[23] ? _GEN2841 : _GEN2827;
wire  _GEN2843 = io_x[2] ? _GEN2842 : _GEN2817;
wire  _GEN2844 = io_x[16] ? _GEN2843 : _GEN2798;
wire  _GEN2845 = io_x[15] ? _GEN2844 : _GEN2771;
wire  _GEN2846 = io_x[12] ? _GEN2845 : _GEN2702;
wire  _GEN2847 = io_x[10] ? _GEN2846 : _GEN2628;
wire  _GEN2848 = io_x[4] ? _GEN2847 : _GEN2476;
wire  _GEN2849 = io_x[8] ? _GEN2848 : _GEN2237;
wire  _GEN2850 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN2851 = io_x[2] ? _GEN140 : _GEN2850;
wire  _GEN2852 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2853 = io_x[11] ? _GEN2852 : _GEN67;
wire  _GEN2854 = io_x[3] ? _GEN2853 : _GEN66;
wire  _GEN2855 = io_x[7] ? _GEN2854 : _GEN65;
wire  _GEN2856 = io_x[23] ? _GEN74 : _GEN2855;
wire  _GEN2857 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2858 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2859 = io_x[11] ? _GEN2858 : _GEN67;
wire  _GEN2860 = io_x[3] ? _GEN2859 : _GEN2857;
wire  _GEN2861 = io_x[7] ? _GEN2860 : _GEN65;
wire  _GEN2862 = io_x[23] ? _GEN74 : _GEN2861;
wire  _GEN2863 = io_x[2] ? _GEN2862 : _GEN2856;
wire  _GEN2864 = io_x[16] ? _GEN2863 : _GEN2851;
wire  _GEN2865 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2866 = io_x[23] ? _GEN2865 : _GEN81;
wire  _GEN2867 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2868 = io_x[11] ? _GEN2867 : _GEN67;
wire  _GEN2869 = io_x[3] ? _GEN2868 : _GEN66;
wire  _GEN2870 = io_x[7] ? _GEN2869 : _GEN65;
wire  _GEN2871 = io_x[23] ? _GEN2870 : _GEN74;
wire  _GEN2872 = io_x[2] ? _GEN2871 : _GEN2866;
wire  _GEN2873 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2874 = io_x[11] ? _GEN2873 : _GEN67;
wire  _GEN2875 = io_x[3] ? _GEN2874 : _GEN66;
wire  _GEN2876 = io_x[7] ? _GEN2875 : _GEN65;
wire  _GEN2877 = io_x[23] ? _GEN81 : _GEN2876;
wire  _GEN2878 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2879 = io_x[11] ? _GEN2878 : _GEN67;
wire  _GEN2880 = io_x[3] ? _GEN2879 : _GEN66;
wire  _GEN2881 = io_x[7] ? _GEN2880 : _GEN65;
wire  _GEN2882 = io_x[23] ? _GEN81 : _GEN2881;
wire  _GEN2883 = io_x[2] ? _GEN2882 : _GEN2877;
wire  _GEN2884 = io_x[16] ? _GEN2883 : _GEN2872;
wire  _GEN2885 = io_x[15] ? _GEN2884 : _GEN2864;
wire  _GEN2886 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN2887 = io_x[23] ? _GEN2886 : _GEN81;
wire  _GEN2888 = io_x[2] ? _GEN573 : _GEN2887;
wire  _GEN2889 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2890 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2891 = io_x[11] ? _GEN2890 : _GEN67;
wire  _GEN2892 = io_x[3] ? _GEN2891 : _GEN66;
wire  _GEN2893 = io_x[7] ? _GEN2892 : _GEN2889;
wire  _GEN2894 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2895 = io_x[11] ? _GEN67 : _GEN2894;
wire  _GEN2896 = io_x[3] ? _GEN2895 : _GEN66;
wire  _GEN2897 = io_x[7] ? _GEN65 : _GEN2896;
wire  _GEN2898 = io_x[23] ? _GEN2897 : _GEN2893;
wire  _GEN2899 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN2900 = io_x[11] ? _GEN2899 : _GEN67;
wire  _GEN2901 = io_x[3] ? _GEN2900 : _GEN78;
wire  _GEN2902 = io_x[7] ? _GEN2901 : _GEN65;
wire  _GEN2903 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN2904 = io_x[23] ? _GEN2903 : _GEN2902;
wire  _GEN2905 = io_x[2] ? _GEN2904 : _GEN2898;
wire  _GEN2906 = io_x[16] ? _GEN2905 : _GEN2888;
wire  _GEN2907 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2908 = io_x[3] ? _GEN78 : _GEN2907;
wire  _GEN2909 = io_x[7] ? _GEN2908 : _GEN65;
wire  _GEN2910 = io_x[23] ? _GEN74 : _GEN2909;
wire  _GEN2911 = io_x[2] ? _GEN2910 : _GEN140;
wire  _GEN2912 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN2913 = io_x[7] ? _GEN2912 : _GEN65;
wire  _GEN2914 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2915 = io_x[23] ? _GEN2914 : _GEN2913;
wire  _GEN2916 = io_x[2] ? _GEN2915 : _GEN140;
wire  _GEN2917 = io_x[16] ? _GEN2916 : _GEN2911;
wire  _GEN2918 = io_x[15] ? _GEN2917 : _GEN2906;
wire  _GEN2919 = io_x[12] ? _GEN2918 : _GEN2885;
wire  _GEN2920 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2921 = io_x[11] ? _GEN2920 : _GEN67;
wire  _GEN2922 = io_x[3] ? _GEN2921 : _GEN66;
wire  _GEN2923 = io_x[7] ? _GEN65 : _GEN2922;
wire  _GEN2924 = io_x[23] ? _GEN2923 : _GEN74;
wire  _GEN2925 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2926 = io_x[7] ? _GEN2925 : _GEN84;
wire  _GEN2927 = io_x[23] ? _GEN81 : _GEN2926;
wire  _GEN2928 = io_x[2] ? _GEN2927 : _GEN2924;
wire  _GEN2929 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN2930 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2931 = io_x[3] ? _GEN2930 : _GEN66;
wire  _GEN2932 = io_x[7] ? _GEN2931 : _GEN2929;
wire  _GEN2933 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2934 = io_x[11] ? _GEN67 : _GEN2933;
wire  _GEN2935 = io_x[3] ? _GEN2934 : _GEN66;
wire  _GEN2936 = io_x[7] ? _GEN2935 : _GEN84;
wire  _GEN2937 = io_x[23] ? _GEN2936 : _GEN2932;
wire  _GEN2938 = io_x[2] ? _GEN140 : _GEN2937;
wire  _GEN2939 = io_x[16] ? _GEN2938 : _GEN2928;
wire  _GEN2940 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2941 = io_x[3] ? _GEN2940 : _GEN78;
wire  _GEN2942 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2943 = io_x[3] ? _GEN66 : _GEN2942;
wire  _GEN2944 = io_x[7] ? _GEN2943 : _GEN2941;
wire  _GEN2945 = io_x[23] ? _GEN74 : _GEN2944;
wire  _GEN2946 = io_x[2] ? _GEN2945 : _GEN573;
wire  _GEN2947 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2948 = io_x[3] ? _GEN66 : _GEN2947;
wire  _GEN2949 = io_x[7] ? _GEN84 : _GEN2948;
wire  _GEN2950 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2951 = io_x[3] ? _GEN2950 : _GEN66;
wire  _GEN2952 = io_x[7] ? _GEN2951 : _GEN65;
wire  _GEN2953 = io_x[23] ? _GEN2952 : _GEN2949;
wire  _GEN2954 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2955 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2956 = io_x[11] ? _GEN2955 : _GEN67;
wire  _GEN2957 = io_x[3] ? _GEN2956 : _GEN2954;
wire  _GEN2958 = io_x[7] ? _GEN2957 : _GEN65;
wire  _GEN2959 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2960 = io_x[3] ? _GEN2959 : _GEN66;
wire  _GEN2961 = io_x[7] ? _GEN2960 : _GEN65;
wire  _GEN2962 = io_x[23] ? _GEN2961 : _GEN2958;
wire  _GEN2963 = io_x[2] ? _GEN2962 : _GEN2953;
wire  _GEN2964 = io_x[16] ? _GEN2963 : _GEN2946;
wire  _GEN2965 = io_x[15] ? _GEN2964 : _GEN2939;
wire  _GEN2966 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2967 = io_x[11] ? _GEN67 : _GEN2966;
wire  _GEN2968 = io_x[3] ? _GEN2967 : _GEN66;
wire  _GEN2969 = io_x[7] ? _GEN2968 : _GEN84;
wire  _GEN2970 = io_x[23] ? _GEN74 : _GEN2969;
wire  _GEN2971 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2972 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN2973 = io_x[11] ? _GEN67 : _GEN2972;
wire  _GEN2974 = io_x[3] ? _GEN2973 : _GEN2971;
wire  _GEN2975 = io_x[7] ? _GEN2974 : _GEN65;
wire  _GEN2976 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2977 = io_x[23] ? _GEN2976 : _GEN2975;
wire  _GEN2978 = io_x[2] ? _GEN2977 : _GEN2970;
wire  _GEN2979 = io_x[16] ? _GEN2978 : _GEN1332;
wire  _GEN2980 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2981 = io_x[7] ? _GEN65 : _GEN2980;
wire  _GEN2982 = io_x[23] ? _GEN81 : _GEN2981;
wire  _GEN2983 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2984 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN2985 = io_x[23] ? _GEN2984 : _GEN2983;
wire  _GEN2986 = io_x[2] ? _GEN2985 : _GEN2982;
wire  _GEN2987 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN2988 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2989 = io_x[3] ? _GEN2988 : _GEN66;
wire  _GEN2990 = io_x[7] ? _GEN2989 : _GEN2987;
wire  _GEN2991 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN2992 = io_x[3] ? _GEN2991 : _GEN66;
wire  _GEN2993 = io_x[7] ? _GEN2992 : _GEN65;
wire  _GEN2994 = io_x[23] ? _GEN2993 : _GEN2990;
wire  _GEN2995 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN2996 = io_x[3] ? _GEN66 : _GEN2995;
wire  _GEN2997 = io_x[7] ? _GEN2996 : _GEN65;
wire  _GEN2998 = io_x[23] ? _GEN74 : _GEN2997;
wire  _GEN2999 = io_x[2] ? _GEN2998 : _GEN2994;
wire  _GEN3000 = io_x[16] ? _GEN2999 : _GEN2986;
wire  _GEN3001 = io_x[15] ? _GEN3000 : _GEN2979;
wire  _GEN3002 = io_x[12] ? _GEN3001 : _GEN2965;
wire  _GEN3003 = io_x[10] ? _GEN3002 : _GEN2919;
wire  _GEN3004 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN3005 = io_x[23] ? _GEN81 : _GEN3004;
wire  _GEN3006 = io_x[2] ? _GEN573 : _GEN3005;
wire  _GEN3007 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN3008 = io_x[23] ? _GEN81 : _GEN3007;
wire  _GEN3009 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3010 = io_x[11] ? _GEN3009 : _GEN67;
wire  _GEN3011 = io_x[3] ? _GEN3010 : _GEN66;
wire  _GEN3012 = io_x[7] ? _GEN3011 : _GEN65;
wire  _GEN3013 = io_x[23] ? _GEN3012 : _GEN81;
wire  _GEN3014 = io_x[2] ? _GEN3013 : _GEN3008;
wire  _GEN3015 = io_x[16] ? _GEN3014 : _GEN3006;
wire  _GEN3016 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3017 = io_x[7] ? _GEN3016 : _GEN65;
wire  _GEN3018 = io_x[23] ? _GEN3017 : _GEN74;
wire  _GEN3019 = io_x[2] ? _GEN3018 : _GEN140;
wire  _GEN3020 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3021 = io_x[11] ? _GEN3020 : _GEN67;
wire  _GEN3022 = io_x[3] ? _GEN3021 : _GEN66;
wire  _GEN3023 = io_x[7] ? _GEN3022 : _GEN65;
wire  _GEN3024 = io_x[23] ? _GEN81 : _GEN3023;
wire  _GEN3025 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN3026 = io_x[2] ? _GEN3025 : _GEN3024;
wire  _GEN3027 = io_x[16] ? _GEN3026 : _GEN3019;
wire  _GEN3028 = io_x[15] ? _GEN3027 : _GEN3015;
wire  _GEN3029 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN3030 = io_x[23] ? _GEN3029 : _GEN81;
wire  _GEN3031 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3032 = io_x[3] ? _GEN66 : _GEN3031;
wire  _GEN3033 = io_x[7] ? _GEN3032 : _GEN84;
wire  _GEN3034 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN3035 = io_x[23] ? _GEN3034 : _GEN3033;
wire  _GEN3036 = io_x[2] ? _GEN3035 : _GEN3030;
wire  _GEN3037 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3038 = io_x[3] ? _GEN3037 : _GEN66;
wire  _GEN3039 = io_x[7] ? _GEN3038 : _GEN65;
wire  _GEN3040 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3041 = io_x[7] ? _GEN3040 : _GEN65;
wire  _GEN3042 = io_x[23] ? _GEN3041 : _GEN3039;
wire  _GEN3043 = io_x[2] ? _GEN3042 : _GEN573;
wire  _GEN3044 = io_x[16] ? _GEN3043 : _GEN3036;
wire  _GEN3045 = io_x[23] ? _GEN74 : _GEN81;
wire  _GEN3046 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3047 = io_x[3] ? _GEN3046 : _GEN78;
wire  _GEN3048 = io_x[7] ? _GEN3047 : _GEN65;
wire  _GEN3049 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN3050 = io_x[23] ? _GEN3049 : _GEN3048;
wire  _GEN3051 = io_x[2] ? _GEN3050 : _GEN3045;
wire  _GEN3052 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3053 = io_x[11] ? _GEN3052 : _GEN76;
wire  _GEN3054 = io_x[3] ? _GEN3053 : _GEN66;
wire  _GEN3055 = io_x[7] ? _GEN3054 : _GEN84;
wire  _GEN3056 = io_x[23] ? _GEN74 : _GEN3055;
wire  _GEN3057 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3058 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3059 = io_x[11] ? _GEN3058 : _GEN3057;
wire  _GEN3060 = io_x[3] ? _GEN3059 : _GEN78;
wire  _GEN3061 = io_x[7] ? _GEN3060 : _GEN65;
wire  _GEN3062 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3063 = io_x[3] ? _GEN3062 : _GEN78;
wire  _GEN3064 = io_x[7] ? _GEN3063 : _GEN65;
wire  _GEN3065 = io_x[23] ? _GEN3064 : _GEN3061;
wire  _GEN3066 = io_x[2] ? _GEN3065 : _GEN3056;
wire  _GEN3067 = io_x[16] ? _GEN3066 : _GEN3051;
wire  _GEN3068 = io_x[15] ? _GEN3067 : _GEN3044;
wire  _GEN3069 = io_x[12] ? _GEN3068 : _GEN3028;
wire  _GEN3070 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3071 = io_x[3] ? _GEN66 : _GEN3070;
wire  _GEN3072 = io_x[7] ? _GEN3071 : _GEN65;
wire  _GEN3073 = io_x[23] ? _GEN81 : _GEN3072;
wire  _GEN3074 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3075 = io_x[11] ? _GEN76 : _GEN3074;
wire  _GEN3076 = io_x[3] ? _GEN78 : _GEN3075;
wire  _GEN3077 = io_x[7] ? _GEN3076 : _GEN65;
wire  _GEN3078 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3079 = io_x[3] ? _GEN66 : _GEN3078;
wire  _GEN3080 = io_x[7] ? _GEN3079 : _GEN65;
wire  _GEN3081 = io_x[23] ? _GEN3080 : _GEN3077;
wire  _GEN3082 = io_x[2] ? _GEN3081 : _GEN3073;
wire  _GEN3083 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN3084 = io_x[23] ? _GEN3083 : _GEN74;
wire  _GEN3085 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3086 = io_x[3] ? _GEN3085 : _GEN66;
wire  _GEN3087 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3088 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3089 = io_x[3] ? _GEN3088 : _GEN3087;
wire  _GEN3090 = io_x[7] ? _GEN3089 : _GEN3086;
wire  _GEN3091 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3092 = io_x[3] ? _GEN78 : _GEN3091;
wire  _GEN3093 = io_x[7] ? _GEN3092 : _GEN65;
wire  _GEN3094 = io_x[23] ? _GEN3093 : _GEN3090;
wire  _GEN3095 = io_x[2] ? _GEN3094 : _GEN3084;
wire  _GEN3096 = io_x[16] ? _GEN3095 : _GEN3082;
wire  _GEN3097 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN3098 = io_x[23] ? _GEN3097 : _GEN81;
wire  _GEN3099 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3100 = io_x[3] ? _GEN66 : _GEN3099;
wire  _GEN3101 = io_x[7] ? _GEN3100 : _GEN84;
wire  _GEN3102 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3103 = io_x[3] ? _GEN66 : _GEN3102;
wire  _GEN3104 = io_x[7] ? _GEN3103 : _GEN65;
wire  _GEN3105 = io_x[23] ? _GEN3104 : _GEN3101;
wire  _GEN3106 = io_x[2] ? _GEN3105 : _GEN3098;
wire  _GEN3107 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3108 = io_x[7] ? _GEN3107 : _GEN65;
wire  _GEN3109 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN3110 = io_x[23] ? _GEN3109 : _GEN3108;
wire  _GEN3111 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3112 = io_x[3] ? _GEN3111 : _GEN66;
wire  _GEN3113 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3114 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3115 = io_x[11] ? _GEN3114 : _GEN67;
wire  _GEN3116 = io_x[3] ? _GEN3115 : _GEN3113;
wire  _GEN3117 = io_x[7] ? _GEN3116 : _GEN3112;
wire  _GEN3118 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3119 = io_x[11] ? _GEN3118 : _GEN76;
wire  _GEN3120 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3121 = io_x[3] ? _GEN3120 : _GEN3119;
wire  _GEN3122 = io_x[7] ? _GEN3121 : _GEN65;
wire  _GEN3123 = io_x[23] ? _GEN3122 : _GEN3117;
wire  _GEN3124 = io_x[2] ? _GEN3123 : _GEN3110;
wire  _GEN3125 = io_x[16] ? _GEN3124 : _GEN3106;
wire  _GEN3126 = io_x[15] ? _GEN3125 : _GEN3096;
wire  _GEN3127 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3128 = io_x[11] ? _GEN67 : _GEN3127;
wire  _GEN3129 = io_x[3] ? _GEN66 : _GEN3128;
wire  _GEN3130 = io_x[7] ? _GEN84 : _GEN3129;
wire  _GEN3131 = io_x[23] ? _GEN74 : _GEN3130;
wire  _GEN3132 = io_x[2] ? _GEN3131 : _GEN140;
wire  _GEN3133 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3134 = io_x[3] ? _GEN3133 : _GEN66;
wire  _GEN3135 = io_x[7] ? _GEN84 : _GEN3134;
wire  _GEN3136 = io_x[23] ? _GEN3135 : _GEN74;
wire  _GEN3137 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3138 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3139 = io_x[3] ? _GEN3138 : _GEN78;
wire  _GEN3140 = io_x[7] ? _GEN3139 : _GEN3137;
wire  _GEN3141 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3142 = io_x[11] ? _GEN3141 : _GEN67;
wire  _GEN3143 = io_x[3] ? _GEN3142 : _GEN78;
wire  _GEN3144 = io_x[7] ? _GEN3143 : _GEN65;
wire  _GEN3145 = io_x[23] ? _GEN3144 : _GEN3140;
wire  _GEN3146 = io_x[2] ? _GEN3145 : _GEN3136;
wire  _GEN3147 = io_x[16] ? _GEN3146 : _GEN3132;
wire  _GEN3148 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3149 = io_x[11] ? _GEN3148 : _GEN67;
wire  _GEN3150 = io_x[3] ? _GEN66 : _GEN3149;
wire  _GEN3151 = io_x[7] ? _GEN3150 : _GEN65;
wire  _GEN3152 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3153 = io_x[7] ? _GEN3152 : _GEN65;
wire  _GEN3154 = io_x[23] ? _GEN3153 : _GEN3151;
wire  _GEN3155 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3156 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3157 = io_x[11] ? _GEN3156 : _GEN67;
wire  _GEN3158 = io_x[3] ? _GEN78 : _GEN3157;
wire  _GEN3159 = io_x[7] ? _GEN3158 : _GEN3155;
wire  _GEN3160 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN3161 = io_x[23] ? _GEN3160 : _GEN3159;
wire  _GEN3162 = io_x[2] ? _GEN3161 : _GEN3154;
wire  _GEN3163 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3164 = io_x[11] ? _GEN3163 : _GEN67;
wire  _GEN3165 = io_x[3] ? _GEN3164 : _GEN66;
wire  _GEN3166 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3167 = io_x[11] ? _GEN3166 : _GEN67;
wire  _GEN3168 = io_x[3] ? _GEN3167 : _GEN66;
wire  _GEN3169 = io_x[7] ? _GEN3168 : _GEN3165;
wire  _GEN3170 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3171 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3172 = io_x[11] ? _GEN3171 : _GEN76;
wire  _GEN3173 = io_x[3] ? _GEN3172 : _GEN66;
wire  _GEN3174 = io_x[7] ? _GEN3173 : _GEN3170;
wire  _GEN3175 = io_x[23] ? _GEN3174 : _GEN3169;
wire  _GEN3176 = io_x[2] ? _GEN3175 : _GEN573;
wire  _GEN3177 = io_x[16] ? _GEN3176 : _GEN3162;
wire  _GEN3178 = io_x[15] ? _GEN3177 : _GEN3147;
wire  _GEN3179 = io_x[12] ? _GEN3178 : _GEN3126;
wire  _GEN3180 = io_x[10] ? _GEN3179 : _GEN3069;
wire  _GEN3181 = io_x[4] ? _GEN3180 : _GEN3003;
wire  _GEN3182 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3183 = io_x[3] ? _GEN3182 : _GEN66;
wire  _GEN3184 = io_x[7] ? _GEN3183 : _GEN65;
wire  _GEN3185 = io_x[23] ? _GEN81 : _GEN3184;
wire  _GEN3186 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3187 = io_x[11] ? _GEN3186 : _GEN67;
wire  _GEN3188 = io_x[3] ? _GEN78 : _GEN3187;
wire  _GEN3189 = io_x[7] ? _GEN65 : _GEN3188;
wire  _GEN3190 = io_x[23] ? _GEN74 : _GEN3189;
wire  _GEN3191 = io_x[2] ? _GEN3190 : _GEN3185;
wire  _GEN3192 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN3193 = io_x[23] ? _GEN3192 : _GEN74;
wire  _GEN3194 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3195 = io_x[11] ? _GEN3194 : _GEN67;
wire  _GEN3196 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3197 = io_x[11] ? _GEN3196 : _GEN67;
wire  _GEN3198 = io_x[3] ? _GEN3197 : _GEN3195;
wire  _GEN3199 = io_x[7] ? _GEN65 : _GEN3198;
wire  _GEN3200 = io_x[23] ? _GEN81 : _GEN3199;
wire  _GEN3201 = io_x[2] ? _GEN3200 : _GEN3193;
wire  _GEN3202 = io_x[16] ? _GEN3201 : _GEN3191;
wire  _GEN3203 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3204 = io_x[7] ? _GEN65 : _GEN3203;
wire  _GEN3205 = io_x[23] ? _GEN81 : _GEN3204;
wire  _GEN3206 = io_x[2] ? _GEN3205 : _GEN140;
wire  _GEN3207 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN3208 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN3209 = io_x[23] ? _GEN3208 : _GEN3207;
wire  _GEN3210 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3211 = io_x[11] ? _GEN3210 : _GEN67;
wire  _GEN3212 = io_x[3] ? _GEN3211 : _GEN78;
wire  _GEN3213 = io_x[7] ? _GEN65 : _GEN3212;
wire  _GEN3214 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3215 = io_x[3] ? _GEN3214 : _GEN78;
wire  _GEN3216 = io_x[7] ? _GEN84 : _GEN3215;
wire  _GEN3217 = io_x[23] ? _GEN3216 : _GEN3213;
wire  _GEN3218 = io_x[2] ? _GEN3217 : _GEN3209;
wire  _GEN3219 = io_x[16] ? _GEN3218 : _GEN3206;
wire  _GEN3220 = io_x[15] ? _GEN3219 : _GEN3202;
wire  _GEN3221 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3222 = io_x[7] ? _GEN84 : _GEN3221;
wire  _GEN3223 = io_x[23] ? _GEN74 : _GEN3222;
wire  _GEN3224 = io_x[2] ? _GEN3223 : _GEN573;
wire  _GEN3225 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3226 = io_x[3] ? _GEN3225 : _GEN66;
wire  _GEN3227 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3228 = io_x[3] ? _GEN3227 : _GEN66;
wire  _GEN3229 = io_x[7] ? _GEN3228 : _GEN3226;
wire  _GEN3230 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3231 = io_x[3] ? _GEN3230 : _GEN66;
wire  _GEN3232 = io_x[7] ? _GEN3231 : _GEN84;
wire  _GEN3233 = io_x[23] ? _GEN3232 : _GEN3229;
wire  _GEN3234 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3235 = io_x[7] ? _GEN65 : _GEN3234;
wire  _GEN3236 = io_x[23] ? _GEN81 : _GEN3235;
wire  _GEN3237 = io_x[2] ? _GEN3236 : _GEN3233;
wire  _GEN3238 = io_x[16] ? _GEN3237 : _GEN3224;
wire  _GEN3239 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN3240 = io_x[23] ? _GEN74 : _GEN3239;
wire  _GEN3241 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3242 = io_x[3] ? _GEN66 : _GEN3241;
wire  _GEN3243 = io_x[7] ? _GEN65 : _GEN3242;
wire  _GEN3244 = io_x[23] ? _GEN81 : _GEN3243;
wire  _GEN3245 = io_x[2] ? _GEN3244 : _GEN3240;
wire  _GEN3246 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3247 = io_x[11] ? _GEN3246 : _GEN67;
wire  _GEN3248 = io_x[3] ? _GEN3247 : _GEN66;
wire  _GEN3249 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3250 = io_x[7] ? _GEN3249 : _GEN3248;
wire  _GEN3251 = io_x[23] ? _GEN81 : _GEN3250;
wire  _GEN3252 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3253 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3254 = io_x[3] ? _GEN3253 : _GEN66;
wire  _GEN3255 = io_x[7] ? _GEN3254 : _GEN3252;
wire  _GEN3256 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3257 = io_x[7] ? _GEN3256 : _GEN84;
wire  _GEN3258 = io_x[23] ? _GEN3257 : _GEN3255;
wire  _GEN3259 = io_x[2] ? _GEN3258 : _GEN3251;
wire  _GEN3260 = io_x[16] ? _GEN3259 : _GEN3245;
wire  _GEN3261 = io_x[15] ? _GEN3260 : _GEN3238;
wire  _GEN3262 = io_x[12] ? _GEN3261 : _GEN3220;
wire  _GEN3263 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3264 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3265 = io_x[7] ? _GEN3264 : _GEN3263;
wire  _GEN3266 = io_x[23] ? _GEN74 : _GEN3265;
wire  _GEN3267 = io_x[2] ? _GEN3266 : _GEN573;
wire  _GEN3268 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3269 = io_x[3] ? _GEN3268 : _GEN66;
wire  _GEN3270 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3271 = io_x[3] ? _GEN3270 : _GEN66;
wire  _GEN3272 = io_x[7] ? _GEN3271 : _GEN3269;
wire  _GEN3273 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3274 = io_x[3] ? _GEN3273 : _GEN66;
wire  _GEN3275 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3276 = io_x[3] ? _GEN3275 : _GEN66;
wire  _GEN3277 = io_x[7] ? _GEN3276 : _GEN3274;
wire  _GEN3278 = io_x[23] ? _GEN3277 : _GEN3272;
wire  _GEN3279 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3280 = io_x[3] ? _GEN78 : _GEN3279;
wire  _GEN3281 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3282 = io_x[7] ? _GEN3281 : _GEN3280;
wire  _GEN3283 = io_x[23] ? _GEN81 : _GEN3282;
wire  _GEN3284 = io_x[2] ? _GEN3283 : _GEN3278;
wire  _GEN3285 = io_x[16] ? _GEN3284 : _GEN3267;
wire  _GEN3286 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN3287 = io_x[23] ? _GEN3286 : _GEN81;
wire  _GEN3288 = io_x[2] ? _GEN3287 : _GEN140;
wire  _GEN3289 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3290 = io_x[3] ? _GEN3289 : _GEN66;
wire  _GEN3291 = io_x[7] ? _GEN3290 : _GEN65;
wire  _GEN3292 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3293 = io_x[3] ? _GEN3292 : _GEN66;
wire  _GEN3294 = io_x[7] ? _GEN3293 : _GEN65;
wire  _GEN3295 = io_x[23] ? _GEN3294 : _GEN3291;
wire  _GEN3296 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3297 = io_x[11] ? _GEN67 : _GEN3296;
wire  _GEN3298 = io_x[3] ? _GEN3297 : _GEN78;
wire  _GEN3299 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3300 = io_x[3] ? _GEN3299 : _GEN78;
wire  _GEN3301 = io_x[7] ? _GEN3300 : _GEN3298;
wire  _GEN3302 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3303 = io_x[7] ? _GEN3302 : _GEN84;
wire  _GEN3304 = io_x[23] ? _GEN3303 : _GEN3301;
wire  _GEN3305 = io_x[2] ? _GEN3304 : _GEN3295;
wire  _GEN3306 = io_x[16] ? _GEN3305 : _GEN3288;
wire  _GEN3307 = io_x[15] ? _GEN3306 : _GEN3285;
wire  _GEN3308 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3309 = io_x[3] ? _GEN66 : _GEN3308;
wire  _GEN3310 = io_x[7] ? _GEN3309 : _GEN65;
wire  _GEN3311 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN3312 = io_x[23] ? _GEN3311 : _GEN3310;
wire  _GEN3313 = io_x[2] ? _GEN3312 : _GEN140;
wire  _GEN3314 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3315 = io_x[11] ? _GEN67 : _GEN3314;
wire  _GEN3316 = io_x[3] ? _GEN3315 : _GEN66;
wire  _GEN3317 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3318 = io_x[11] ? _GEN67 : _GEN3317;
wire  _GEN3319 = io_x[3] ? _GEN3318 : _GEN66;
wire  _GEN3320 = io_x[7] ? _GEN3319 : _GEN3316;
wire  _GEN3321 = io_x[23] ? _GEN81 : _GEN3320;
wire  _GEN3322 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3323 = io_x[3] ? _GEN66 : _GEN3322;
wire  _GEN3324 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3325 = io_x[3] ? _GEN66 : _GEN3324;
wire  _GEN3326 = io_x[7] ? _GEN3325 : _GEN3323;
wire  _GEN3327 = io_x[23] ? _GEN74 : _GEN3326;
wire  _GEN3328 = io_x[2] ? _GEN3327 : _GEN3321;
wire  _GEN3329 = io_x[16] ? _GEN3328 : _GEN3313;
wire  _GEN3330 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3331 = io_x[7] ? _GEN3330 : _GEN65;
wire  _GEN3332 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3333 = io_x[3] ? _GEN3332 : _GEN66;
wire  _GEN3334 = io_x[7] ? _GEN3333 : _GEN65;
wire  _GEN3335 = io_x[23] ? _GEN3334 : _GEN3331;
wire  _GEN3336 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3337 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3338 = io_x[11] ? _GEN3337 : _GEN67;
wire  _GEN3339 = io_x[3] ? _GEN3338 : _GEN66;
wire  _GEN3340 = io_x[7] ? _GEN3339 : _GEN3336;
wire  _GEN3341 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3342 = io_x[11] ? _GEN67 : _GEN3341;
wire  _GEN3343 = io_x[3] ? _GEN78 : _GEN3342;
wire  _GEN3344 = io_x[7] ? _GEN65 : _GEN3343;
wire  _GEN3345 = io_x[23] ? _GEN3344 : _GEN3340;
wire  _GEN3346 = io_x[2] ? _GEN3345 : _GEN3335;
wire  _GEN3347 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3348 = io_x[3] ? _GEN3347 : _GEN66;
wire  _GEN3349 = io_x[7] ? _GEN3348 : _GEN84;
wire  _GEN3350 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3351 = io_x[11] ? _GEN3350 : _GEN67;
wire  _GEN3352 = io_x[3] ? _GEN3351 : _GEN66;
wire  _GEN3353 = io_x[7] ? _GEN3352 : _GEN84;
wire  _GEN3354 = io_x[23] ? _GEN3353 : _GEN3349;
wire  _GEN3355 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3356 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3357 = io_x[3] ? _GEN3356 : _GEN3355;
wire  _GEN3358 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3359 = io_x[11] ? _GEN3358 : _GEN67;
wire  _GEN3360 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3361 = io_x[11] ? _GEN3360 : _GEN67;
wire  _GEN3362 = io_x[3] ? _GEN3361 : _GEN3359;
wire  _GEN3363 = io_x[7] ? _GEN3362 : _GEN3357;
wire  _GEN3364 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3365 = io_x[11] ? _GEN67 : _GEN3364;
wire  _GEN3366 = io_x[3] ? _GEN78 : _GEN3365;
wire  _GEN3367 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3368 = io_x[11] ? _GEN3367 : _GEN67;
wire  _GEN3369 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3370 = io_x[11] ? _GEN3369 : _GEN67;
wire  _GEN3371 = io_x[3] ? _GEN3370 : _GEN3368;
wire  _GEN3372 = io_x[7] ? _GEN3371 : _GEN3366;
wire  _GEN3373 = io_x[23] ? _GEN3372 : _GEN3363;
wire  _GEN3374 = io_x[2] ? _GEN3373 : _GEN3354;
wire  _GEN3375 = io_x[16] ? _GEN3374 : _GEN3346;
wire  _GEN3376 = io_x[15] ? _GEN3375 : _GEN3329;
wire  _GEN3377 = io_x[12] ? _GEN3376 : _GEN3307;
wire  _GEN3378 = io_x[10] ? _GEN3377 : _GEN3262;
wire  _GEN3379 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3380 = io_x[11] ? _GEN3379 : _GEN67;
wire  _GEN3381 = io_x[3] ? _GEN66 : _GEN3380;
wire  _GEN3382 = io_x[7] ? _GEN84 : _GEN3381;
wire  _GEN3383 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3384 = io_x[7] ? _GEN3383 : _GEN65;
wire  _GEN3385 = io_x[23] ? _GEN3384 : _GEN3382;
wire  _GEN3386 = io_x[2] ? _GEN3385 : _GEN140;
wire  _GEN3387 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN3388 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3389 = io_x[7] ? _GEN65 : _GEN3388;
wire  _GEN3390 = io_x[23] ? _GEN3389 : _GEN3387;
wire  _GEN3391 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3392 = io_x[11] ? _GEN3391 : _GEN67;
wire  _GEN3393 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3394 = io_x[3] ? _GEN3393 : _GEN3392;
wire  _GEN3395 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3396 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3397 = io_x[3] ? _GEN3396 : _GEN3395;
wire  _GEN3398 = io_x[7] ? _GEN3397 : _GEN3394;
wire  _GEN3399 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3400 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3401 = io_x[11] ? _GEN3400 : _GEN67;
wire  _GEN3402 = io_x[3] ? _GEN3401 : _GEN78;
wire  _GEN3403 = io_x[7] ? _GEN3402 : _GEN3399;
wire  _GEN3404 = io_x[23] ? _GEN3403 : _GEN3398;
wire  _GEN3405 = io_x[2] ? _GEN3404 : _GEN3390;
wire  _GEN3406 = io_x[16] ? _GEN3405 : _GEN3386;
wire  _GEN3407 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN3408 = io_x[23] ? _GEN81 : _GEN3407;
wire  _GEN3409 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN3410 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3411 = io_x[11] ? _GEN3410 : _GEN67;
wire  _GEN3412 = io_x[3] ? _GEN66 : _GEN3411;
wire  _GEN3413 = io_x[7] ? _GEN65 : _GEN3412;
wire  _GEN3414 = io_x[23] ? _GEN3413 : _GEN3409;
wire  _GEN3415 = io_x[2] ? _GEN3414 : _GEN3408;
wire  _GEN3416 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3417 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3418 = io_x[3] ? _GEN3417 : _GEN3416;
wire  _GEN3419 = io_x[7] ? _GEN3418 : _GEN65;
wire  _GEN3420 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3421 = io_x[7] ? _GEN3420 : _GEN65;
wire  _GEN3422 = io_x[23] ? _GEN3421 : _GEN3419;
wire  _GEN3423 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3424 = io_x[3] ? _GEN3423 : _GEN78;
wire  _GEN3425 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3426 = io_x[3] ? _GEN3425 : _GEN66;
wire  _GEN3427 = io_x[7] ? _GEN3426 : _GEN3424;
wire  _GEN3428 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3429 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3430 = io_x[7] ? _GEN3429 : _GEN3428;
wire  _GEN3431 = io_x[23] ? _GEN3430 : _GEN3427;
wire  _GEN3432 = io_x[2] ? _GEN3431 : _GEN3422;
wire  _GEN3433 = io_x[16] ? _GEN3432 : _GEN3415;
wire  _GEN3434 = io_x[15] ? _GEN3433 : _GEN3406;
wire  _GEN3435 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3436 = io_x[3] ? _GEN3435 : _GEN78;
wire  _GEN3437 = io_x[7] ? _GEN3436 : _GEN65;
wire  _GEN3438 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3439 = io_x[11] ? _GEN3438 : _GEN67;
wire  _GEN3440 = io_x[3] ? _GEN66 : _GEN3439;
wire  _GEN3441 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3442 = io_x[7] ? _GEN3441 : _GEN3440;
wire  _GEN3443 = io_x[23] ? _GEN3442 : _GEN3437;
wire  _GEN3444 = io_x[2] ? _GEN3443 : _GEN140;
wire  _GEN3445 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3446 = io_x[3] ? _GEN3445 : _GEN78;
wire  _GEN3447 = io_x[7] ? _GEN3446 : _GEN65;
wire  _GEN3448 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3449 = io_x[3] ? _GEN3448 : _GEN66;
wire  _GEN3450 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3451 = io_x[7] ? _GEN3450 : _GEN3449;
wire  _GEN3452 = io_x[23] ? _GEN3451 : _GEN3447;
wire  _GEN3453 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3454 = io_x[3] ? _GEN3453 : _GEN66;
wire  _GEN3455 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3456 = io_x[3] ? _GEN3455 : _GEN78;
wire  _GEN3457 = io_x[7] ? _GEN3456 : _GEN3454;
wire  _GEN3458 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3459 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3460 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3461 = io_x[3] ? _GEN3460 : _GEN3459;
wire  _GEN3462 = io_x[7] ? _GEN3461 : _GEN3458;
wire  _GEN3463 = io_x[23] ? _GEN3462 : _GEN3457;
wire  _GEN3464 = io_x[2] ? _GEN3463 : _GEN3452;
wire  _GEN3465 = io_x[16] ? _GEN3464 : _GEN3444;
wire  _GEN3466 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3467 = io_x[3] ? _GEN3466 : _GEN66;
wire  _GEN3468 = io_x[7] ? _GEN3467 : _GEN65;
wire  _GEN3469 = io_x[23] ? _GEN81 : _GEN3468;
wire  _GEN3470 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3471 = io_x[3] ? _GEN66 : _GEN3470;
wire  _GEN3472 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3473 = io_x[3] ? _GEN66 : _GEN3472;
wire  _GEN3474 = io_x[7] ? _GEN3473 : _GEN3471;
wire  _GEN3475 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3476 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3477 = io_x[11] ? _GEN3476 : _GEN3475;
wire  _GEN3478 = io_x[3] ? _GEN3477 : _GEN66;
wire  _GEN3479 = io_x[7] ? _GEN3478 : _GEN84;
wire  _GEN3480 = io_x[23] ? _GEN3479 : _GEN3474;
wire  _GEN3481 = io_x[2] ? _GEN3480 : _GEN3469;
wire  _GEN3482 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3483 = io_x[11] ? _GEN3482 : _GEN67;
wire  _GEN3484 = io_x[3] ? _GEN78 : _GEN3483;
wire  _GEN3485 = io_x[7] ? _GEN3484 : _GEN65;
wire  _GEN3486 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3487 = io_x[3] ? _GEN3486 : _GEN66;
wire  _GEN3488 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3489 = io_x[3] ? _GEN3488 : _GEN66;
wire  _GEN3490 = io_x[7] ? _GEN3489 : _GEN3487;
wire  _GEN3491 = io_x[23] ? _GEN3490 : _GEN3485;
wire  _GEN3492 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3493 = io_x[11] ? _GEN3492 : _GEN76;
wire  _GEN3494 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3495 = io_x[11] ? _GEN67 : _GEN3494;
wire  _GEN3496 = io_x[3] ? _GEN3495 : _GEN3493;
wire  _GEN3497 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3498 = io_x[11] ? _GEN67 : _GEN3497;
wire  _GEN3499 = io_x[3] ? _GEN3498 : _GEN66;
wire  _GEN3500 = io_x[7] ? _GEN3499 : _GEN3496;
wire  _GEN3501 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3502 = io_x[11] ? _GEN67 : _GEN3501;
wire  _GEN3503 = io_x[3] ? _GEN66 : _GEN3502;
wire  _GEN3504 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3505 = io_x[11] ? _GEN3504 : _GEN67;
wire  _GEN3506 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3507 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3508 = io_x[11] ? _GEN3507 : _GEN3506;
wire  _GEN3509 = io_x[3] ? _GEN3508 : _GEN3505;
wire  _GEN3510 = io_x[7] ? _GEN3509 : _GEN3503;
wire  _GEN3511 = io_x[23] ? _GEN3510 : _GEN3500;
wire  _GEN3512 = io_x[2] ? _GEN3511 : _GEN3491;
wire  _GEN3513 = io_x[16] ? _GEN3512 : _GEN3481;
wire  _GEN3514 = io_x[15] ? _GEN3513 : _GEN3465;
wire  _GEN3515 = io_x[12] ? _GEN3514 : _GEN3434;
wire  _GEN3516 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3517 = io_x[3] ? _GEN66 : _GEN3516;
wire  _GEN3518 = io_x[7] ? _GEN65 : _GEN3517;
wire  _GEN3519 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3520 = io_x[3] ? _GEN66 : _GEN3519;
wire  _GEN3521 = io_x[7] ? _GEN65 : _GEN3520;
wire  _GEN3522 = io_x[23] ? _GEN3521 : _GEN3518;
wire  _GEN3523 = io_x[2] ? _GEN3522 : _GEN140;
wire  _GEN3524 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3525 = io_x[3] ? _GEN3524 : _GEN78;
wire  _GEN3526 = io_x[7] ? _GEN3525 : _GEN84;
wire  _GEN3527 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN3528 = io_x[23] ? _GEN3527 : _GEN3526;
wire  _GEN3529 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3530 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3531 = io_x[3] ? _GEN3530 : _GEN3529;
wire  _GEN3532 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3533 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3534 = io_x[11] ? _GEN3533 : _GEN67;
wire  _GEN3535 = io_x[3] ? _GEN3534 : _GEN3532;
wire  _GEN3536 = io_x[7] ? _GEN3535 : _GEN3531;
wire  _GEN3537 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3538 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3539 = io_x[3] ? _GEN3538 : _GEN3537;
wire  _GEN3540 = io_x[7] ? _GEN65 : _GEN3539;
wire  _GEN3541 = io_x[23] ? _GEN3540 : _GEN3536;
wire  _GEN3542 = io_x[2] ? _GEN3541 : _GEN3528;
wire  _GEN3543 = io_x[16] ? _GEN3542 : _GEN3523;
wire  _GEN3544 = io_x[7] ? _GEN65 : _GEN84;
wire  _GEN3545 = io_x[3] ? _GEN66 : _GEN78;
wire  _GEN3546 = io_x[7] ? _GEN3545 : _GEN65;
wire  _GEN3547 = io_x[23] ? _GEN3546 : _GEN3544;
wire  _GEN3548 = io_x[7] ? _GEN84 : _GEN65;
wire  _GEN3549 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3550 = io_x[11] ? _GEN3549 : _GEN67;
wire  _GEN3551 = io_x[3] ? _GEN66 : _GEN3550;
wire  _GEN3552 = io_x[3] ? _GEN78 : _GEN66;
wire  _GEN3553 = io_x[7] ? _GEN3552 : _GEN3551;
wire  _GEN3554 = io_x[23] ? _GEN3553 : _GEN3548;
wire  _GEN3555 = io_x[2] ? _GEN3554 : _GEN3547;
wire  _GEN3556 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3557 = io_x[11] ? _GEN3556 : _GEN67;
wire  _GEN3558 = io_x[3] ? _GEN3557 : _GEN66;
wire  _GEN3559 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3560 = io_x[3] ? _GEN3559 : _GEN66;
wire  _GEN3561 = io_x[7] ? _GEN3560 : _GEN3558;
wire  _GEN3562 = io_x[23] ? _GEN81 : _GEN3561;
wire  _GEN3563 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3564 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3565 = io_x[11] ? _GEN3564 : _GEN76;
wire  _GEN3566 = io_x[3] ? _GEN3565 : _GEN3563;
wire  _GEN3567 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3568 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3569 = io_x[11] ? _GEN3568 : _GEN3567;
wire  _GEN3570 = io_x[3] ? _GEN3569 : _GEN78;
wire  _GEN3571 = io_x[7] ? _GEN3570 : _GEN3566;
wire  _GEN3572 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3573 = io_x[3] ? _GEN3572 : _GEN78;
wire  _GEN3574 = io_x[7] ? _GEN65 : _GEN3573;
wire  _GEN3575 = io_x[23] ? _GEN3574 : _GEN3571;
wire  _GEN3576 = io_x[2] ? _GEN3575 : _GEN3562;
wire  _GEN3577 = io_x[16] ? _GEN3576 : _GEN3555;
wire  _GEN3578 = io_x[15] ? _GEN3577 : _GEN3543;
wire  _GEN3579 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3580 = io_x[11] ? _GEN3579 : _GEN67;
wire  _GEN3581 = io_x[3] ? _GEN3580 : _GEN66;
wire  _GEN3582 = io_x[7] ? _GEN3581 : _GEN65;
wire  _GEN3583 = io_x[23] ? _GEN3582 : _GEN81;
wire  _GEN3584 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3585 = io_x[3] ? _GEN3584 : _GEN66;
wire  _GEN3586 = io_x[7] ? _GEN3585 : _GEN65;
wire  _GEN3587 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3588 = io_x[11] ? _GEN67 : _GEN3587;
wire  _GEN3589 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3590 = io_x[11] ? _GEN67 : _GEN3589;
wire  _GEN3591 = io_x[3] ? _GEN3590 : _GEN3588;
wire  _GEN3592 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3593 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3594 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3595 = io_x[11] ? _GEN3594 : _GEN3593;
wire  _GEN3596 = io_x[3] ? _GEN3595 : _GEN3592;
wire  _GEN3597 = io_x[7] ? _GEN3596 : _GEN3591;
wire  _GEN3598 = io_x[23] ? _GEN3597 : _GEN3586;
wire  _GEN3599 = io_x[2] ? _GEN3598 : _GEN3583;
wire  _GEN3600 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3601 = io_x[11] ? _GEN76 : _GEN3600;
wire  _GEN3602 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3603 = io_x[11] ? _GEN3602 : _GEN76;
wire  _GEN3604 = io_x[3] ? _GEN3603 : _GEN3601;
wire  _GEN3605 = io_x[7] ? _GEN3604 : _GEN84;
wire  _GEN3606 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3607 = io_x[3] ? _GEN66 : _GEN3606;
wire  _GEN3608 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3609 = io_x[3] ? _GEN3608 : _GEN66;
wire  _GEN3610 = io_x[7] ? _GEN3609 : _GEN3607;
wire  _GEN3611 = io_x[23] ? _GEN3610 : _GEN3605;
wire  _GEN3612 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3613 = io_x[11] ? _GEN67 : _GEN3612;
wire  _GEN3614 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3615 = io_x[11] ? _GEN76 : _GEN3614;
wire  _GEN3616 = io_x[3] ? _GEN3615 : _GEN3613;
wire  _GEN3617 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3618 = io_x[11] ? _GEN3617 : _GEN76;
wire  _GEN3619 = io_x[3] ? _GEN3618 : _GEN66;
wire  _GEN3620 = io_x[7] ? _GEN3619 : _GEN3616;
wire  _GEN3621 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3622 = io_x[11] ? _GEN67 : _GEN3621;
wire  _GEN3623 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3624 = io_x[11] ? _GEN76 : _GEN3623;
wire  _GEN3625 = io_x[3] ? _GEN3624 : _GEN3622;
wire  _GEN3626 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3627 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3628 = io_x[11] ? _GEN3627 : _GEN3626;
wire  _GEN3629 = io_x[3] ? _GEN3628 : _GEN66;
wire  _GEN3630 = io_x[7] ? _GEN3629 : _GEN3625;
wire  _GEN3631 = io_x[23] ? _GEN3630 : _GEN3620;
wire  _GEN3632 = io_x[2] ? _GEN3631 : _GEN3611;
wire  _GEN3633 = io_x[16] ? _GEN3632 : _GEN3599;
wire  _GEN3634 = io_x[11] ? _GEN67 : _GEN76;
wire  _GEN3635 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3636 = io_x[11] ? _GEN3635 : _GEN67;
wire  _GEN3637 = io_x[3] ? _GEN3636 : _GEN3634;
wire  _GEN3638 = io_x[7] ? _GEN3637 : _GEN84;
wire  _GEN3639 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3640 = io_x[11] ? _GEN3639 : _GEN67;
wire  _GEN3641 = io_x[3] ? _GEN3640 : _GEN78;
wire  _GEN3642 = io_x[7] ? _GEN3641 : _GEN84;
wire  _GEN3643 = io_x[23] ? _GEN3642 : _GEN3638;
wire  _GEN3644 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3645 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3646 = io_x[11] ? _GEN3645 : _GEN3644;
wire  _GEN3647 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3648 = io_x[11] ? _GEN3647 : _GEN67;
wire  _GEN3649 = io_x[3] ? _GEN3648 : _GEN3646;
wire  _GEN3650 = io_x[7] ? _GEN3649 : _GEN84;
wire  _GEN3651 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3652 = io_x[11] ? _GEN76 : _GEN3651;
wire  _GEN3653 = io_x[3] ? _GEN78 : _GEN3652;
wire  _GEN3654 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3655 = io_x[11] ? _GEN3654 : _GEN67;
wire  _GEN3656 = io_x[3] ? _GEN3655 : _GEN78;
wire  _GEN3657 = io_x[7] ? _GEN3656 : _GEN3653;
wire  _GEN3658 = io_x[23] ? _GEN3657 : _GEN3650;
wire  _GEN3659 = io_x[2] ? _GEN3658 : _GEN3643;
wire  _GEN3660 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3661 = io_x[3] ? _GEN66 : _GEN3660;
wire  _GEN3662 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3663 = io_x[11] ? _GEN3662 : _GEN76;
wire  _GEN3664 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3665 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3666 = io_x[11] ? _GEN3665 : _GEN3664;
wire  _GEN3667 = io_x[3] ? _GEN3666 : _GEN3663;
wire  _GEN3668 = io_x[7] ? _GEN3667 : _GEN3661;
wire  _GEN3669 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3670 = io_x[11] ? _GEN3669 : _GEN76;
wire  _GEN3671 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3672 = io_x[11] ? _GEN3671 : _GEN67;
wire  _GEN3673 = io_x[3] ? _GEN3672 : _GEN3670;
wire  _GEN3674 = io_x[7] ? _GEN3673 : _GEN84;
wire  _GEN3675 = io_x[23] ? _GEN3674 : _GEN3668;
wire  _GEN3676 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3677 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3678 = io_x[11] ? _GEN3677 : _GEN76;
wire  _GEN3679 = io_x[3] ? _GEN3678 : _GEN3676;
wire  _GEN3680 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3681 = io_x[11] ? _GEN67 : _GEN3680;
wire  _GEN3682 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3683 = io_x[11] ? _GEN3682 : _GEN67;
wire  _GEN3684 = io_x[3] ? _GEN3683 : _GEN3681;
wire  _GEN3685 = io_x[7] ? _GEN3684 : _GEN3679;
wire  _GEN3686 = io_x[11] ? _GEN76 : _GEN67;
wire  _GEN3687 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3688 = io_x[11] ? _GEN3687 : _GEN67;
wire  _GEN3689 = io_x[3] ? _GEN3688 : _GEN3686;
wire  _GEN3690 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3691 = io_x[11] ? _GEN76 : _GEN3690;
wire  _GEN3692 = io_x[27] ? _GEN69 : _GEN68;
wire  _GEN3693 = io_x[27] ? _GEN68 : _GEN69;
wire  _GEN3694 = io_x[11] ? _GEN3693 : _GEN3692;
wire  _GEN3695 = io_x[3] ? _GEN3694 : _GEN3691;
wire  _GEN3696 = io_x[7] ? _GEN3695 : _GEN3689;
wire  _GEN3697 = io_x[23] ? _GEN3696 : _GEN3685;
wire  _GEN3698 = io_x[2] ? _GEN3697 : _GEN3675;
wire  _GEN3699 = io_x[16] ? _GEN3698 : _GEN3659;
wire  _GEN3700 = io_x[15] ? _GEN3699 : _GEN3633;
wire  _GEN3701 = io_x[12] ? _GEN3700 : _GEN3578;
wire  _GEN3702 = io_x[10] ? _GEN3701 : _GEN3515;
wire  _GEN3703 = io_x[4] ? _GEN3702 : _GEN3378;
wire  _GEN3704 = io_x[8] ? _GEN3703 : _GEN3181;
wire  _GEN3705 = io_x[28] ? _GEN3704 : _GEN2849;
wire  _GEN3706 = io_x[22] ? _GEN3705 : _GEN1797;
assign io_y[9] = _GEN3706;
wire  _GEN3707 = 1'b1;
wire  _GEN3708 = 1'b0;
wire  _GEN3709 = 1'b1;
wire  _GEN3710 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN3711 = 1'b1;
wire  _GEN3712 = io_x[10] ? _GEN3711 : _GEN3710;
wire  _GEN3713 = 1'b1;
wire  _GEN3714 = io_x[23] ? _GEN3713 : _GEN3712;
wire  _GEN3715 = io_x[16] ? _GEN3714 : _GEN3707;
wire  _GEN3716 = 1'b0;
wire  _GEN3717 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN3718 = io_x[23] ? _GEN3713 : _GEN3717;
wire  _GEN3719 = 1'b0;
wire  _GEN3720 = 1'b1;
wire  _GEN3721 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3722 = io_x[14] ? _GEN3721 : _GEN3709;
wire  _GEN3723 = io_x[10] ? _GEN3722 : _GEN3716;
wire  _GEN3724 = io_x[23] ? _GEN3713 : _GEN3723;
wire  _GEN3725 = io_x[16] ? _GEN3724 : _GEN3718;
wire  _GEN3726 = io_x[12] ? _GEN3725 : _GEN3715;
wire  _GEN3727 = 1'b0;
wire  _GEN3728 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN3729 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3730 = io_x[14] ? _GEN3729 : _GEN3709;
wire  _GEN3731 = io_x[10] ? _GEN3716 : _GEN3730;
wire  _GEN3732 = io_x[23] ? _GEN3731 : _GEN3728;
wire  _GEN3733 = io_x[16] ? _GEN3732 : _GEN3727;
wire  _GEN3734 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN3735 = io_x[10] ? _GEN3734 : _GEN3711;
wire  _GEN3736 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN3737 = io_x[23] ? _GEN3736 : _GEN3735;
wire  _GEN3738 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3739 = io_x[14] ? _GEN3738 : _GEN3709;
wire  _GEN3740 = io_x[10] ? _GEN3739 : _GEN3711;
wire  _GEN3741 = 1'b0;
wire  _GEN3742 = io_x[23] ? _GEN3741 : _GEN3740;
wire  _GEN3743 = io_x[16] ? _GEN3742 : _GEN3737;
wire  _GEN3744 = io_x[12] ? _GEN3743 : _GEN3733;
wire  _GEN3745 = io_x[2] ? _GEN3744 : _GEN3726;
wire  _GEN3746 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN3747 = io_x[10] ? _GEN3746 : _GEN3711;
wire  _GEN3748 = io_x[23] ? _GEN3713 : _GEN3747;
wire  _GEN3749 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3750 = io_x[14] ? _GEN3749 : _GEN3708;
wire  _GEN3751 = io_x[10] ? _GEN3750 : _GEN3711;
wire  _GEN3752 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN3753 = io_x[10] ? _GEN3752 : _GEN3711;
wire  _GEN3754 = io_x[23] ? _GEN3753 : _GEN3751;
wire  _GEN3755 = io_x[16] ? _GEN3754 : _GEN3748;
wire  _GEN3756 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN3757 = io_x[10] ? _GEN3756 : _GEN3716;
wire  _GEN3758 = io_x[23] ? _GEN3713 : _GEN3757;
wire  _GEN3759 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3760 = io_x[14] ? _GEN3759 : _GEN3709;
wire  _GEN3761 = io_x[10] ? _GEN3760 : _GEN3716;
wire  _GEN3762 = io_x[23] ? _GEN3741 : _GEN3761;
wire  _GEN3763 = io_x[16] ? _GEN3762 : _GEN3758;
wire  _GEN3764 = io_x[12] ? _GEN3763 : _GEN3755;
wire  _GEN3765 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3766 = io_x[14] ? _GEN3765 : _GEN3709;
wire  _GEN3767 = io_x[10] ? _GEN3711 : _GEN3766;
wire  _GEN3768 = io_x[23] ? _GEN3713 : _GEN3767;
wire  _GEN3769 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3770 = io_x[14] ? _GEN3769 : _GEN3709;
wire  _GEN3771 = io_x[10] ? _GEN3770 : _GEN3711;
wire  _GEN3772 = io_x[23] ? _GEN3741 : _GEN3771;
wire  _GEN3773 = io_x[16] ? _GEN3772 : _GEN3768;
wire  _GEN3774 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN3775 = io_x[10] ? _GEN3774 : _GEN3716;
wire  _GEN3776 = io_x[23] ? _GEN3775 : _GEN3741;
wire  _GEN3777 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3778 = io_x[14] ? _GEN3777 : _GEN3709;
wire  _GEN3779 = io_x[10] ? _GEN3778 : _GEN3716;
wire  _GEN3780 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3781 = io_x[14] ? _GEN3780 : _GEN3709;
wire  _GEN3782 = io_x[10] ? _GEN3716 : _GEN3781;
wire  _GEN3783 = io_x[23] ? _GEN3782 : _GEN3779;
wire  _GEN3784 = io_x[16] ? _GEN3783 : _GEN3776;
wire  _GEN3785 = io_x[12] ? _GEN3784 : _GEN3773;
wire  _GEN3786 = io_x[2] ? _GEN3785 : _GEN3764;
wire  _GEN3787 = io_x[9] ? _GEN3786 : _GEN3745;
wire  _GEN3788 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN3789 = io_x[10] ? _GEN3711 : _GEN3788;
wire  _GEN3790 = io_x[23] ? _GEN3741 : _GEN3789;
wire  _GEN3791 = io_x[16] ? _GEN3727 : _GEN3790;
wire  _GEN3792 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3793 = io_x[14] ? _GEN3709 : _GEN3792;
wire  _GEN3794 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN3795 = io_x[10] ? _GEN3794 : _GEN3793;
wire  _GEN3796 = io_x[23] ? _GEN3713 : _GEN3795;
wire  _GEN3797 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3798 = io_x[14] ? _GEN3709 : _GEN3797;
wire  _GEN3799 = io_x[10] ? _GEN3716 : _GEN3798;
wire  _GEN3800 = io_x[23] ? _GEN3741 : _GEN3799;
wire  _GEN3801 = io_x[16] ? _GEN3800 : _GEN3796;
wire  _GEN3802 = io_x[12] ? _GEN3801 : _GEN3791;
wire  _GEN3803 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3804 = io_x[14] ? _GEN3803 : _GEN3709;
wire  _GEN3805 = io_x[10] ? _GEN3804 : _GEN3711;
wire  _GEN3806 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN3807 = io_x[10] ? _GEN3806 : _GEN3711;
wire  _GEN3808 = io_x[23] ? _GEN3807 : _GEN3805;
wire  _GEN3809 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN3810 = io_x[10] ? _GEN3716 : _GEN3809;
wire  _GEN3811 = io_x[23] ? _GEN3741 : _GEN3810;
wire  _GEN3812 = io_x[16] ? _GEN3811 : _GEN3808;
wire  _GEN3813 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN3814 = io_x[10] ? _GEN3813 : _GEN3716;
wire  _GEN3815 = io_x[23] ? _GEN3814 : _GEN3741;
wire  _GEN3816 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3817 = io_x[14] ? _GEN3816 : _GEN3709;
wire  _GEN3818 = io_x[10] ? _GEN3817 : _GEN3711;
wire  _GEN3819 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN3820 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN3821 = io_x[10] ? _GEN3820 : _GEN3819;
wire  _GEN3822 = io_x[23] ? _GEN3821 : _GEN3818;
wire  _GEN3823 = io_x[16] ? _GEN3822 : _GEN3815;
wire  _GEN3824 = io_x[12] ? _GEN3823 : _GEN3812;
wire  _GEN3825 = io_x[2] ? _GEN3824 : _GEN3802;
wire  _GEN3826 = io_x[23] ? _GEN3741 : _GEN3713;
wire  _GEN3827 = io_x[16] ? _GEN3826 : _GEN3727;
wire  _GEN3828 = io_x[23] ? _GEN3713 : _GEN3741;
wire  _GEN3829 = io_x[16] ? _GEN3828 : _GEN3707;
wire  _GEN3830 = io_x[12] ? _GEN3829 : _GEN3827;
wire  _GEN3831 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3832 = io_x[14] ? _GEN3708 : _GEN3831;
wire  _GEN3833 = io_x[10] ? _GEN3832 : _GEN3711;
wire  _GEN3834 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3835 = io_x[14] ? _GEN3709 : _GEN3834;
wire  _GEN3836 = io_x[10] ? _GEN3835 : _GEN3711;
wire  _GEN3837 = io_x[23] ? _GEN3836 : _GEN3833;
wire  _GEN3838 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3839 = io_x[14] ? _GEN3838 : _GEN3709;
wire  _GEN3840 = io_x[10] ? _GEN3716 : _GEN3839;
wire  _GEN3841 = io_x[23] ? _GEN3741 : _GEN3840;
wire  _GEN3842 = io_x[16] ? _GEN3841 : _GEN3837;
wire  _GEN3843 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN3844 = io_x[10] ? _GEN3843 : _GEN3711;
wire  _GEN3845 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3846 = io_x[14] ? _GEN3709 : _GEN3845;
wire  _GEN3847 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN3848 = io_x[10] ? _GEN3847 : _GEN3846;
wire  _GEN3849 = io_x[23] ? _GEN3848 : _GEN3844;
wire  _GEN3850 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3851 = io_x[14] ? _GEN3850 : _GEN3709;
wire  _GEN3852 = io_x[10] ? _GEN3851 : _GEN3711;
wire  _GEN3853 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3854 = io_x[14] ? _GEN3853 : _GEN3708;
wire  _GEN3855 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN3856 = io_x[10] ? _GEN3855 : _GEN3854;
wire  _GEN3857 = io_x[23] ? _GEN3856 : _GEN3852;
wire  _GEN3858 = io_x[16] ? _GEN3857 : _GEN3849;
wire  _GEN3859 = io_x[12] ? _GEN3858 : _GEN3842;
wire  _GEN3860 = io_x[2] ? _GEN3859 : _GEN3830;
wire  _GEN3861 = io_x[9] ? _GEN3860 : _GEN3825;
wire  _GEN3862 = io_x[13] ? _GEN3861 : _GEN3787;
wire  _GEN3863 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN3864 = io_x[23] ? _GEN3713 : _GEN3863;
wire  _GEN3865 = io_x[16] ? _GEN3707 : _GEN3864;
wire  _GEN3866 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN3867 = io_x[23] ? _GEN3713 : _GEN3866;
wire  _GEN3868 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3869 = io_x[14] ? _GEN3868 : _GEN3709;
wire  _GEN3870 = io_x[10] ? _GEN3716 : _GEN3869;
wire  _GEN3871 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN3872 = io_x[23] ? _GEN3871 : _GEN3870;
wire  _GEN3873 = io_x[16] ? _GEN3872 : _GEN3867;
wire  _GEN3874 = io_x[12] ? _GEN3873 : _GEN3865;
wire  _GEN3875 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN3876 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN3877 = io_x[23] ? _GEN3876 : _GEN3875;
wire  _GEN3878 = io_x[16] ? _GEN3877 : _GEN3727;
wire  _GEN3879 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3880 = io_x[14] ? _GEN3708 : _GEN3879;
wire  _GEN3881 = io_x[10] ? _GEN3880 : _GEN3716;
wire  _GEN3882 = io_x[23] ? _GEN3881 : _GEN3741;
wire  _GEN3883 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3884 = io_x[14] ? _GEN3883 : _GEN3709;
wire  _GEN3885 = io_x[10] ? _GEN3884 : _GEN3711;
wire  _GEN3886 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3887 = io_x[14] ? _GEN3708 : _GEN3886;
wire  _GEN3888 = io_x[10] ? _GEN3887 : _GEN3711;
wire  _GEN3889 = io_x[23] ? _GEN3888 : _GEN3885;
wire  _GEN3890 = io_x[16] ? _GEN3889 : _GEN3882;
wire  _GEN3891 = io_x[12] ? _GEN3890 : _GEN3878;
wire  _GEN3892 = io_x[2] ? _GEN3891 : _GEN3874;
wire  _GEN3893 = 1'b1;
wire  _GEN3894 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3895 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3896 = io_x[14] ? _GEN3895 : _GEN3894;
wire  _GEN3897 = io_x[10] ? _GEN3896 : _GEN3711;
wire  _GEN3898 = io_x[23] ? _GEN3713 : _GEN3897;
wire  _GEN3899 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN3900 = io_x[23] ? _GEN3899 : _GEN3713;
wire  _GEN3901 = io_x[16] ? _GEN3900 : _GEN3898;
wire  _GEN3902 = io_x[12] ? _GEN3901 : _GEN3893;
wire  _GEN3903 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN3904 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN3905 = io_x[23] ? _GEN3904 : _GEN3903;
wire  _GEN3906 = io_x[16] ? _GEN3905 : _GEN3727;
wire  _GEN3907 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3908 = io_x[14] ? _GEN3907 : _GEN3708;
wire  _GEN3909 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN3910 = io_x[10] ? _GEN3909 : _GEN3908;
wire  _GEN3911 = io_x[23] ? _GEN3741 : _GEN3910;
wire  _GEN3912 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3913 = io_x[14] ? _GEN3708 : _GEN3912;
wire  _GEN3914 = io_x[10] ? _GEN3913 : _GEN3711;
wire  _GEN3915 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN3916 = io_x[23] ? _GEN3915 : _GEN3914;
wire  _GEN3917 = io_x[16] ? _GEN3916 : _GEN3911;
wire  _GEN3918 = io_x[12] ? _GEN3917 : _GEN3906;
wire  _GEN3919 = io_x[2] ? _GEN3918 : _GEN3902;
wire  _GEN3920 = io_x[9] ? _GEN3919 : _GEN3892;
wire  _GEN3921 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3922 = io_x[14] ? _GEN3708 : _GEN3921;
wire  _GEN3923 = io_x[10] ? _GEN3922 : _GEN3711;
wire  _GEN3924 = io_x[23] ? _GEN3713 : _GEN3923;
wire  _GEN3925 = io_x[16] ? _GEN3707 : _GEN3924;
wire  _GEN3926 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3927 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3928 = io_x[14] ? _GEN3927 : _GEN3926;
wire  _GEN3929 = io_x[10] ? _GEN3928 : _GEN3711;
wire  _GEN3930 = io_x[23] ? _GEN3713 : _GEN3929;
wire  _GEN3931 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3932 = io_x[14] ? _GEN3931 : _GEN3708;
wire  _GEN3933 = io_x[10] ? _GEN3932 : _GEN3716;
wire  _GEN3934 = io_x[23] ? _GEN3933 : _GEN3741;
wire  _GEN3935 = io_x[16] ? _GEN3934 : _GEN3930;
wire  _GEN3936 = io_x[12] ? _GEN3935 : _GEN3925;
wire  _GEN3937 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN3938 = io_x[23] ? _GEN3937 : _GEN3741;
wire  _GEN3939 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3940 = io_x[14] ? _GEN3939 : _GEN3709;
wire  _GEN3941 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN3942 = io_x[10] ? _GEN3941 : _GEN3940;
wire  _GEN3943 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN3944 = io_x[10] ? _GEN3943 : _GEN3711;
wire  _GEN3945 = io_x[23] ? _GEN3944 : _GEN3942;
wire  _GEN3946 = io_x[16] ? _GEN3945 : _GEN3938;
wire  _GEN3947 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3948 = io_x[14] ? _GEN3947 : _GEN3709;
wire  _GEN3949 = io_x[10] ? _GEN3948 : _GEN3711;
wire  _GEN3950 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3951 = io_x[14] ? _GEN3950 : _GEN3709;
wire  _GEN3952 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3953 = io_x[14] ? _GEN3952 : _GEN3709;
wire  _GEN3954 = io_x[10] ? _GEN3953 : _GEN3951;
wire  _GEN3955 = io_x[23] ? _GEN3954 : _GEN3949;
wire  _GEN3956 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3957 = io_x[14] ? _GEN3956 : _GEN3709;
wire  _GEN3958 = io_x[10] ? _GEN3957 : _GEN3711;
wire  _GEN3959 = io_x[23] ? _GEN3958 : _GEN3741;
wire  _GEN3960 = io_x[16] ? _GEN3959 : _GEN3955;
wire  _GEN3961 = io_x[12] ? _GEN3960 : _GEN3946;
wire  _GEN3962 = io_x[2] ? _GEN3961 : _GEN3936;
wire  _GEN3963 = io_x[23] ? _GEN3713 : _GEN3741;
wire  _GEN3964 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3965 = io_x[14] ? _GEN3708 : _GEN3964;
wire  _GEN3966 = io_x[10] ? _GEN3711 : _GEN3965;
wire  _GEN3967 = io_x[23] ? _GEN3713 : _GEN3966;
wire  _GEN3968 = io_x[16] ? _GEN3967 : _GEN3963;
wire  _GEN3969 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN3970 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN3971 = io_x[10] ? _GEN3970 : _GEN3969;
wire  _GEN3972 = io_x[23] ? _GEN3741 : _GEN3971;
wire  _GEN3973 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3974 = io_x[14] ? _GEN3973 : _GEN3708;
wire  _GEN3975 = io_x[10] ? _GEN3974 : _GEN3711;
wire  _GEN3976 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN3977 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN3978 = io_x[10] ? _GEN3977 : _GEN3976;
wire  _GEN3979 = io_x[23] ? _GEN3978 : _GEN3975;
wire  _GEN3980 = io_x[16] ? _GEN3979 : _GEN3972;
wire  _GEN3981 = io_x[12] ? _GEN3980 : _GEN3968;
wire  _GEN3982 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3983 = io_x[14] ? _GEN3982 : _GEN3709;
wire  _GEN3984 = io_x[10] ? _GEN3716 : _GEN3983;
wire  _GEN3985 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3986 = io_x[14] ? _GEN3709 : _GEN3985;
wire  _GEN3987 = io_x[10] ? _GEN3711 : _GEN3986;
wire  _GEN3988 = io_x[23] ? _GEN3987 : _GEN3984;
wire  _GEN3989 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3990 = io_x[14] ? _GEN3709 : _GEN3989;
wire  _GEN3991 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN3992 = io_x[14] ? _GEN3708 : _GEN3991;
wire  _GEN3993 = io_x[10] ? _GEN3992 : _GEN3990;
wire  _GEN3994 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN3995 = io_x[23] ? _GEN3994 : _GEN3993;
wire  _GEN3996 = io_x[16] ? _GEN3995 : _GEN3988;
wire  _GEN3997 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN3998 = io_x[14] ? _GEN3997 : _GEN3709;
wire  _GEN3999 = io_x[10] ? _GEN3998 : _GEN3711;
wire  _GEN4000 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4001 = io_x[14] ? _GEN4000 : _GEN3709;
wire  _GEN4002 = io_x[10] ? _GEN4001 : _GEN3711;
wire  _GEN4003 = io_x[23] ? _GEN4002 : _GEN3999;
wire  _GEN4004 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4005 = io_x[14] ? _GEN4004 : _GEN3709;
wire  _GEN4006 = io_x[10] ? _GEN4005 : _GEN3711;
wire  _GEN4007 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4008 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4009 = io_x[14] ? _GEN4008 : _GEN3709;
wire  _GEN4010 = io_x[10] ? _GEN4009 : _GEN4007;
wire  _GEN4011 = io_x[23] ? _GEN4010 : _GEN4006;
wire  _GEN4012 = io_x[16] ? _GEN4011 : _GEN4003;
wire  _GEN4013 = io_x[12] ? _GEN4012 : _GEN3996;
wire  _GEN4014 = io_x[2] ? _GEN4013 : _GEN3981;
wire  _GEN4015 = io_x[9] ? _GEN4014 : _GEN3962;
wire  _GEN4016 = io_x[13] ? _GEN4015 : _GEN3920;
wire  _GEN4017 = io_x[7] ? _GEN4016 : _GEN3862;
wire  _GEN4018 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4019 = io_x[10] ? _GEN4018 : _GEN3716;
wire  _GEN4020 = io_x[23] ? _GEN4019 : _GEN3741;
wire  _GEN4021 = io_x[16] ? _GEN4020 : _GEN3727;
wire  _GEN4022 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN4023 = io_x[23] ? _GEN3713 : _GEN4022;
wire  _GEN4024 = io_x[16] ? _GEN3727 : _GEN4023;
wire  _GEN4025 = io_x[12] ? _GEN4024 : _GEN4021;
wire  _GEN4026 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4027 = io_x[10] ? _GEN4026 : _GEN3716;
wire  _GEN4028 = io_x[23] ? _GEN3741 : _GEN4027;
wire  _GEN4029 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN4030 = io_x[23] ? _GEN4029 : _GEN3713;
wire  _GEN4031 = io_x[16] ? _GEN4030 : _GEN4028;
wire  _GEN4032 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4033 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4034 = io_x[14] ? _GEN4033 : _GEN3709;
wire  _GEN4035 = io_x[10] ? _GEN4034 : _GEN4032;
wire  _GEN4036 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4037 = io_x[10] ? _GEN4036 : _GEN3716;
wire  _GEN4038 = io_x[23] ? _GEN4037 : _GEN4035;
wire  _GEN4039 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4040 = io_x[14] ? _GEN4039 : _GEN3709;
wire  _GEN4041 = io_x[10] ? _GEN4040 : _GEN3711;
wire  _GEN4042 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4043 = io_x[10] ? _GEN3716 : _GEN4042;
wire  _GEN4044 = io_x[23] ? _GEN4043 : _GEN4041;
wire  _GEN4045 = io_x[16] ? _GEN4044 : _GEN4038;
wire  _GEN4046 = io_x[12] ? _GEN4045 : _GEN4031;
wire  _GEN4047 = io_x[2] ? _GEN4046 : _GEN4025;
wire  _GEN4048 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4049 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4050 = io_x[14] ? _GEN4049 : _GEN4048;
wire  _GEN4051 = io_x[10] ? _GEN4050 : _GEN3711;
wire  _GEN4052 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN4053 = io_x[23] ? _GEN4052 : _GEN4051;
wire  _GEN4054 = io_x[16] ? _GEN4053 : _GEN3707;
wire  _GEN4055 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4056 = io_x[14] ? _GEN3709 : _GEN4055;
wire  _GEN4057 = io_x[10] ? _GEN3716 : _GEN4056;
wire  _GEN4058 = io_x[23] ? _GEN3713 : _GEN4057;
wire  _GEN4059 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4060 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4061 = io_x[10] ? _GEN4060 : _GEN4059;
wire  _GEN4062 = io_x[23] ? _GEN3713 : _GEN4061;
wire  _GEN4063 = io_x[16] ? _GEN4062 : _GEN4058;
wire  _GEN4064 = io_x[12] ? _GEN4063 : _GEN4054;
wire  _GEN4065 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN4066 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4067 = io_x[10] ? _GEN3711 : _GEN4066;
wire  _GEN4068 = io_x[23] ? _GEN4067 : _GEN4065;
wire  _GEN4069 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4070 = io_x[14] ? _GEN4069 : _GEN3709;
wire  _GEN4071 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4072 = io_x[14] ? _GEN4071 : _GEN3708;
wire  _GEN4073 = io_x[10] ? _GEN4072 : _GEN4070;
wire  _GEN4074 = io_x[23] ? _GEN4073 : _GEN3713;
wire  _GEN4075 = io_x[16] ? _GEN4074 : _GEN4068;
wire  _GEN4076 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4077 = io_x[10] ? _GEN4076 : _GEN3711;
wire  _GEN4078 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4079 = io_x[10] ? _GEN3711 : _GEN4078;
wire  _GEN4080 = io_x[23] ? _GEN4079 : _GEN4077;
wire  _GEN4081 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4082 = io_x[14] ? _GEN4081 : _GEN3709;
wire  _GEN4083 = io_x[10] ? _GEN4082 : _GEN3711;
wire  _GEN4084 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4085 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4086 = io_x[10] ? _GEN4085 : _GEN4084;
wire  _GEN4087 = io_x[23] ? _GEN4086 : _GEN4083;
wire  _GEN4088 = io_x[16] ? _GEN4087 : _GEN4080;
wire  _GEN4089 = io_x[12] ? _GEN4088 : _GEN4075;
wire  _GEN4090 = io_x[2] ? _GEN4089 : _GEN4064;
wire  _GEN4091 = io_x[9] ? _GEN4090 : _GEN4047;
wire  _GEN4092 = io_x[23] ? _GEN3713 : _GEN3741;
wire  _GEN4093 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4094 = io_x[10] ? _GEN3711 : _GEN4093;
wire  _GEN4095 = io_x[23] ? _GEN4094 : _GEN3741;
wire  _GEN4096 = io_x[16] ? _GEN4095 : _GEN4092;
wire  _GEN4097 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4098 = io_x[14] ? _GEN4097 : _GEN3709;
wire  _GEN4099 = io_x[10] ? _GEN4098 : _GEN3711;
wire  _GEN4100 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4101 = io_x[10] ? _GEN4100 : _GEN3711;
wire  _GEN4102 = io_x[23] ? _GEN4101 : _GEN4099;
wire  _GEN4103 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN4104 = io_x[23] ? _GEN4103 : _GEN3741;
wire  _GEN4105 = io_x[16] ? _GEN4104 : _GEN4102;
wire  _GEN4106 = io_x[12] ? _GEN4105 : _GEN4096;
wire  _GEN4107 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4108 = io_x[14] ? _GEN4107 : _GEN3709;
wire  _GEN4109 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4110 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4111 = io_x[14] ? _GEN4110 : _GEN4109;
wire  _GEN4112 = io_x[10] ? _GEN4111 : _GEN4108;
wire  _GEN4113 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4114 = io_x[10] ? _GEN4113 : _GEN3711;
wire  _GEN4115 = io_x[23] ? _GEN4114 : _GEN4112;
wire  _GEN4116 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4117 = io_x[10] ? _GEN3711 : _GEN4116;
wire  _GEN4118 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4119 = io_x[10] ? _GEN4118 : _GEN3716;
wire  _GEN4120 = io_x[23] ? _GEN4119 : _GEN4117;
wire  _GEN4121 = io_x[16] ? _GEN4120 : _GEN4115;
wire  _GEN4122 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4123 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4124 = io_x[14] ? _GEN4123 : _GEN4122;
wire  _GEN4125 = io_x[10] ? _GEN4124 : _GEN3711;
wire  _GEN4126 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4127 = io_x[10] ? _GEN4126 : _GEN3711;
wire  _GEN4128 = io_x[23] ? _GEN4127 : _GEN4125;
wire  _GEN4129 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4130 = io_x[14] ? _GEN4129 : _GEN3709;
wire  _GEN4131 = io_x[10] ? _GEN4130 : _GEN3716;
wire  _GEN4132 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4133 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4134 = io_x[14] ? _GEN4133 : _GEN3709;
wire  _GEN4135 = io_x[10] ? _GEN4134 : _GEN4132;
wire  _GEN4136 = io_x[23] ? _GEN4135 : _GEN4131;
wire  _GEN4137 = io_x[16] ? _GEN4136 : _GEN4128;
wire  _GEN4138 = io_x[12] ? _GEN4137 : _GEN4121;
wire  _GEN4139 = io_x[2] ? _GEN4138 : _GEN4106;
wire  _GEN4140 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4141 = io_x[14] ? _GEN4140 : _GEN3709;
wire  _GEN4142 = io_x[10] ? _GEN4141 : _GEN3711;
wire  _GEN4143 = io_x[23] ? _GEN3741 : _GEN4142;
wire  _GEN4144 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4145 = io_x[14] ? _GEN4144 : _GEN3709;
wire  _GEN4146 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4147 = io_x[14] ? _GEN4146 : _GEN4048;
wire  _GEN4148 = io_x[10] ? _GEN4147 : _GEN4145;
wire  _GEN4149 = io_x[23] ? _GEN3741 : _GEN4148;
wire  _GEN4150 = io_x[16] ? _GEN4149 : _GEN4143;
wire  _GEN4151 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4152 = io_x[14] ? _GEN4151 : _GEN3709;
wire  _GEN4153 = io_x[10] ? _GEN4152 : _GEN3711;
wire  _GEN4154 = io_x[23] ? _GEN3741 : _GEN4153;
wire  _GEN4155 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4156 = io_x[14] ? _GEN4155 : _GEN3709;
wire  _GEN4157 = io_x[10] ? _GEN4156 : _GEN3711;
wire  _GEN4158 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4159 = io_x[14] ? _GEN4158 : _GEN3709;
wire  _GEN4160 = io_x[10] ? _GEN4159 : _GEN3711;
wire  _GEN4161 = io_x[23] ? _GEN4160 : _GEN4157;
wire  _GEN4162 = io_x[16] ? _GEN4161 : _GEN4154;
wire  _GEN4163 = io_x[12] ? _GEN4162 : _GEN4150;
wire  _GEN4164 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4165 = io_x[14] ? _GEN4164 : _GEN3709;
wire  _GEN4166 = io_x[10] ? _GEN4165 : _GEN3716;
wire  _GEN4167 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4168 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4169 = io_x[10] ? _GEN4168 : _GEN4167;
wire  _GEN4170 = io_x[23] ? _GEN4169 : _GEN4166;
wire  _GEN4171 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4172 = io_x[14] ? _GEN3709 : _GEN4171;
wire  _GEN4173 = io_x[10] ? _GEN3711 : _GEN4172;
wire  _GEN4174 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4175 = io_x[14] ? _GEN3708 : _GEN4174;
wire  _GEN4176 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4177 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4178 = io_x[14] ? _GEN4177 : _GEN4176;
wire  _GEN4179 = io_x[10] ? _GEN4178 : _GEN4175;
wire  _GEN4180 = io_x[23] ? _GEN4179 : _GEN4173;
wire  _GEN4181 = io_x[16] ? _GEN4180 : _GEN4170;
wire  _GEN4182 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4183 = io_x[14] ? _GEN4182 : _GEN3709;
wire  _GEN4184 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4185 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4186 = io_x[14] ? _GEN4185 : _GEN4184;
wire  _GEN4187 = io_x[10] ? _GEN4186 : _GEN4183;
wire  _GEN4188 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4189 = io_x[14] ? _GEN4188 : _GEN3709;
wire  _GEN4190 = io_x[10] ? _GEN4189 : _GEN3716;
wire  _GEN4191 = io_x[23] ? _GEN4190 : _GEN4187;
wire  _GEN4192 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4193 = io_x[10] ? _GEN4192 : _GEN3716;
wire  _GEN4194 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4195 = io_x[14] ? _GEN4194 : _GEN3709;
wire  _GEN4196 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4197 = io_x[14] ? _GEN4196 : _GEN3709;
wire  _GEN4198 = io_x[10] ? _GEN4197 : _GEN4195;
wire  _GEN4199 = io_x[23] ? _GEN4198 : _GEN4193;
wire  _GEN4200 = io_x[16] ? _GEN4199 : _GEN4191;
wire  _GEN4201 = io_x[12] ? _GEN4200 : _GEN4181;
wire  _GEN4202 = io_x[2] ? _GEN4201 : _GEN4163;
wire  _GEN4203 = io_x[9] ? _GEN4202 : _GEN4139;
wire  _GEN4204 = io_x[13] ? _GEN4203 : _GEN4091;
wire  _GEN4205 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4206 = io_x[10] ? _GEN4205 : _GEN3711;
wire  _GEN4207 = io_x[23] ? _GEN3713 : _GEN4206;
wire  _GEN4208 = io_x[16] ? _GEN4207 : _GEN3707;
wire  _GEN4209 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4210 = io_x[14] ? _GEN4209 : _GEN3708;
wire  _GEN4211 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4212 = io_x[14] ? _GEN3709 : _GEN4211;
wire  _GEN4213 = io_x[10] ? _GEN4212 : _GEN4210;
wire  _GEN4214 = io_x[23] ? _GEN3713 : _GEN4213;
wire  _GEN4215 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4216 = io_x[14] ? _GEN3709 : _GEN4215;
wire  _GEN4217 = io_x[10] ? _GEN4216 : _GEN3716;
wire  _GEN4218 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN4219 = io_x[23] ? _GEN4218 : _GEN4217;
wire  _GEN4220 = io_x[16] ? _GEN4219 : _GEN4214;
wire  _GEN4221 = io_x[12] ? _GEN4220 : _GEN4208;
wire  _GEN4222 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4223 = io_x[14] ? _GEN4222 : _GEN3709;
wire  _GEN4224 = io_x[10] ? _GEN4223 : _GEN3711;
wire  _GEN4225 = io_x[23] ? _GEN4224 : _GEN3713;
wire  _GEN4226 = io_x[16] ? _GEN4225 : _GEN3727;
wire  _GEN4227 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4228 = io_x[14] ? _GEN4227 : _GEN3708;
wire  _GEN4229 = io_x[10] ? _GEN4228 : _GEN3711;
wire  _GEN4230 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4231 = io_x[14] ? _GEN3709 : _GEN4230;
wire  _GEN4232 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4233 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4234 = io_x[14] ? _GEN4233 : _GEN4232;
wire  _GEN4235 = io_x[10] ? _GEN4234 : _GEN4231;
wire  _GEN4236 = io_x[23] ? _GEN4235 : _GEN4229;
wire  _GEN4237 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4238 = io_x[14] ? _GEN4237 : _GEN3709;
wire  _GEN4239 = io_x[10] ? _GEN4238 : _GEN3711;
wire  _GEN4240 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4241 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4242 = io_x[14] ? _GEN4241 : _GEN4240;
wire  _GEN4243 = io_x[10] ? _GEN4242 : _GEN3716;
wire  _GEN4244 = io_x[23] ? _GEN4243 : _GEN4239;
wire  _GEN4245 = io_x[16] ? _GEN4244 : _GEN4236;
wire  _GEN4246 = io_x[12] ? _GEN4245 : _GEN4226;
wire  _GEN4247 = io_x[2] ? _GEN4246 : _GEN4221;
wire  _GEN4248 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4249 = io_x[10] ? _GEN4248 : _GEN3711;
wire  _GEN4250 = io_x[23] ? _GEN3713 : _GEN4249;
wire  _GEN4251 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4252 = io_x[14] ? _GEN3709 : _GEN4251;
wire  _GEN4253 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4254 = io_x[10] ? _GEN4253 : _GEN4252;
wire  _GEN4255 = io_x[23] ? _GEN3713 : _GEN4254;
wire  _GEN4256 = io_x[16] ? _GEN4255 : _GEN4250;
wire  _GEN4257 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4258 = io_x[14] ? _GEN4257 : _GEN3709;
wire  _GEN4259 = io_x[10] ? _GEN4258 : _GEN3716;
wire  _GEN4260 = io_x[23] ? _GEN3713 : _GEN4259;
wire  _GEN4261 = io_x[16] ? _GEN3707 : _GEN4260;
wire  _GEN4262 = io_x[12] ? _GEN4261 : _GEN4256;
wire  _GEN4263 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4264 = io_x[14] ? _GEN4263 : _GEN3709;
wire  _GEN4265 = io_x[10] ? _GEN4264 : _GEN3711;
wire  _GEN4266 = io_x[23] ? _GEN4265 : _GEN3741;
wire  _GEN4267 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN4268 = io_x[23] ? _GEN3741 : _GEN4267;
wire  _GEN4269 = io_x[16] ? _GEN4268 : _GEN4266;
wire  _GEN4270 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4271 = io_x[14] ? _GEN4270 : _GEN3709;
wire  _GEN4272 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4273 = io_x[14] ? _GEN4272 : _GEN3709;
wire  _GEN4274 = io_x[10] ? _GEN4273 : _GEN4271;
wire  _GEN4275 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4276 = io_x[14] ? _GEN4275 : _GEN3709;
wire  _GEN4277 = io_x[10] ? _GEN4276 : _GEN3711;
wire  _GEN4278 = io_x[23] ? _GEN4277 : _GEN4274;
wire  _GEN4279 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4280 = io_x[14] ? _GEN4279 : _GEN3709;
wire  _GEN4281 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4282 = io_x[10] ? _GEN4281 : _GEN4280;
wire  _GEN4283 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4284 = io_x[14] ? _GEN4283 : _GEN3708;
wire  _GEN4285 = io_x[10] ? _GEN4284 : _GEN3711;
wire  _GEN4286 = io_x[23] ? _GEN4285 : _GEN4282;
wire  _GEN4287 = io_x[16] ? _GEN4286 : _GEN4278;
wire  _GEN4288 = io_x[12] ? _GEN4287 : _GEN4269;
wire  _GEN4289 = io_x[2] ? _GEN4288 : _GEN4262;
wire  _GEN4290 = io_x[9] ? _GEN4289 : _GEN4247;
wire  _GEN4291 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4292 = io_x[14] ? _GEN4291 : _GEN3709;
wire  _GEN4293 = io_x[10] ? _GEN3716 : _GEN4292;
wire  _GEN4294 = io_x[23] ? _GEN3713 : _GEN4293;
wire  _GEN4295 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4296 = io_x[10] ? _GEN3711 : _GEN4295;
wire  _GEN4297 = io_x[23] ? _GEN4296 : _GEN3741;
wire  _GEN4298 = io_x[16] ? _GEN4297 : _GEN4294;
wire  _GEN4299 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4300 = io_x[14] ? _GEN4299 : _GEN3709;
wire  _GEN4301 = io_x[10] ? _GEN3711 : _GEN4300;
wire  _GEN4302 = io_x[23] ? _GEN3713 : _GEN4301;
wire  _GEN4303 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4304 = io_x[14] ? _GEN4303 : _GEN3709;
wire  _GEN4305 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4306 = io_x[14] ? _GEN4305 : _GEN3708;
wire  _GEN4307 = io_x[10] ? _GEN4306 : _GEN4304;
wire  _GEN4308 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN4309 = io_x[23] ? _GEN4308 : _GEN4307;
wire  _GEN4310 = io_x[16] ? _GEN4309 : _GEN4302;
wire  _GEN4311 = io_x[12] ? _GEN4310 : _GEN4298;
wire  _GEN4312 = io_x[23] ? _GEN3713 : _GEN3741;
wire  _GEN4313 = io_x[16] ? _GEN4312 : _GEN3707;
wire  _GEN4314 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4315 = io_x[14] ? _GEN3708 : _GEN4314;
wire  _GEN4316 = io_x[10] ? _GEN4315 : _GEN3711;
wire  _GEN4317 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4318 = io_x[10] ? _GEN4317 : _GEN3711;
wire  _GEN4319 = io_x[23] ? _GEN4318 : _GEN4316;
wire  _GEN4320 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4321 = io_x[14] ? _GEN3708 : _GEN4320;
wire  _GEN4322 = io_x[10] ? _GEN4321 : _GEN3711;
wire  _GEN4323 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4324 = io_x[10] ? _GEN4323 : _GEN3711;
wire  _GEN4325 = io_x[23] ? _GEN4324 : _GEN4322;
wire  _GEN4326 = io_x[16] ? _GEN4325 : _GEN4319;
wire  _GEN4327 = io_x[12] ? _GEN4326 : _GEN4313;
wire  _GEN4328 = io_x[2] ? _GEN4327 : _GEN4311;
wire  _GEN4329 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4330 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4331 = io_x[14] ? _GEN4330 : _GEN4329;
wire  _GEN4332 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4333 = io_x[10] ? _GEN4332 : _GEN4331;
wire  _GEN4334 = io_x[23] ? _GEN3713 : _GEN4333;
wire  _GEN4335 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4336 = io_x[14] ? _GEN3709 : _GEN4335;
wire  _GEN4337 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4338 = io_x[10] ? _GEN4337 : _GEN4336;
wire  _GEN4339 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN4340 = io_x[23] ? _GEN4339 : _GEN4338;
wire  _GEN4341 = io_x[16] ? _GEN4340 : _GEN4334;
wire  _GEN4342 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4343 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4344 = io_x[14] ? _GEN4343 : _GEN4342;
wire  _GEN4345 = io_x[10] ? _GEN4344 : _GEN3711;
wire  _GEN4346 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4347 = io_x[14] ? _GEN4346 : _GEN3709;
wire  _GEN4348 = io_x[10] ? _GEN4347 : _GEN3711;
wire  _GEN4349 = io_x[23] ? _GEN4348 : _GEN4345;
wire  _GEN4350 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4351 = io_x[14] ? _GEN4350 : _GEN3708;
wire  _GEN4352 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4353 = io_x[14] ? _GEN4352 : _GEN3708;
wire  _GEN4354 = io_x[10] ? _GEN4353 : _GEN4351;
wire  _GEN4355 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4356 = io_x[14] ? _GEN4355 : _GEN3708;
wire  _GEN4357 = io_x[10] ? _GEN4356 : _GEN3716;
wire  _GEN4358 = io_x[23] ? _GEN4357 : _GEN4354;
wire  _GEN4359 = io_x[16] ? _GEN4358 : _GEN4349;
wire  _GEN4360 = io_x[12] ? _GEN4359 : _GEN4341;
wire  _GEN4361 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4362 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4363 = io_x[14] ? _GEN4362 : _GEN4361;
wire  _GEN4364 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4365 = io_x[14] ? _GEN3708 : _GEN4364;
wire  _GEN4366 = io_x[10] ? _GEN4365 : _GEN4363;
wire  _GEN4367 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4368 = io_x[14] ? _GEN3709 : _GEN4367;
wire  _GEN4369 = io_x[10] ? _GEN3716 : _GEN4368;
wire  _GEN4370 = io_x[23] ? _GEN4369 : _GEN4366;
wire  _GEN4371 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4372 = io_x[14] ? _GEN4371 : _GEN3709;
wire  _GEN4373 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4374 = io_x[14] ? _GEN4373 : _GEN3709;
wire  _GEN4375 = io_x[10] ? _GEN4374 : _GEN4372;
wire  _GEN4376 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4377 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4378 = io_x[14] ? _GEN4377 : _GEN4376;
wire  _GEN4379 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4380 = io_x[14] ? _GEN3708 : _GEN4379;
wire  _GEN4381 = io_x[10] ? _GEN4380 : _GEN4378;
wire  _GEN4382 = io_x[23] ? _GEN4381 : _GEN4375;
wire  _GEN4383 = io_x[16] ? _GEN4382 : _GEN4370;
wire  _GEN4384 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4385 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4386 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4387 = io_x[14] ? _GEN4386 : _GEN4385;
wire  _GEN4388 = io_x[10] ? _GEN4387 : _GEN4384;
wire  _GEN4389 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4390 = io_x[10] ? _GEN4389 : _GEN3711;
wire  _GEN4391 = io_x[23] ? _GEN4390 : _GEN4388;
wire  _GEN4392 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4393 = io_x[14] ? _GEN4392 : _GEN3709;
wire  _GEN4394 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4395 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4396 = io_x[14] ? _GEN4395 : _GEN4394;
wire  _GEN4397 = io_x[10] ? _GEN4396 : _GEN4393;
wire  _GEN4398 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4399 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4400 = io_x[14] ? _GEN4399 : _GEN4398;
wire  _GEN4401 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4402 = io_x[14] ? _GEN4401 : _GEN3709;
wire  _GEN4403 = io_x[10] ? _GEN4402 : _GEN4400;
wire  _GEN4404 = io_x[23] ? _GEN4403 : _GEN4397;
wire  _GEN4405 = io_x[16] ? _GEN4404 : _GEN4391;
wire  _GEN4406 = io_x[12] ? _GEN4405 : _GEN4383;
wire  _GEN4407 = io_x[2] ? _GEN4406 : _GEN4360;
wire  _GEN4408 = io_x[9] ? _GEN4407 : _GEN4328;
wire  _GEN4409 = io_x[13] ? _GEN4408 : _GEN4290;
wire  _GEN4410 = io_x[7] ? _GEN4409 : _GEN4204;
wire  _GEN4411 = io_x[15] ? _GEN4410 : _GEN4017;
wire  _GEN4412 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4413 = io_x[14] ? _GEN4412 : _GEN3709;
wire  _GEN4414 = io_x[10] ? _GEN4413 : _GEN3711;
wire  _GEN4415 = io_x[23] ? _GEN3713 : _GEN4414;
wire  _GEN4416 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4417 = io_x[14] ? _GEN4416 : _GEN3709;
wire  _GEN4418 = io_x[10] ? _GEN4417 : _GEN3711;
wire  _GEN4419 = io_x[23] ? _GEN3713 : _GEN4418;
wire  _GEN4420 = io_x[16] ? _GEN4419 : _GEN4415;
wire  _GEN4421 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4422 = io_x[14] ? _GEN3709 : _GEN4421;
wire  _GEN4423 = io_x[10] ? _GEN4422 : _GEN3711;
wire  _GEN4424 = io_x[23] ? _GEN3741 : _GEN4423;
wire  _GEN4425 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4426 = io_x[10] ? _GEN4425 : _GEN3711;
wire  _GEN4427 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4428 = io_x[14] ? _GEN4427 : _GEN3709;
wire  _GEN4429 = io_x[10] ? _GEN4428 : _GEN3711;
wire  _GEN4430 = io_x[23] ? _GEN4429 : _GEN4426;
wire  _GEN4431 = io_x[16] ? _GEN4430 : _GEN4424;
wire  _GEN4432 = io_x[12] ? _GEN4431 : _GEN4420;
wire  _GEN4433 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN4434 = io_x[23] ? _GEN4433 : _GEN3741;
wire  _GEN4435 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4436 = io_x[14] ? _GEN4435 : _GEN3709;
wire  _GEN4437 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4438 = io_x[14] ? _GEN4437 : _GEN3709;
wire  _GEN4439 = io_x[10] ? _GEN4438 : _GEN4436;
wire  _GEN4440 = io_x[23] ? _GEN4439 : _GEN3713;
wire  _GEN4441 = io_x[16] ? _GEN4440 : _GEN4434;
wire  _GEN4442 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN4443 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN4444 = io_x[23] ? _GEN4443 : _GEN4442;
wire  _GEN4445 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4446 = io_x[14] ? _GEN4445 : _GEN3709;
wire  _GEN4447 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4448 = io_x[14] ? _GEN4447 : _GEN3709;
wire  _GEN4449 = io_x[10] ? _GEN4448 : _GEN4446;
wire  _GEN4450 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4451 = io_x[14] ? _GEN4450 : _GEN3709;
wire  _GEN4452 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4453 = io_x[14] ? _GEN4452 : _GEN3709;
wire  _GEN4454 = io_x[10] ? _GEN4453 : _GEN4451;
wire  _GEN4455 = io_x[23] ? _GEN4454 : _GEN4449;
wire  _GEN4456 = io_x[16] ? _GEN4455 : _GEN4444;
wire  _GEN4457 = io_x[12] ? _GEN4456 : _GEN4441;
wire  _GEN4458 = io_x[2] ? _GEN4457 : _GEN4432;
wire  _GEN4459 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN4460 = io_x[23] ? _GEN4459 : _GEN3713;
wire  _GEN4461 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4462 = io_x[10] ? _GEN4461 : _GEN3711;
wire  _GEN4463 = io_x[23] ? _GEN3713 : _GEN4462;
wire  _GEN4464 = io_x[16] ? _GEN4463 : _GEN4460;
wire  _GEN4465 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4466 = io_x[14] ? _GEN4465 : _GEN3709;
wire  _GEN4467 = io_x[10] ? _GEN3716 : _GEN4466;
wire  _GEN4468 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4469 = io_x[14] ? _GEN4468 : _GEN3709;
wire  _GEN4470 = io_x[10] ? _GEN3711 : _GEN4469;
wire  _GEN4471 = io_x[23] ? _GEN4470 : _GEN4467;
wire  _GEN4472 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4473 = io_x[14] ? _GEN4472 : _GEN3708;
wire  _GEN4474 = io_x[10] ? _GEN4473 : _GEN3716;
wire  _GEN4475 = io_x[23] ? _GEN3713 : _GEN4474;
wire  _GEN4476 = io_x[16] ? _GEN4475 : _GEN4471;
wire  _GEN4477 = io_x[12] ? _GEN4476 : _GEN4464;
wire  _GEN4478 = 1'b0;
wire  _GEN4479 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4480 = io_x[14] ? _GEN4479 : _GEN3709;
wire  _GEN4481 = io_x[10] ? _GEN4480 : _GEN3716;
wire  _GEN4482 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4483 = io_x[10] ? _GEN4482 : _GEN3711;
wire  _GEN4484 = io_x[23] ? _GEN4483 : _GEN4481;
wire  _GEN4485 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4486 = io_x[14] ? _GEN4485 : _GEN3709;
wire  _GEN4487 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4488 = io_x[14] ? _GEN4487 : _GEN3709;
wire  _GEN4489 = io_x[10] ? _GEN4488 : _GEN4486;
wire  _GEN4490 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4491 = io_x[10] ? _GEN3711 : _GEN4490;
wire  _GEN4492 = io_x[23] ? _GEN4491 : _GEN4489;
wire  _GEN4493 = io_x[16] ? _GEN4492 : _GEN4484;
wire  _GEN4494 = io_x[12] ? _GEN4493 : _GEN4478;
wire  _GEN4495 = io_x[2] ? _GEN4494 : _GEN4477;
wire  _GEN4496 = io_x[9] ? _GEN4495 : _GEN4458;
wire  _GEN4497 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4498 = io_x[10] ? _GEN4497 : _GEN3711;
wire  _GEN4499 = io_x[23] ? _GEN3713 : _GEN4498;
wire  _GEN4500 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN4501 = io_x[23] ? _GEN4500 : _GEN3713;
wire  _GEN4502 = io_x[16] ? _GEN4501 : _GEN4499;
wire  _GEN4503 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN4504 = io_x[23] ? _GEN4503 : _GEN3713;
wire  _GEN4505 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4506 = io_x[14] ? _GEN4505 : _GEN3709;
wire  _GEN4507 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4508 = io_x[10] ? _GEN4507 : _GEN4506;
wire  _GEN4509 = io_x[23] ? _GEN3713 : _GEN4508;
wire  _GEN4510 = io_x[16] ? _GEN4509 : _GEN4504;
wire  _GEN4511 = io_x[12] ? _GEN4510 : _GEN4502;
wire  _GEN4512 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4513 = io_x[10] ? _GEN4512 : _GEN3711;
wire  _GEN4514 = io_x[23] ? _GEN4513 : _GEN3741;
wire  _GEN4515 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4516 = io_x[14] ? _GEN4515 : _GEN3709;
wire  _GEN4517 = io_x[10] ? _GEN4516 : _GEN3716;
wire  _GEN4518 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4519 = io_x[14] ? _GEN3709 : _GEN4518;
wire  _GEN4520 = io_x[10] ? _GEN4519 : _GEN3711;
wire  _GEN4521 = io_x[23] ? _GEN4520 : _GEN4517;
wire  _GEN4522 = io_x[16] ? _GEN4521 : _GEN4514;
wire  _GEN4523 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4524 = io_x[10] ? _GEN4523 : _GEN3711;
wire  _GEN4525 = io_x[23] ? _GEN4524 : _GEN3741;
wire  _GEN4526 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4527 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4528 = io_x[10] ? _GEN4527 : _GEN4526;
wire  _GEN4529 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4530 = io_x[10] ? _GEN4529 : _GEN3711;
wire  _GEN4531 = io_x[23] ? _GEN4530 : _GEN4528;
wire  _GEN4532 = io_x[16] ? _GEN4531 : _GEN4525;
wire  _GEN4533 = io_x[12] ? _GEN4532 : _GEN4522;
wire  _GEN4534 = io_x[2] ? _GEN4533 : _GEN4511;
wire  _GEN4535 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4536 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4537 = io_x[10] ? _GEN4536 : _GEN4535;
wire  _GEN4538 = io_x[23] ? _GEN4537 : _GEN3741;
wire  _GEN4539 = io_x[16] ? _GEN4538 : _GEN3727;
wire  _GEN4540 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN4541 = io_x[23] ? _GEN4540 : _GEN3713;
wire  _GEN4542 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4543 = io_x[10] ? _GEN4542 : _GEN3711;
wire  _GEN4544 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4545 = io_x[14] ? _GEN3708 : _GEN4544;
wire  _GEN4546 = io_x[10] ? _GEN4545 : _GEN3711;
wire  _GEN4547 = io_x[23] ? _GEN4546 : _GEN4543;
wire  _GEN4548 = io_x[16] ? _GEN4547 : _GEN4541;
wire  _GEN4549 = io_x[12] ? _GEN4548 : _GEN4539;
wire  _GEN4550 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4551 = io_x[10] ? _GEN4550 : _GEN3711;
wire  _GEN4552 = io_x[23] ? _GEN4551 : _GEN3713;
wire  _GEN4553 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4554 = io_x[10] ? _GEN3711 : _GEN4553;
wire  _GEN4555 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4556 = io_x[10] ? _GEN3711 : _GEN4555;
wire  _GEN4557 = io_x[23] ? _GEN4556 : _GEN4554;
wire  _GEN4558 = io_x[16] ? _GEN4557 : _GEN4552;
wire  _GEN4559 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4560 = io_x[14] ? _GEN4559 : _GEN3709;
wire  _GEN4561 = io_x[10] ? _GEN4560 : _GEN3711;
wire  _GEN4562 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4563 = io_x[10] ? _GEN4562 : _GEN3711;
wire  _GEN4564 = io_x[23] ? _GEN4563 : _GEN4561;
wire  _GEN4565 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4566 = io_x[14] ? _GEN4565 : _GEN3709;
wire  _GEN4567 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4568 = io_x[14] ? _GEN4567 : _GEN3708;
wire  _GEN4569 = io_x[10] ? _GEN4568 : _GEN4566;
wire  _GEN4570 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4571 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4572 = io_x[14] ? _GEN4571 : _GEN4570;
wire  _GEN4573 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4574 = io_x[14] ? _GEN4573 : _GEN3709;
wire  _GEN4575 = io_x[10] ? _GEN4574 : _GEN4572;
wire  _GEN4576 = io_x[23] ? _GEN4575 : _GEN4569;
wire  _GEN4577 = io_x[16] ? _GEN4576 : _GEN4564;
wire  _GEN4578 = io_x[12] ? _GEN4577 : _GEN4558;
wire  _GEN4579 = io_x[2] ? _GEN4578 : _GEN4549;
wire  _GEN4580 = io_x[9] ? _GEN4579 : _GEN4534;
wire  _GEN4581 = io_x[13] ? _GEN4580 : _GEN4496;
wire  _GEN4582 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4583 = io_x[10] ? _GEN4582 : _GEN3711;
wire  _GEN4584 = io_x[23] ? _GEN4583 : _GEN3713;
wire  _GEN4585 = io_x[16] ? _GEN4584 : _GEN3707;
wire  _GEN4586 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN4587 = io_x[23] ? _GEN3713 : _GEN4586;
wire  _GEN4588 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4589 = io_x[14] ? _GEN4588 : _GEN3709;
wire  _GEN4590 = io_x[10] ? _GEN4589 : _GEN3711;
wire  _GEN4591 = io_x[23] ? _GEN3741 : _GEN4590;
wire  _GEN4592 = io_x[16] ? _GEN4591 : _GEN4587;
wire  _GEN4593 = io_x[12] ? _GEN4592 : _GEN4585;
wire  _GEN4594 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4595 = io_x[14] ? _GEN4594 : _GEN3709;
wire  _GEN4596 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4597 = io_x[14] ? _GEN4596 : _GEN3709;
wire  _GEN4598 = io_x[10] ? _GEN4597 : _GEN4595;
wire  _GEN4599 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4600 = io_x[14] ? _GEN4599 : _GEN3709;
wire  _GEN4601 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4602 = io_x[14] ? _GEN4601 : _GEN3709;
wire  _GEN4603 = io_x[10] ? _GEN4602 : _GEN4600;
wire  _GEN4604 = io_x[23] ? _GEN4603 : _GEN4598;
wire  _GEN4605 = io_x[16] ? _GEN4604 : _GEN3727;
wire  _GEN4606 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4607 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4608 = io_x[14] ? _GEN4607 : _GEN3708;
wire  _GEN4609 = io_x[10] ? _GEN4608 : _GEN4606;
wire  _GEN4610 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4611 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4612 = io_x[14] ? _GEN4611 : _GEN4610;
wire  _GEN4613 = io_x[10] ? _GEN4612 : _GEN3711;
wire  _GEN4614 = io_x[23] ? _GEN4613 : _GEN4609;
wire  _GEN4615 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4616 = io_x[14] ? _GEN3709 : _GEN4615;
wire  _GEN4617 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4618 = io_x[14] ? _GEN4617 : _GEN3709;
wire  _GEN4619 = io_x[10] ? _GEN4618 : _GEN4616;
wire  _GEN4620 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4621 = io_x[14] ? _GEN4620 : _GEN3709;
wire  _GEN4622 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4623 = io_x[10] ? _GEN4622 : _GEN4621;
wire  _GEN4624 = io_x[23] ? _GEN4623 : _GEN4619;
wire  _GEN4625 = io_x[16] ? _GEN4624 : _GEN4614;
wire  _GEN4626 = io_x[12] ? _GEN4625 : _GEN4605;
wire  _GEN4627 = io_x[2] ? _GEN4626 : _GEN4593;
wire  _GEN4628 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4629 = io_x[14] ? _GEN4628 : _GEN3709;
wire  _GEN4630 = io_x[10] ? _GEN3716 : _GEN4629;
wire  _GEN4631 = io_x[23] ? _GEN4630 : _GEN3741;
wire  _GEN4632 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4633 = io_x[14] ? _GEN3709 : _GEN4632;
wire  _GEN4634 = io_x[10] ? _GEN3711 : _GEN4633;
wire  _GEN4635 = io_x[23] ? _GEN3713 : _GEN4634;
wire  _GEN4636 = io_x[16] ? _GEN4635 : _GEN4631;
wire  _GEN4637 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4638 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4639 = io_x[14] ? _GEN4638 : _GEN3708;
wire  _GEN4640 = io_x[10] ? _GEN4639 : _GEN4637;
wire  _GEN4641 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4642 = io_x[10] ? _GEN4641 : _GEN3711;
wire  _GEN4643 = io_x[23] ? _GEN4642 : _GEN4640;
wire  _GEN4644 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4645 = io_x[14] ? _GEN4644 : _GEN3708;
wire  _GEN4646 = io_x[10] ? _GEN4645 : _GEN3716;
wire  _GEN4647 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4648 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4649 = io_x[10] ? _GEN4648 : _GEN4647;
wire  _GEN4650 = io_x[23] ? _GEN4649 : _GEN4646;
wire  _GEN4651 = io_x[16] ? _GEN4650 : _GEN4643;
wire  _GEN4652 = io_x[12] ? _GEN4651 : _GEN4636;
wire  _GEN4653 = io_x[23] ? _GEN3713 : _GEN3741;
wire  _GEN4654 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4655 = io_x[14] ? _GEN4654 : _GEN3709;
wire  _GEN4656 = io_x[10] ? _GEN4655 : _GEN3711;
wire  _GEN4657 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4658 = io_x[14] ? _GEN4657 : _GEN3708;
wire  _GEN4659 = io_x[10] ? _GEN3716 : _GEN4658;
wire  _GEN4660 = io_x[23] ? _GEN4659 : _GEN4656;
wire  _GEN4661 = io_x[16] ? _GEN4660 : _GEN4653;
wire  _GEN4662 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4663 = io_x[14] ? _GEN4662 : _GEN3708;
wire  _GEN4664 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4665 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4666 = io_x[14] ? _GEN4665 : _GEN4664;
wire  _GEN4667 = io_x[10] ? _GEN4666 : _GEN4663;
wire  _GEN4668 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4669 = io_x[14] ? _GEN3709 : _GEN4668;
wire  _GEN4670 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4671 = io_x[14] ? _GEN3708 : _GEN4670;
wire  _GEN4672 = io_x[10] ? _GEN4671 : _GEN4669;
wire  _GEN4673 = io_x[23] ? _GEN4672 : _GEN4667;
wire  _GEN4674 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4675 = io_x[14] ? _GEN4674 : _GEN3708;
wire  _GEN4676 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4677 = io_x[14] ? _GEN4676 : _GEN3709;
wire  _GEN4678 = io_x[10] ? _GEN4677 : _GEN4675;
wire  _GEN4679 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4680 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4681 = io_x[14] ? _GEN4680 : _GEN4679;
wire  _GEN4682 = io_x[10] ? _GEN4681 : _GEN3716;
wire  _GEN4683 = io_x[23] ? _GEN4682 : _GEN4678;
wire  _GEN4684 = io_x[16] ? _GEN4683 : _GEN4673;
wire  _GEN4685 = io_x[12] ? _GEN4684 : _GEN4661;
wire  _GEN4686 = io_x[2] ? _GEN4685 : _GEN4652;
wire  _GEN4687 = io_x[9] ? _GEN4686 : _GEN4627;
wire  _GEN4688 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4689 = io_x[14] ? _GEN3708 : _GEN4688;
wire  _GEN4690 = io_x[10] ? _GEN4689 : _GEN3711;
wire  _GEN4691 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4692 = io_x[10] ? _GEN3711 : _GEN4691;
wire  _GEN4693 = io_x[23] ? _GEN4692 : _GEN4690;
wire  _GEN4694 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4695 = io_x[14] ? _GEN4694 : _GEN3709;
wire  _GEN4696 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4697 = io_x[14] ? _GEN3709 : _GEN4696;
wire  _GEN4698 = io_x[10] ? _GEN4697 : _GEN4695;
wire  _GEN4699 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4700 = io_x[10] ? _GEN4699 : _GEN3711;
wire  _GEN4701 = io_x[23] ? _GEN4700 : _GEN4698;
wire  _GEN4702 = io_x[16] ? _GEN4701 : _GEN4693;
wire  _GEN4703 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4704 = io_x[10] ? _GEN4703 : _GEN3711;
wire  _GEN4705 = io_x[23] ? _GEN4704 : _GEN3741;
wire  _GEN4706 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4707 = io_x[14] ? _GEN4706 : _GEN3708;
wire  _GEN4708 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4709 = io_x[14] ? _GEN4708 : _GEN3709;
wire  _GEN4710 = io_x[10] ? _GEN4709 : _GEN4707;
wire  _GEN4711 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN4712 = io_x[23] ? _GEN4711 : _GEN4710;
wire  _GEN4713 = io_x[16] ? _GEN4712 : _GEN4705;
wire  _GEN4714 = io_x[12] ? _GEN4713 : _GEN4702;
wire  _GEN4715 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4716 = io_x[14] ? _GEN4715 : _GEN3709;
wire  _GEN4717 = io_x[10] ? _GEN4716 : _GEN3711;
wire  _GEN4718 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4719 = io_x[10] ? _GEN3711 : _GEN4718;
wire  _GEN4720 = io_x[23] ? _GEN4719 : _GEN4717;
wire  _GEN4721 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4722 = io_x[10] ? _GEN4721 : _GEN3711;
wire  _GEN4723 = io_x[23] ? _GEN4722 : _GEN3741;
wire  _GEN4724 = io_x[16] ? _GEN4723 : _GEN4720;
wire  _GEN4725 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4726 = io_x[14] ? _GEN3708 : _GEN4725;
wire  _GEN4727 = io_x[10] ? _GEN4726 : _GEN3716;
wire  _GEN4728 = io_x[23] ? _GEN3741 : _GEN4727;
wire  _GEN4729 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4730 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4731 = io_x[14] ? _GEN4730 : _GEN4729;
wire  _GEN4732 = io_x[10] ? _GEN3716 : _GEN4731;
wire  _GEN4733 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4734 = io_x[10] ? _GEN4733 : _GEN3716;
wire  _GEN4735 = io_x[23] ? _GEN4734 : _GEN4732;
wire  _GEN4736 = io_x[16] ? _GEN4735 : _GEN4728;
wire  _GEN4737 = io_x[12] ? _GEN4736 : _GEN4724;
wire  _GEN4738 = io_x[2] ? _GEN4737 : _GEN4714;
wire  _GEN4739 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4740 = io_x[14] ? _GEN4739 : _GEN3709;
wire  _GEN4741 = io_x[10] ? _GEN3711 : _GEN4740;
wire  _GEN4742 = io_x[23] ? _GEN3741 : _GEN4741;
wire  _GEN4743 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4744 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4745 = io_x[14] ? _GEN4744 : _GEN4743;
wire  _GEN4746 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4747 = io_x[14] ? _GEN4746 : _GEN3709;
wire  _GEN4748 = io_x[10] ? _GEN4747 : _GEN4745;
wire  _GEN4749 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4750 = io_x[14] ? _GEN4749 : _GEN3709;
wire  _GEN4751 = io_x[10] ? _GEN4750 : _GEN3716;
wire  _GEN4752 = io_x[23] ? _GEN4751 : _GEN4748;
wire  _GEN4753 = io_x[16] ? _GEN4752 : _GEN4742;
wire  _GEN4754 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4755 = io_x[14] ? _GEN4754 : _GEN3709;
wire  _GEN4756 = io_x[10] ? _GEN4755 : _GEN3716;
wire  _GEN4757 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4758 = io_x[14] ? _GEN4757 : _GEN3709;
wire  _GEN4759 = io_x[10] ? _GEN4758 : _GEN3711;
wire  _GEN4760 = io_x[23] ? _GEN4759 : _GEN4756;
wire  _GEN4761 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4762 = io_x[14] ? _GEN4761 : _GEN3708;
wire  _GEN4763 = io_x[10] ? _GEN4762 : _GEN3716;
wire  _GEN4764 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4765 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4766 = io_x[14] ? _GEN4765 : _GEN4764;
wire  _GEN4767 = io_x[10] ? _GEN4766 : _GEN3711;
wire  _GEN4768 = io_x[23] ? _GEN4767 : _GEN4763;
wire  _GEN4769 = io_x[16] ? _GEN4768 : _GEN4760;
wire  _GEN4770 = io_x[12] ? _GEN4769 : _GEN4753;
wire  _GEN4771 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4772 = io_x[10] ? _GEN4771 : _GEN3711;
wire  _GEN4773 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4774 = io_x[14] ? _GEN3709 : _GEN4773;
wire  _GEN4775 = io_x[10] ? _GEN3711 : _GEN4774;
wire  _GEN4776 = io_x[23] ? _GEN4775 : _GEN4772;
wire  _GEN4777 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4778 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4779 = io_x[10] ? _GEN4778 : _GEN4777;
wire  _GEN4780 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4781 = io_x[10] ? _GEN4780 : _GEN3711;
wire  _GEN4782 = io_x[23] ? _GEN4781 : _GEN4779;
wire  _GEN4783 = io_x[16] ? _GEN4782 : _GEN4776;
wire  _GEN4784 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4785 = io_x[14] ? _GEN4784 : _GEN3709;
wire  _GEN4786 = io_x[10] ? _GEN4785 : _GEN3711;
wire  _GEN4787 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4788 = io_x[14] ? _GEN4787 : _GEN3709;
wire  _GEN4789 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4790 = io_x[10] ? _GEN4789 : _GEN4788;
wire  _GEN4791 = io_x[23] ? _GEN4790 : _GEN4786;
wire  _GEN4792 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4793 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4794 = io_x[14] ? _GEN4793 : _GEN4792;
wire  _GEN4795 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4796 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4797 = io_x[14] ? _GEN4796 : _GEN4795;
wire  _GEN4798 = io_x[10] ? _GEN4797 : _GEN4794;
wire  _GEN4799 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4800 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4801 = io_x[14] ? _GEN4800 : _GEN4799;
wire  _GEN4802 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4803 = io_x[14] ? _GEN4802 : _GEN3709;
wire  _GEN4804 = io_x[10] ? _GEN4803 : _GEN4801;
wire  _GEN4805 = io_x[23] ? _GEN4804 : _GEN4798;
wire  _GEN4806 = io_x[16] ? _GEN4805 : _GEN4791;
wire  _GEN4807 = io_x[12] ? _GEN4806 : _GEN4783;
wire  _GEN4808 = io_x[2] ? _GEN4807 : _GEN4770;
wire  _GEN4809 = io_x[9] ? _GEN4808 : _GEN4738;
wire  _GEN4810 = io_x[13] ? _GEN4809 : _GEN4687;
wire  _GEN4811 = io_x[7] ? _GEN4810 : _GEN4581;
wire  _GEN4812 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4813 = io_x[10] ? _GEN4812 : _GEN3711;
wire  _GEN4814 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4815 = io_x[10] ? _GEN3711 : _GEN4814;
wire  _GEN4816 = io_x[23] ? _GEN4815 : _GEN4813;
wire  _GEN4817 = io_x[16] ? _GEN4816 : _GEN3727;
wire  _GEN4818 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4819 = io_x[10] ? _GEN4818 : _GEN3711;
wire  _GEN4820 = io_x[23] ? _GEN3713 : _GEN4819;
wire  _GEN4821 = io_x[16] ? _GEN4820 : _GEN3707;
wire  _GEN4822 = io_x[12] ? _GEN4821 : _GEN4817;
wire  _GEN4823 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4824 = io_x[10] ? _GEN4823 : _GEN3711;
wire  _GEN4825 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4826 = io_x[14] ? _GEN4825 : _GEN3709;
wire  _GEN4827 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4828 = io_x[10] ? _GEN4827 : _GEN4826;
wire  _GEN4829 = io_x[23] ? _GEN4828 : _GEN4824;
wire  _GEN4830 = io_x[16] ? _GEN4829 : _GEN3727;
wire  _GEN4831 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN4832 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4833 = io_x[14] ? _GEN4832 : _GEN3709;
wire  _GEN4834 = io_x[10] ? _GEN4833 : _GEN3711;
wire  _GEN4835 = io_x[23] ? _GEN4834 : _GEN4831;
wire  _GEN4836 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4837 = io_x[14] ? _GEN4836 : _GEN3708;
wire  _GEN4838 = io_x[10] ? _GEN4837 : _GEN3716;
wire  _GEN4839 = io_x[23] ? _GEN4838 : _GEN3741;
wire  _GEN4840 = io_x[16] ? _GEN4839 : _GEN4835;
wire  _GEN4841 = io_x[12] ? _GEN4840 : _GEN4830;
wire  _GEN4842 = io_x[2] ? _GEN4841 : _GEN4822;
wire  _GEN4843 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN4844 = io_x[23] ? _GEN3741 : _GEN4843;
wire  _GEN4845 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4846 = io_x[14] ? _GEN4845 : _GEN3709;
wire  _GEN4847 = io_x[10] ? _GEN3711 : _GEN4846;
wire  _GEN4848 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4849 = io_x[10] ? _GEN3716 : _GEN4848;
wire  _GEN4850 = io_x[23] ? _GEN4849 : _GEN4847;
wire  _GEN4851 = io_x[16] ? _GEN4850 : _GEN4844;
wire  _GEN4852 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4853 = io_x[14] ? _GEN4852 : _GEN3709;
wire  _GEN4854 = io_x[10] ? _GEN3716 : _GEN4853;
wire  _GEN4855 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4856 = io_x[14] ? _GEN3709 : _GEN4855;
wire  _GEN4857 = io_x[10] ? _GEN3711 : _GEN4856;
wire  _GEN4858 = io_x[23] ? _GEN4857 : _GEN4854;
wire  _GEN4859 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4860 = io_x[14] ? _GEN4859 : _GEN3709;
wire  _GEN4861 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4862 = io_x[14] ? _GEN4861 : _GEN3709;
wire  _GEN4863 = io_x[10] ? _GEN4862 : _GEN4860;
wire  _GEN4864 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4865 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4866 = io_x[14] ? _GEN4865 : _GEN3709;
wire  _GEN4867 = io_x[10] ? _GEN4866 : _GEN4864;
wire  _GEN4868 = io_x[23] ? _GEN4867 : _GEN4863;
wire  _GEN4869 = io_x[16] ? _GEN4868 : _GEN4858;
wire  _GEN4870 = io_x[12] ? _GEN4869 : _GEN4851;
wire  _GEN4871 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4872 = io_x[14] ? _GEN4871 : _GEN3709;
wire  _GEN4873 = io_x[10] ? _GEN4872 : _GEN3711;
wire  _GEN4874 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4875 = io_x[10] ? _GEN3716 : _GEN4874;
wire  _GEN4876 = io_x[23] ? _GEN4875 : _GEN4873;
wire  _GEN4877 = io_x[16] ? _GEN4876 : _GEN3707;
wire  _GEN4878 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4879 = io_x[14] ? _GEN3709 : _GEN4878;
wire  _GEN4880 = io_x[10] ? _GEN3716 : _GEN4879;
wire  _GEN4881 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4882 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4883 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4884 = io_x[14] ? _GEN4883 : _GEN4882;
wire  _GEN4885 = io_x[10] ? _GEN4884 : _GEN4881;
wire  _GEN4886 = io_x[23] ? _GEN4885 : _GEN4880;
wire  _GEN4887 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4888 = io_x[10] ? _GEN4887 : _GEN3711;
wire  _GEN4889 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4890 = io_x[14] ? _GEN3709 : _GEN4889;
wire  _GEN4891 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4892 = io_x[14] ? _GEN4891 : _GEN3709;
wire  _GEN4893 = io_x[10] ? _GEN4892 : _GEN4890;
wire  _GEN4894 = io_x[23] ? _GEN4893 : _GEN4888;
wire  _GEN4895 = io_x[16] ? _GEN4894 : _GEN4886;
wire  _GEN4896 = io_x[12] ? _GEN4895 : _GEN4877;
wire  _GEN4897 = io_x[2] ? _GEN4896 : _GEN4870;
wire  _GEN4898 = io_x[9] ? _GEN4897 : _GEN4842;
wire  _GEN4899 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4900 = io_x[14] ? _GEN4899 : _GEN3708;
wire  _GEN4901 = io_x[10] ? _GEN4900 : _GEN3711;
wire  _GEN4902 = io_x[23] ? _GEN3713 : _GEN4901;
wire  _GEN4903 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4904 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4905 = io_x[14] ? _GEN4904 : _GEN4903;
wire  _GEN4906 = io_x[10] ? _GEN4905 : _GEN3711;
wire  _GEN4907 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4908 = io_x[14] ? _GEN3709 : _GEN4907;
wire  _GEN4909 = io_x[10] ? _GEN4908 : _GEN3711;
wire  _GEN4910 = io_x[23] ? _GEN4909 : _GEN4906;
wire  _GEN4911 = io_x[16] ? _GEN4910 : _GEN4902;
wire  _GEN4912 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN4913 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4914 = io_x[10] ? _GEN3711 : _GEN4913;
wire  _GEN4915 = io_x[23] ? _GEN4914 : _GEN4912;
wire  _GEN4916 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4917 = io_x[14] ? _GEN4916 : _GEN3708;
wire  _GEN4918 = io_x[10] ? _GEN4917 : _GEN3716;
wire  _GEN4919 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4920 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4921 = io_x[14] ? _GEN4920 : _GEN4919;
wire  _GEN4922 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4923 = io_x[10] ? _GEN4922 : _GEN4921;
wire  _GEN4924 = io_x[23] ? _GEN4923 : _GEN4918;
wire  _GEN4925 = io_x[16] ? _GEN4924 : _GEN4915;
wire  _GEN4926 = io_x[12] ? _GEN4925 : _GEN4911;
wire  _GEN4927 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4928 = io_x[14] ? _GEN4927 : _GEN3709;
wire  _GEN4929 = io_x[10] ? _GEN4928 : _GEN3711;
wire  _GEN4930 = io_x[23] ? _GEN3713 : _GEN4929;
wire  _GEN4931 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4932 = io_x[10] ? _GEN4931 : _GEN3711;
wire  _GEN4933 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4934 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4935 = io_x[14] ? _GEN3708 : _GEN4934;
wire  _GEN4936 = io_x[10] ? _GEN4935 : _GEN4933;
wire  _GEN4937 = io_x[23] ? _GEN4936 : _GEN4932;
wire  _GEN4938 = io_x[16] ? _GEN4937 : _GEN4930;
wire  _GEN4939 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4940 = io_x[14] ? _GEN4939 : _GEN3709;
wire  _GEN4941 = io_x[10] ? _GEN4940 : _GEN3716;
wire  _GEN4942 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4943 = io_x[14] ? _GEN4942 : _GEN3708;
wire  _GEN4944 = io_x[10] ? _GEN4943 : _GEN3711;
wire  _GEN4945 = io_x[23] ? _GEN4944 : _GEN4941;
wire  _GEN4946 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4947 = io_x[14] ? _GEN4946 : _GEN3709;
wire  _GEN4948 = io_x[10] ? _GEN4947 : _GEN3711;
wire  _GEN4949 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4950 = io_x[14] ? _GEN4949 : _GEN3709;
wire  _GEN4951 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4952 = io_x[14] ? _GEN3708 : _GEN4951;
wire  _GEN4953 = io_x[10] ? _GEN4952 : _GEN4950;
wire  _GEN4954 = io_x[23] ? _GEN4953 : _GEN4948;
wire  _GEN4955 = io_x[16] ? _GEN4954 : _GEN4945;
wire  _GEN4956 = io_x[12] ? _GEN4955 : _GEN4938;
wire  _GEN4957 = io_x[2] ? _GEN4956 : _GEN4926;
wire  _GEN4958 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN4959 = io_x[10] ? _GEN4958 : _GEN3716;
wire  _GEN4960 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4961 = io_x[14] ? _GEN3709 : _GEN4960;
wire  _GEN4962 = io_x[10] ? _GEN3711 : _GEN4961;
wire  _GEN4963 = io_x[23] ? _GEN4962 : _GEN4959;
wire  _GEN4964 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4965 = io_x[14] ? _GEN3709 : _GEN4964;
wire  _GEN4966 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4967 = io_x[14] ? _GEN4966 : _GEN3709;
wire  _GEN4968 = io_x[10] ? _GEN4967 : _GEN4965;
wire  _GEN4969 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4970 = io_x[14] ? _GEN3709 : _GEN4969;
wire  _GEN4971 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4972 = io_x[10] ? _GEN4971 : _GEN4970;
wire  _GEN4973 = io_x[23] ? _GEN4972 : _GEN4968;
wire  _GEN4974 = io_x[16] ? _GEN4973 : _GEN4963;
wire  _GEN4975 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4976 = io_x[14] ? _GEN4975 : _GEN3708;
wire  _GEN4977 = io_x[10] ? _GEN4976 : _GEN3711;
wire  _GEN4978 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4979 = io_x[14] ? _GEN3709 : _GEN4978;
wire  _GEN4980 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN4981 = io_x[10] ? _GEN4980 : _GEN4979;
wire  _GEN4982 = io_x[23] ? _GEN4981 : _GEN4977;
wire  _GEN4983 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4984 = io_x[14] ? _GEN4983 : _GEN3709;
wire  _GEN4985 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4986 = io_x[14] ? _GEN4985 : _GEN3708;
wire  _GEN4987 = io_x[10] ? _GEN4986 : _GEN4984;
wire  _GEN4988 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4989 = io_x[14] ? _GEN4988 : _GEN3709;
wire  _GEN4990 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN4991 = io_x[14] ? _GEN4990 : _GEN3708;
wire  _GEN4992 = io_x[10] ? _GEN4991 : _GEN4989;
wire  _GEN4993 = io_x[23] ? _GEN4992 : _GEN4987;
wire  _GEN4994 = io_x[16] ? _GEN4993 : _GEN4982;
wire  _GEN4995 = io_x[12] ? _GEN4994 : _GEN4974;
wire  _GEN4996 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN4997 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN4998 = io_x[14] ? _GEN4997 : _GEN3709;
wire  _GEN4999 = io_x[10] ? _GEN4998 : _GEN3716;
wire  _GEN5000 = io_x[23] ? _GEN4999 : _GEN4996;
wire  _GEN5001 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5002 = io_x[14] ? _GEN3709 : _GEN5001;
wire  _GEN5003 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5004 = io_x[14] ? _GEN5003 : _GEN3709;
wire  _GEN5005 = io_x[10] ? _GEN5004 : _GEN5002;
wire  _GEN5006 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5007 = io_x[10] ? _GEN3716 : _GEN5006;
wire  _GEN5008 = io_x[23] ? _GEN5007 : _GEN5005;
wire  _GEN5009 = io_x[16] ? _GEN5008 : _GEN5000;
wire  _GEN5010 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5011 = io_x[14] ? _GEN5010 : _GEN3708;
wire  _GEN5012 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5013 = io_x[14] ? _GEN5012 : _GEN3709;
wire  _GEN5014 = io_x[10] ? _GEN5013 : _GEN5011;
wire  _GEN5015 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5016 = io_x[14] ? _GEN3709 : _GEN5015;
wire  _GEN5017 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5018 = io_x[14] ? _GEN5017 : _GEN3709;
wire  _GEN5019 = io_x[10] ? _GEN5018 : _GEN5016;
wire  _GEN5020 = io_x[23] ? _GEN5019 : _GEN5014;
wire  _GEN5021 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5022 = io_x[14] ? _GEN5021 : _GEN3709;
wire  _GEN5023 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5024 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5025 = io_x[14] ? _GEN5024 : _GEN5023;
wire  _GEN5026 = io_x[10] ? _GEN5025 : _GEN5022;
wire  _GEN5027 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5028 = io_x[14] ? _GEN5027 : _GEN3708;
wire  _GEN5029 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5030 = io_x[14] ? _GEN5029 : _GEN3709;
wire  _GEN5031 = io_x[10] ? _GEN5030 : _GEN5028;
wire  _GEN5032 = io_x[23] ? _GEN5031 : _GEN5026;
wire  _GEN5033 = io_x[16] ? _GEN5032 : _GEN5020;
wire  _GEN5034 = io_x[12] ? _GEN5033 : _GEN5009;
wire  _GEN5035 = io_x[2] ? _GEN5034 : _GEN4995;
wire  _GEN5036 = io_x[9] ? _GEN5035 : _GEN4957;
wire  _GEN5037 = io_x[13] ? _GEN5036 : _GEN4898;
wire  _GEN5038 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5039 = io_x[14] ? _GEN5038 : _GEN3709;
wire  _GEN5040 = io_x[10] ? _GEN5039 : _GEN3711;
wire  _GEN5041 = io_x[23] ? _GEN5040 : _GEN3741;
wire  _GEN5042 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5043 = io_x[14] ? _GEN3709 : _GEN5042;
wire  _GEN5044 = io_x[10] ? _GEN3711 : _GEN5043;
wire  _GEN5045 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN5046 = io_x[23] ? _GEN5045 : _GEN5044;
wire  _GEN5047 = io_x[16] ? _GEN5046 : _GEN5041;
wire  _GEN5048 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5049 = io_x[10] ? _GEN5048 : _GEN3716;
wire  _GEN5050 = io_x[23] ? _GEN3713 : _GEN5049;
wire  _GEN5051 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN5052 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5053 = io_x[10] ? _GEN5052 : _GEN3716;
wire  _GEN5054 = io_x[23] ? _GEN5053 : _GEN5051;
wire  _GEN5055 = io_x[16] ? _GEN5054 : _GEN5050;
wire  _GEN5056 = io_x[12] ? _GEN5055 : _GEN5047;
wire  _GEN5057 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5058 = io_x[14] ? _GEN3709 : _GEN5057;
wire  _GEN5059 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5060 = io_x[10] ? _GEN5059 : _GEN5058;
wire  _GEN5061 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5062 = io_x[10] ? _GEN5061 : _GEN3711;
wire  _GEN5063 = io_x[23] ? _GEN5062 : _GEN5060;
wire  _GEN5064 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5065 = io_x[14] ? _GEN5064 : _GEN3708;
wire  _GEN5066 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5067 = io_x[10] ? _GEN5066 : _GEN5065;
wire  _GEN5068 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5069 = io_x[10] ? _GEN5068 : _GEN3716;
wire  _GEN5070 = io_x[23] ? _GEN5069 : _GEN5067;
wire  _GEN5071 = io_x[16] ? _GEN5070 : _GEN5063;
wire  _GEN5072 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5073 = io_x[14] ? _GEN5072 : _GEN3709;
wire  _GEN5074 = io_x[10] ? _GEN5073 : _GEN3716;
wire  _GEN5075 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5076 = io_x[14] ? _GEN5075 : _GEN3708;
wire  _GEN5077 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5078 = io_x[10] ? _GEN5077 : _GEN5076;
wire  _GEN5079 = io_x[23] ? _GEN5078 : _GEN5074;
wire  _GEN5080 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5081 = io_x[14] ? _GEN5080 : _GEN3708;
wire  _GEN5082 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5083 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5084 = io_x[14] ? _GEN5083 : _GEN5082;
wire  _GEN5085 = io_x[10] ? _GEN5084 : _GEN5081;
wire  _GEN5086 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5087 = io_x[14] ? _GEN3708 : _GEN5086;
wire  _GEN5088 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5089 = io_x[10] ? _GEN5088 : _GEN5087;
wire  _GEN5090 = io_x[23] ? _GEN5089 : _GEN5085;
wire  _GEN5091 = io_x[16] ? _GEN5090 : _GEN5079;
wire  _GEN5092 = io_x[12] ? _GEN5091 : _GEN5071;
wire  _GEN5093 = io_x[2] ? _GEN5092 : _GEN5056;
wire  _GEN5094 = io_x[23] ? _GEN3741 : _GEN3713;
wire  _GEN5095 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5096 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5097 = io_x[14] ? _GEN5096 : _GEN5095;
wire  _GEN5098 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5099 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5100 = io_x[14] ? _GEN5099 : _GEN5098;
wire  _GEN5101 = io_x[10] ? _GEN5100 : _GEN5097;
wire  _GEN5102 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5103 = io_x[14] ? _GEN5102 : _GEN3709;
wire  _GEN5104 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5105 = io_x[10] ? _GEN5104 : _GEN5103;
wire  _GEN5106 = io_x[23] ? _GEN5105 : _GEN5101;
wire  _GEN5107 = io_x[16] ? _GEN5106 : _GEN5094;
wire  _GEN5108 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5109 = io_x[10] ? _GEN3711 : _GEN5108;
wire  _GEN5110 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5111 = io_x[10] ? _GEN5110 : _GEN3711;
wire  _GEN5112 = io_x[23] ? _GEN5111 : _GEN5109;
wire  _GEN5113 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5114 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5115 = io_x[14] ? _GEN5114 : _GEN5113;
wire  _GEN5116 = io_x[10] ? _GEN5115 : _GEN3716;
wire  _GEN5117 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5118 = io_x[10] ? _GEN5117 : _GEN3711;
wire  _GEN5119 = io_x[23] ? _GEN5118 : _GEN5116;
wire  _GEN5120 = io_x[16] ? _GEN5119 : _GEN5112;
wire  _GEN5121 = io_x[12] ? _GEN5120 : _GEN5107;
wire  _GEN5122 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5123 = io_x[14] ? _GEN5122 : _GEN3709;
wire  _GEN5124 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5125 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5126 = io_x[14] ? _GEN5125 : _GEN5124;
wire  _GEN5127 = io_x[10] ? _GEN5126 : _GEN5123;
wire  _GEN5128 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5129 = io_x[14] ? _GEN5128 : _GEN3709;
wire  _GEN5130 = io_x[10] ? _GEN5129 : _GEN3711;
wire  _GEN5131 = io_x[23] ? _GEN5130 : _GEN5127;
wire  _GEN5132 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5133 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5134 = io_x[14] ? _GEN5133 : _GEN3709;
wire  _GEN5135 = io_x[10] ? _GEN5134 : _GEN5132;
wire  _GEN5136 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5137 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5138 = io_x[14] ? _GEN3708 : _GEN5137;
wire  _GEN5139 = io_x[10] ? _GEN5138 : _GEN5136;
wire  _GEN5140 = io_x[23] ? _GEN5139 : _GEN5135;
wire  _GEN5141 = io_x[16] ? _GEN5140 : _GEN5131;
wire  _GEN5142 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5143 = io_x[14] ? _GEN5142 : _GEN3709;
wire  _GEN5144 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5145 = io_x[14] ? _GEN5144 : _GEN3709;
wire  _GEN5146 = io_x[10] ? _GEN5145 : _GEN5143;
wire  _GEN5147 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5148 = io_x[14] ? _GEN3709 : _GEN5147;
wire  _GEN5149 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5150 = io_x[14] ? _GEN5149 : _GEN3709;
wire  _GEN5151 = io_x[10] ? _GEN5150 : _GEN5148;
wire  _GEN5152 = io_x[23] ? _GEN5151 : _GEN5146;
wire  _GEN5153 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5154 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5155 = io_x[14] ? _GEN5154 : _GEN5153;
wire  _GEN5156 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5157 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5158 = io_x[14] ? _GEN5157 : _GEN5156;
wire  _GEN5159 = io_x[10] ? _GEN5158 : _GEN5155;
wire  _GEN5160 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5161 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5162 = io_x[14] ? _GEN5161 : _GEN5160;
wire  _GEN5163 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5164 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5165 = io_x[14] ? _GEN5164 : _GEN5163;
wire  _GEN5166 = io_x[10] ? _GEN5165 : _GEN5162;
wire  _GEN5167 = io_x[23] ? _GEN5166 : _GEN5159;
wire  _GEN5168 = io_x[16] ? _GEN5167 : _GEN5152;
wire  _GEN5169 = io_x[12] ? _GEN5168 : _GEN5141;
wire  _GEN5170 = io_x[2] ? _GEN5169 : _GEN5121;
wire  _GEN5171 = io_x[9] ? _GEN5170 : _GEN5093;
wire  _GEN5172 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5173 = io_x[14] ? _GEN5172 : _GEN3709;
wire  _GEN5174 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5175 = io_x[14] ? _GEN3709 : _GEN5174;
wire  _GEN5176 = io_x[10] ? _GEN5175 : _GEN5173;
wire  _GEN5177 = io_x[23] ? _GEN3713 : _GEN5176;
wire  _GEN5178 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5179 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5180 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5181 = io_x[14] ? _GEN5180 : _GEN5179;
wire  _GEN5182 = io_x[10] ? _GEN5181 : _GEN5178;
wire  _GEN5183 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5184 = io_x[14] ? _GEN5183 : _GEN3709;
wire  _GEN5185 = io_x[10] ? _GEN5184 : _GEN3716;
wire  _GEN5186 = io_x[23] ? _GEN5185 : _GEN5182;
wire  _GEN5187 = io_x[16] ? _GEN5186 : _GEN5177;
wire  _GEN5188 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5189 = io_x[14] ? _GEN5188 : _GEN3709;
wire  _GEN5190 = io_x[10] ? _GEN5189 : _GEN3711;
wire  _GEN5191 = io_x[23] ? _GEN3741 : _GEN5190;
wire  _GEN5192 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5193 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5194 = io_x[14] ? _GEN5193 : _GEN5192;
wire  _GEN5195 = io_x[10] ? _GEN5194 : _GEN3711;
wire  _GEN5196 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5197 = io_x[14] ? _GEN5196 : _GEN3709;
wire  _GEN5198 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5199 = io_x[14] ? _GEN5198 : _GEN3708;
wire  _GEN5200 = io_x[10] ? _GEN5199 : _GEN5197;
wire  _GEN5201 = io_x[23] ? _GEN5200 : _GEN5195;
wire  _GEN5202 = io_x[16] ? _GEN5201 : _GEN5191;
wire  _GEN5203 = io_x[12] ? _GEN5202 : _GEN5187;
wire  _GEN5204 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5205 = io_x[10] ? _GEN3716 : _GEN5204;
wire  _GEN5206 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5207 = io_x[14] ? _GEN3708 : _GEN5206;
wire  _GEN5208 = io_x[10] ? _GEN5207 : _GEN3711;
wire  _GEN5209 = io_x[23] ? _GEN5208 : _GEN5205;
wire  _GEN5210 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5211 = io_x[14] ? _GEN5210 : _GEN3709;
wire  _GEN5212 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5213 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5214 = io_x[14] ? _GEN5213 : _GEN5212;
wire  _GEN5215 = io_x[10] ? _GEN5214 : _GEN5211;
wire  _GEN5216 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5217 = io_x[10] ? _GEN3716 : _GEN5216;
wire  _GEN5218 = io_x[23] ? _GEN5217 : _GEN5215;
wire  _GEN5219 = io_x[16] ? _GEN5218 : _GEN5209;
wire  _GEN5220 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5221 = io_x[14] ? _GEN5220 : _GEN3708;
wire  _GEN5222 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5223 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5224 = io_x[14] ? _GEN5223 : _GEN5222;
wire  _GEN5225 = io_x[10] ? _GEN5224 : _GEN5221;
wire  _GEN5226 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5227 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5228 = io_x[14] ? _GEN5227 : _GEN5226;
wire  _GEN5229 = io_x[10] ? _GEN5228 : _GEN3711;
wire  _GEN5230 = io_x[23] ? _GEN5229 : _GEN5225;
wire  _GEN5231 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5232 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5233 = io_x[14] ? _GEN5232 : _GEN5231;
wire  _GEN5234 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5235 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5236 = io_x[14] ? _GEN5235 : _GEN5234;
wire  _GEN5237 = io_x[10] ? _GEN5236 : _GEN5233;
wire  _GEN5238 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5239 = io_x[14] ? _GEN5238 : _GEN3709;
wire  _GEN5240 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5241 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5242 = io_x[14] ? _GEN5241 : _GEN5240;
wire  _GEN5243 = io_x[10] ? _GEN5242 : _GEN5239;
wire  _GEN5244 = io_x[23] ? _GEN5243 : _GEN5237;
wire  _GEN5245 = io_x[16] ? _GEN5244 : _GEN5230;
wire  _GEN5246 = io_x[12] ? _GEN5245 : _GEN5219;
wire  _GEN5247 = io_x[2] ? _GEN5246 : _GEN5203;
wire  _GEN5248 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5249 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5250 = io_x[14] ? _GEN5249 : _GEN5248;
wire  _GEN5251 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5252 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5253 = io_x[14] ? _GEN5252 : _GEN5251;
wire  _GEN5254 = io_x[10] ? _GEN5253 : _GEN5250;
wire  _GEN5255 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5256 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5257 = io_x[14] ? _GEN3708 : _GEN5256;
wire  _GEN5258 = io_x[10] ? _GEN5257 : _GEN5255;
wire  _GEN5259 = io_x[23] ? _GEN5258 : _GEN5254;
wire  _GEN5260 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5261 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5262 = io_x[14] ? _GEN5261 : _GEN5260;
wire  _GEN5263 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5264 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5265 = io_x[14] ? _GEN5264 : _GEN5263;
wire  _GEN5266 = io_x[10] ? _GEN5265 : _GEN5262;
wire  _GEN5267 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5268 = io_x[14] ? _GEN3709 : _GEN5267;
wire  _GEN5269 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5270 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5271 = io_x[14] ? _GEN5270 : _GEN5269;
wire  _GEN5272 = io_x[10] ? _GEN5271 : _GEN5268;
wire  _GEN5273 = io_x[23] ? _GEN5272 : _GEN5266;
wire  _GEN5274 = io_x[16] ? _GEN5273 : _GEN5259;
wire  _GEN5275 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5276 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5277 = io_x[14] ? _GEN5276 : _GEN5275;
wire  _GEN5278 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5279 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5280 = io_x[14] ? _GEN5279 : _GEN5278;
wire  _GEN5281 = io_x[10] ? _GEN5280 : _GEN5277;
wire  _GEN5282 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5283 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5284 = io_x[10] ? _GEN5283 : _GEN5282;
wire  _GEN5285 = io_x[23] ? _GEN5284 : _GEN5281;
wire  _GEN5286 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5287 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5288 = io_x[14] ? _GEN5287 : _GEN5286;
wire  _GEN5289 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5290 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5291 = io_x[14] ? _GEN5290 : _GEN5289;
wire  _GEN5292 = io_x[10] ? _GEN5291 : _GEN5288;
wire  _GEN5293 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5294 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5295 = io_x[14] ? _GEN5294 : _GEN5293;
wire  _GEN5296 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5297 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5298 = io_x[14] ? _GEN5297 : _GEN5296;
wire  _GEN5299 = io_x[10] ? _GEN5298 : _GEN5295;
wire  _GEN5300 = io_x[23] ? _GEN5299 : _GEN5292;
wire  _GEN5301 = io_x[16] ? _GEN5300 : _GEN5285;
wire  _GEN5302 = io_x[12] ? _GEN5301 : _GEN5274;
wire  _GEN5303 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5304 = io_x[14] ? _GEN5303 : _GEN3708;
wire  _GEN5305 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5306 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5307 = io_x[14] ? _GEN5306 : _GEN5305;
wire  _GEN5308 = io_x[10] ? _GEN5307 : _GEN5304;
wire  _GEN5309 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5310 = io_x[14] ? _GEN3709 : _GEN5309;
wire  _GEN5311 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5312 = io_x[14] ? _GEN5311 : _GEN3709;
wire  _GEN5313 = io_x[10] ? _GEN5312 : _GEN5310;
wire  _GEN5314 = io_x[23] ? _GEN5313 : _GEN5308;
wire  _GEN5315 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5316 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5317 = io_x[14] ? _GEN5316 : _GEN5315;
wire  _GEN5318 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5319 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5320 = io_x[14] ? _GEN5319 : _GEN5318;
wire  _GEN5321 = io_x[10] ? _GEN5320 : _GEN5317;
wire  _GEN5322 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5323 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5324 = io_x[14] ? _GEN5323 : _GEN5322;
wire  _GEN5325 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5326 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5327 = io_x[14] ? _GEN5326 : _GEN5325;
wire  _GEN5328 = io_x[10] ? _GEN5327 : _GEN5324;
wire  _GEN5329 = io_x[23] ? _GEN5328 : _GEN5321;
wire  _GEN5330 = io_x[16] ? _GEN5329 : _GEN5314;
wire  _GEN5331 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5332 = io_x[14] ? _GEN5331 : _GEN3709;
wire  _GEN5333 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5334 = io_x[14] ? _GEN5333 : _GEN3709;
wire  _GEN5335 = io_x[10] ? _GEN5334 : _GEN5332;
wire  _GEN5336 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5337 = io_x[14] ? _GEN5336 : _GEN3709;
wire  _GEN5338 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5339 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5340 = io_x[14] ? _GEN5339 : _GEN5338;
wire  _GEN5341 = io_x[10] ? _GEN5340 : _GEN5337;
wire  _GEN5342 = io_x[23] ? _GEN5341 : _GEN5335;
wire  _GEN5343 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5344 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5345 = io_x[14] ? _GEN5344 : _GEN5343;
wire  _GEN5346 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5347 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5348 = io_x[14] ? _GEN5347 : _GEN5346;
wire  _GEN5349 = io_x[10] ? _GEN5348 : _GEN5345;
wire  _GEN5350 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5351 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5352 = io_x[14] ? _GEN5351 : _GEN5350;
wire  _GEN5353 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5354 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5355 = io_x[14] ? _GEN5354 : _GEN5353;
wire  _GEN5356 = io_x[10] ? _GEN5355 : _GEN5352;
wire  _GEN5357 = io_x[23] ? _GEN5356 : _GEN5349;
wire  _GEN5358 = io_x[16] ? _GEN5357 : _GEN5342;
wire  _GEN5359 = io_x[12] ? _GEN5358 : _GEN5330;
wire  _GEN5360 = io_x[2] ? _GEN5359 : _GEN5302;
wire  _GEN5361 = io_x[9] ? _GEN5360 : _GEN5247;
wire  _GEN5362 = io_x[13] ? _GEN5361 : _GEN5171;
wire  _GEN5363 = io_x[7] ? _GEN5362 : _GEN5037;
wire  _GEN5364 = io_x[15] ? _GEN5363 : _GEN4811;
wire  _GEN5365 = io_x[3] ? _GEN5364 : _GEN4411;
wire  _GEN5366 = io_x[23] ? _GEN3713 : _GEN3741;
wire  _GEN5367 = io_x[16] ? _GEN5366 : _GEN3707;
wire  _GEN5368 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5369 = io_x[14] ? _GEN5368 : _GEN3709;
wire  _GEN5370 = io_x[10] ? _GEN5369 : _GEN3711;
wire  _GEN5371 = io_x[23] ? _GEN5370 : _GEN3741;
wire  _GEN5372 = io_x[16] ? _GEN5371 : _GEN3727;
wire  _GEN5373 = io_x[12] ? _GEN5372 : _GEN5367;
wire  _GEN5374 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN5375 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5376 = io_x[14] ? _GEN5375 : _GEN3709;
wire  _GEN5377 = io_x[10] ? _GEN5376 : _GEN3711;
wire  _GEN5378 = io_x[23] ? _GEN5377 : _GEN5374;
wire  _GEN5379 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5380 = io_x[10] ? _GEN3716 : _GEN5379;
wire  _GEN5381 = io_x[23] ? _GEN5380 : _GEN3713;
wire  _GEN5382 = io_x[16] ? _GEN5381 : _GEN5378;
wire  _GEN5383 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5384 = io_x[14] ? _GEN5383 : _GEN3709;
wire  _GEN5385 = io_x[10] ? _GEN5384 : _GEN3711;
wire  _GEN5386 = io_x[23] ? _GEN3713 : _GEN5385;
wire  _GEN5387 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5388 = io_x[14] ? _GEN5387 : _GEN3709;
wire  _GEN5389 = io_x[10] ? _GEN5388 : _GEN3716;
wire  _GEN5390 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN5391 = io_x[23] ? _GEN5390 : _GEN5389;
wire  _GEN5392 = io_x[16] ? _GEN5391 : _GEN5386;
wire  _GEN5393 = io_x[12] ? _GEN5392 : _GEN5382;
wire  _GEN5394 = io_x[2] ? _GEN5393 : _GEN5373;
wire  _GEN5395 = io_x[23] ? _GEN3741 : _GEN3713;
wire  _GEN5396 = io_x[16] ? _GEN3707 : _GEN5395;
wire  _GEN5397 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5398 = io_x[10] ? _GEN5397 : _GEN3716;
wire  _GEN5399 = io_x[23] ? _GEN5398 : _GEN3713;
wire  _GEN5400 = io_x[16] ? _GEN5399 : _GEN3727;
wire  _GEN5401 = io_x[12] ? _GEN5400 : _GEN5396;
wire  _GEN5402 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN5403 = io_x[23] ? _GEN3741 : _GEN5402;
wire  _GEN5404 = io_x[16] ? _GEN3727 : _GEN5403;
wire  _GEN5405 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5406 = io_x[14] ? _GEN3709 : _GEN5405;
wire  _GEN5407 = io_x[10] ? _GEN5406 : _GEN3716;
wire  _GEN5408 = io_x[23] ? _GEN3741 : _GEN5407;
wire  _GEN5409 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5410 = io_x[14] ? _GEN5409 : _GEN3709;
wire  _GEN5411 = io_x[10] ? _GEN5410 : _GEN3711;
wire  _GEN5412 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5413 = io_x[14] ? _GEN5412 : _GEN3709;
wire  _GEN5414 = io_x[10] ? _GEN5413 : _GEN3716;
wire  _GEN5415 = io_x[23] ? _GEN5414 : _GEN5411;
wire  _GEN5416 = io_x[16] ? _GEN5415 : _GEN5408;
wire  _GEN5417 = io_x[12] ? _GEN5416 : _GEN5404;
wire  _GEN5418 = io_x[2] ? _GEN5417 : _GEN5401;
wire  _GEN5419 = io_x[9] ? _GEN5418 : _GEN5394;
wire  _GEN5420 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5421 = io_x[14] ? _GEN5420 : _GEN3709;
wire  _GEN5422 = io_x[10] ? _GEN3711 : _GEN5421;
wire  _GEN5423 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN5424 = io_x[23] ? _GEN5423 : _GEN5422;
wire  _GEN5425 = io_x[16] ? _GEN5424 : _GEN3707;
wire  _GEN5426 = io_x[12] ? _GEN4478 : _GEN5425;
wire  _GEN5427 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5428 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5429 = io_x[14] ? _GEN5428 : _GEN3708;
wire  _GEN5430 = io_x[10] ? _GEN5429 : _GEN5427;
wire  _GEN5431 = io_x[23] ? _GEN3741 : _GEN5430;
wire  _GEN5432 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5433 = io_x[10] ? _GEN5432 : _GEN3711;
wire  _GEN5434 = io_x[23] ? _GEN5433 : _GEN3741;
wire  _GEN5435 = io_x[16] ? _GEN5434 : _GEN5431;
wire  _GEN5436 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5437 = io_x[10] ? _GEN5436 : _GEN3711;
wire  _GEN5438 = io_x[23] ? _GEN3713 : _GEN5437;
wire  _GEN5439 = io_x[16] ? _GEN3707 : _GEN5438;
wire  _GEN5440 = io_x[12] ? _GEN5439 : _GEN5435;
wire  _GEN5441 = io_x[2] ? _GEN5440 : _GEN5426;
wire  _GEN5442 = io_x[23] ? _GEN3741 : _GEN3713;
wire  _GEN5443 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN5444 = io_x[23] ? _GEN3713 : _GEN5443;
wire  _GEN5445 = io_x[16] ? _GEN5444 : _GEN5442;
wire  _GEN5446 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN5447 = io_x[23] ? _GEN3713 : _GEN5446;
wire  _GEN5448 = io_x[16] ? _GEN5447 : _GEN3707;
wire  _GEN5449 = io_x[12] ? _GEN5448 : _GEN5445;
wire  _GEN5450 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5451 = io_x[14] ? _GEN3709 : _GEN5450;
wire  _GEN5452 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5453 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5454 = io_x[14] ? _GEN5453 : _GEN5452;
wire  _GEN5455 = io_x[10] ? _GEN5454 : _GEN5451;
wire  _GEN5456 = io_x[23] ? _GEN3741 : _GEN5455;
wire  _GEN5457 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5458 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5459 = io_x[14] ? _GEN3709 : _GEN5458;
wire  _GEN5460 = io_x[10] ? _GEN5459 : _GEN5457;
wire  _GEN5461 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5462 = io_x[14] ? _GEN3709 : _GEN5461;
wire  _GEN5463 = io_x[10] ? _GEN5462 : _GEN3716;
wire  _GEN5464 = io_x[23] ? _GEN5463 : _GEN5460;
wire  _GEN5465 = io_x[16] ? _GEN5464 : _GEN5456;
wire  _GEN5466 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN5467 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN5468 = io_x[23] ? _GEN5467 : _GEN5466;
wire  _GEN5469 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5470 = io_x[10] ? _GEN5469 : _GEN3716;
wire  _GEN5471 = io_x[23] ? _GEN5470 : _GEN3741;
wire  _GEN5472 = io_x[16] ? _GEN5471 : _GEN5468;
wire  _GEN5473 = io_x[12] ? _GEN5472 : _GEN5465;
wire  _GEN5474 = io_x[2] ? _GEN5473 : _GEN5449;
wire  _GEN5475 = io_x[9] ? _GEN5474 : _GEN5441;
wire  _GEN5476 = io_x[13] ? _GEN5475 : _GEN5419;
wire  _GEN5477 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5478 = io_x[14] ? _GEN5477 : _GEN3709;
wire  _GEN5479 = io_x[10] ? _GEN5478 : _GEN3711;
wire  _GEN5480 = io_x[23] ? _GEN3741 : _GEN5479;
wire  _GEN5481 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5482 = io_x[10] ? _GEN5481 : _GEN3716;
wire  _GEN5483 = io_x[23] ? _GEN3713 : _GEN5482;
wire  _GEN5484 = io_x[16] ? _GEN5483 : _GEN5480;
wire  _GEN5485 = io_x[12] ? _GEN5484 : _GEN3893;
wire  _GEN5486 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5487 = io_x[14] ? _GEN5486 : _GEN3708;
wire  _GEN5488 = io_x[10] ? _GEN3716 : _GEN5487;
wire  _GEN5489 = io_x[23] ? _GEN3713 : _GEN5488;
wire  _GEN5490 = io_x[16] ? _GEN5489 : _GEN3727;
wire  _GEN5491 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5492 = io_x[14] ? _GEN5491 : _GEN3709;
wire  _GEN5493 = io_x[10] ? _GEN5492 : _GEN3711;
wire  _GEN5494 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5495 = io_x[14] ? _GEN5494 : _GEN3709;
wire  _GEN5496 = io_x[10] ? _GEN5495 : _GEN3711;
wire  _GEN5497 = io_x[23] ? _GEN5496 : _GEN5493;
wire  _GEN5498 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5499 = io_x[14] ? _GEN5498 : _GEN3709;
wire  _GEN5500 = io_x[10] ? _GEN5499 : _GEN3716;
wire  _GEN5501 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5502 = io_x[14] ? _GEN5501 : _GEN3709;
wire  _GEN5503 = io_x[10] ? _GEN5502 : _GEN3711;
wire  _GEN5504 = io_x[23] ? _GEN5503 : _GEN5500;
wire  _GEN5505 = io_x[16] ? _GEN5504 : _GEN5497;
wire  _GEN5506 = io_x[12] ? _GEN5505 : _GEN5490;
wire  _GEN5507 = io_x[2] ? _GEN5506 : _GEN5485;
wire  _GEN5508 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5509 = io_x[10] ? _GEN3716 : _GEN5508;
wire  _GEN5510 = io_x[23] ? _GEN5509 : _GEN3741;
wire  _GEN5511 = io_x[16] ? _GEN5510 : _GEN3727;
wire  _GEN5512 = io_x[12] ? _GEN5511 : _GEN4478;
wire  _GEN5513 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5514 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5515 = io_x[14] ? _GEN5514 : _GEN3709;
wire  _GEN5516 = io_x[10] ? _GEN5515 : _GEN5513;
wire  _GEN5517 = io_x[23] ? _GEN3713 : _GEN5516;
wire  _GEN5518 = io_x[16] ? _GEN3707 : _GEN5517;
wire  _GEN5519 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5520 = io_x[14] ? _GEN5519 : _GEN3708;
wire  _GEN5521 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5522 = io_x[14] ? _GEN5521 : _GEN3709;
wire  _GEN5523 = io_x[10] ? _GEN5522 : _GEN5520;
wire  _GEN5524 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5525 = io_x[14] ? _GEN5524 : _GEN3709;
wire  _GEN5526 = io_x[10] ? _GEN3711 : _GEN5525;
wire  _GEN5527 = io_x[23] ? _GEN5526 : _GEN5523;
wire  _GEN5528 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5529 = io_x[14] ? _GEN5528 : _GEN3708;
wire  _GEN5530 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5531 = io_x[14] ? _GEN5530 : _GEN3709;
wire  _GEN5532 = io_x[10] ? _GEN5531 : _GEN5529;
wire  _GEN5533 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5534 = io_x[14] ? _GEN5533 : _GEN3708;
wire  _GEN5535 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5536 = io_x[14] ? _GEN5535 : _GEN3709;
wire  _GEN5537 = io_x[10] ? _GEN5536 : _GEN5534;
wire  _GEN5538 = io_x[23] ? _GEN5537 : _GEN5532;
wire  _GEN5539 = io_x[16] ? _GEN5538 : _GEN5527;
wire  _GEN5540 = io_x[12] ? _GEN5539 : _GEN5518;
wire  _GEN5541 = io_x[2] ? _GEN5540 : _GEN5512;
wire  _GEN5542 = io_x[9] ? _GEN5541 : _GEN5507;
wire  _GEN5543 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5544 = io_x[14] ? _GEN3709 : _GEN5543;
wire  _GEN5545 = io_x[10] ? _GEN5544 : _GEN3711;
wire  _GEN5546 = io_x[23] ? _GEN3713 : _GEN5545;
wire  _GEN5547 = io_x[16] ? _GEN3727 : _GEN5546;
wire  _GEN5548 = io_x[12] ? _GEN3893 : _GEN5547;
wire  _GEN5549 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5550 = io_x[14] ? _GEN3709 : _GEN5549;
wire  _GEN5551 = io_x[10] ? _GEN5550 : _GEN3711;
wire  _GEN5552 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5553 = io_x[10] ? _GEN5552 : _GEN3711;
wire  _GEN5554 = io_x[23] ? _GEN5553 : _GEN5551;
wire  _GEN5555 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5556 = io_x[14] ? _GEN3709 : _GEN5555;
wire  _GEN5557 = io_x[10] ? _GEN5556 : _GEN3711;
wire  _GEN5558 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5559 = io_x[14] ? _GEN3709 : _GEN5558;
wire  _GEN5560 = io_x[10] ? _GEN5559 : _GEN3711;
wire  _GEN5561 = io_x[23] ? _GEN5560 : _GEN5557;
wire  _GEN5562 = io_x[16] ? _GEN5561 : _GEN5554;
wire  _GEN5563 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5564 = io_x[14] ? _GEN5563 : _GEN3709;
wire  _GEN5565 = io_x[10] ? _GEN3716 : _GEN5564;
wire  _GEN5566 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5567 = io_x[14] ? _GEN3708 : _GEN5566;
wire  _GEN5568 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5569 = io_x[14] ? _GEN5568 : _GEN3709;
wire  _GEN5570 = io_x[10] ? _GEN5569 : _GEN5567;
wire  _GEN5571 = io_x[23] ? _GEN5570 : _GEN5565;
wire  _GEN5572 = io_x[16] ? _GEN3727 : _GEN5571;
wire  _GEN5573 = io_x[12] ? _GEN5572 : _GEN5562;
wire  _GEN5574 = io_x[2] ? _GEN5573 : _GEN5548;
wire  _GEN5575 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5576 = io_x[14] ? _GEN5575 : _GEN3709;
wire  _GEN5577 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5578 = io_x[14] ? _GEN5577 : _GEN3709;
wire  _GEN5579 = io_x[10] ? _GEN5578 : _GEN5576;
wire  _GEN5580 = io_x[23] ? _GEN3741 : _GEN5579;
wire  _GEN5581 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5582 = io_x[14] ? _GEN5581 : _GEN3709;
wire  _GEN5583 = io_x[10] ? _GEN3711 : _GEN5582;
wire  _GEN5584 = io_x[23] ? _GEN3741 : _GEN5583;
wire  _GEN5585 = io_x[16] ? _GEN5584 : _GEN5580;
wire  _GEN5586 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5587 = io_x[10] ? _GEN3711 : _GEN5586;
wire  _GEN5588 = io_x[23] ? _GEN3741 : _GEN5587;
wire  _GEN5589 = io_x[16] ? _GEN5588 : _GEN3707;
wire  _GEN5590 = io_x[12] ? _GEN5589 : _GEN5585;
wire  _GEN5591 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5592 = io_x[10] ? _GEN3711 : _GEN5591;
wire  _GEN5593 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5594 = io_x[14] ? _GEN5593 : _GEN3709;
wire  _GEN5595 = io_x[10] ? _GEN3711 : _GEN5594;
wire  _GEN5596 = io_x[23] ? _GEN5595 : _GEN5592;
wire  _GEN5597 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5598 = io_x[14] ? _GEN5597 : _GEN3709;
wire  _GEN5599 = io_x[10] ? _GEN3711 : _GEN5598;
wire  _GEN5600 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5601 = io_x[14] ? _GEN5600 : _GEN3709;
wire  _GEN5602 = io_x[10] ? _GEN3711 : _GEN5601;
wire  _GEN5603 = io_x[23] ? _GEN5602 : _GEN5599;
wire  _GEN5604 = io_x[16] ? _GEN5603 : _GEN5596;
wire  _GEN5605 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5606 = io_x[14] ? _GEN5605 : _GEN3708;
wire  _GEN5607 = io_x[10] ? _GEN5606 : _GEN3716;
wire  _GEN5608 = io_x[23] ? _GEN3741 : _GEN5607;
wire  _GEN5609 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5610 = io_x[14] ? _GEN5609 : _GEN3709;
wire  _GEN5611 = io_x[10] ? _GEN5610 : _GEN3716;
wire  _GEN5612 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5613 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5614 = io_x[14] ? _GEN5613 : _GEN3709;
wire  _GEN5615 = io_x[10] ? _GEN5614 : _GEN5612;
wire  _GEN5616 = io_x[23] ? _GEN5615 : _GEN5611;
wire  _GEN5617 = io_x[16] ? _GEN5616 : _GEN5608;
wire  _GEN5618 = io_x[12] ? _GEN5617 : _GEN5604;
wire  _GEN5619 = io_x[2] ? _GEN5618 : _GEN5590;
wire  _GEN5620 = io_x[9] ? _GEN5619 : _GEN5574;
wire  _GEN5621 = io_x[13] ? _GEN5620 : _GEN5542;
wire  _GEN5622 = io_x[7] ? _GEN5621 : _GEN5476;
wire  _GEN5623 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5624 = io_x[14] ? _GEN3709 : _GEN5623;
wire  _GEN5625 = io_x[10] ? _GEN5624 : _GEN3711;
wire  _GEN5626 = io_x[23] ? _GEN5625 : _GEN3713;
wire  _GEN5627 = io_x[16] ? _GEN5626 : _GEN3707;
wire  _GEN5628 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5629 = io_x[10] ? _GEN5628 : _GEN3711;
wire  _GEN5630 = io_x[23] ? _GEN3713 : _GEN5629;
wire  _GEN5631 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5632 = io_x[10] ? _GEN5631 : _GEN3711;
wire  _GEN5633 = io_x[23] ? _GEN3713 : _GEN5632;
wire  _GEN5634 = io_x[16] ? _GEN5633 : _GEN5630;
wire  _GEN5635 = io_x[12] ? _GEN5634 : _GEN5627;
wire  _GEN5636 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5637 = io_x[10] ? _GEN5636 : _GEN3711;
wire  _GEN5638 = io_x[23] ? _GEN3713 : _GEN5637;
wire  _GEN5639 = io_x[16] ? _GEN3707 : _GEN5638;
wire  _GEN5640 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5641 = io_x[14] ? _GEN5640 : _GEN3708;
wire  _GEN5642 = io_x[10] ? _GEN5641 : _GEN3711;
wire  _GEN5643 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5644 = io_x[14] ? _GEN5643 : _GEN3708;
wire  _GEN5645 = io_x[10] ? _GEN5644 : _GEN3711;
wire  _GEN5646 = io_x[23] ? _GEN5645 : _GEN5642;
wire  _GEN5647 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5648 = io_x[14] ? _GEN5647 : _GEN3708;
wire  _GEN5649 = io_x[10] ? _GEN5648 : _GEN3711;
wire  _GEN5650 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5651 = io_x[10] ? _GEN5650 : _GEN3711;
wire  _GEN5652 = io_x[23] ? _GEN5651 : _GEN5649;
wire  _GEN5653 = io_x[16] ? _GEN5652 : _GEN5646;
wire  _GEN5654 = io_x[12] ? _GEN5653 : _GEN5639;
wire  _GEN5655 = io_x[2] ? _GEN5654 : _GEN5635;
wire  _GEN5656 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5657 = io_x[14] ? _GEN5656 : _GEN3709;
wire  _GEN5658 = io_x[10] ? _GEN5657 : _GEN3711;
wire  _GEN5659 = io_x[23] ? _GEN5658 : _GEN3713;
wire  _GEN5660 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5661 = io_x[10] ? _GEN5660 : _GEN3711;
wire  _GEN5662 = io_x[23] ? _GEN5661 : _GEN3713;
wire  _GEN5663 = io_x[16] ? _GEN5662 : _GEN5659;
wire  _GEN5664 = io_x[12] ? _GEN4478 : _GEN5663;
wire  _GEN5665 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5666 = io_x[14] ? _GEN5665 : _GEN3708;
wire  _GEN5667 = io_x[10] ? _GEN3711 : _GEN5666;
wire  _GEN5668 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5669 = io_x[14] ? _GEN5668 : _GEN3709;
wire  _GEN5670 = io_x[10] ? _GEN3711 : _GEN5669;
wire  _GEN5671 = io_x[23] ? _GEN5670 : _GEN5667;
wire  _GEN5672 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN5673 = io_x[23] ? _GEN3713 : _GEN5672;
wire  _GEN5674 = io_x[16] ? _GEN5673 : _GEN5671;
wire  _GEN5675 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5676 = io_x[14] ? _GEN3708 : _GEN5675;
wire  _GEN5677 = io_x[10] ? _GEN3716 : _GEN5676;
wire  _GEN5678 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5679 = io_x[14] ? _GEN3708 : _GEN5678;
wire  _GEN5680 = io_x[10] ? _GEN3711 : _GEN5679;
wire  _GEN5681 = io_x[23] ? _GEN5680 : _GEN5677;
wire  _GEN5682 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5683 = io_x[14] ? _GEN5682 : _GEN3708;
wire  _GEN5684 = io_x[10] ? _GEN5683 : _GEN3711;
wire  _GEN5685 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5686 = io_x[14] ? _GEN5685 : _GEN3709;
wire  _GEN5687 = io_x[10] ? _GEN5686 : _GEN3711;
wire  _GEN5688 = io_x[23] ? _GEN5687 : _GEN5684;
wire  _GEN5689 = io_x[16] ? _GEN5688 : _GEN5681;
wire  _GEN5690 = io_x[12] ? _GEN5689 : _GEN5674;
wire  _GEN5691 = io_x[2] ? _GEN5690 : _GEN5664;
wire  _GEN5692 = io_x[9] ? _GEN5691 : _GEN5655;
wire  _GEN5693 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5694 = io_x[10] ? _GEN5693 : _GEN3711;
wire  _GEN5695 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5696 = io_x[14] ? _GEN5695 : _GEN3709;
wire  _GEN5697 = io_x[10] ? _GEN5696 : _GEN3711;
wire  _GEN5698 = io_x[23] ? _GEN5697 : _GEN5694;
wire  _GEN5699 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5700 = io_x[10] ? _GEN5699 : _GEN3716;
wire  _GEN5701 = io_x[23] ? _GEN3713 : _GEN5700;
wire  _GEN5702 = io_x[16] ? _GEN5701 : _GEN5698;
wire  _GEN5703 = io_x[23] ? _GEN3741 : _GEN3713;
wire  _GEN5704 = io_x[16] ? _GEN3707 : _GEN5703;
wire  _GEN5705 = io_x[12] ? _GEN5704 : _GEN5702;
wire  _GEN5706 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5707 = io_x[10] ? _GEN5706 : _GEN3711;
wire  _GEN5708 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5709 = io_x[14] ? _GEN5708 : _GEN3709;
wire  _GEN5710 = io_x[10] ? _GEN5709 : _GEN3711;
wire  _GEN5711 = io_x[23] ? _GEN5710 : _GEN5707;
wire  _GEN5712 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5713 = io_x[14] ? _GEN5712 : _GEN3709;
wire  _GEN5714 = io_x[10] ? _GEN3711 : _GEN5713;
wire  _GEN5715 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5716 = io_x[10] ? _GEN5715 : _GEN3711;
wire  _GEN5717 = io_x[23] ? _GEN5716 : _GEN5714;
wire  _GEN5718 = io_x[16] ? _GEN5717 : _GEN5711;
wire  _GEN5719 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5720 = io_x[14] ? _GEN3708 : _GEN5719;
wire  _GEN5721 = io_x[10] ? _GEN3716 : _GEN5720;
wire  _GEN5722 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN5723 = io_x[23] ? _GEN5722 : _GEN5721;
wire  _GEN5724 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5725 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5726 = io_x[14] ? _GEN5725 : _GEN5724;
wire  _GEN5727 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5728 = io_x[10] ? _GEN5727 : _GEN5726;
wire  _GEN5729 = io_x[23] ? _GEN3741 : _GEN5728;
wire  _GEN5730 = io_x[16] ? _GEN5729 : _GEN5723;
wire  _GEN5731 = io_x[12] ? _GEN5730 : _GEN5718;
wire  _GEN5732 = io_x[2] ? _GEN5731 : _GEN5705;
wire  _GEN5733 = io_x[23] ? _GEN3741 : _GEN3713;
wire  _GEN5734 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5735 = io_x[14] ? _GEN5734 : _GEN3709;
wire  _GEN5736 = io_x[10] ? _GEN5735 : _GEN3711;
wire  _GEN5737 = io_x[23] ? _GEN3713 : _GEN5736;
wire  _GEN5738 = io_x[16] ? _GEN5737 : _GEN5733;
wire  _GEN5739 = io_x[23] ? _GEN3713 : _GEN3741;
wire  _GEN5740 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5741 = io_x[14] ? _GEN5740 : _GEN3708;
wire  _GEN5742 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5743 = io_x[14] ? _GEN5742 : _GEN3709;
wire  _GEN5744 = io_x[10] ? _GEN5743 : _GEN5741;
wire  _GEN5745 = io_x[23] ? _GEN5744 : _GEN3741;
wire  _GEN5746 = io_x[16] ? _GEN5745 : _GEN5739;
wire  _GEN5747 = io_x[12] ? _GEN5746 : _GEN5738;
wire  _GEN5748 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5749 = io_x[14] ? _GEN3708 : _GEN5748;
wire  _GEN5750 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5751 = io_x[14] ? _GEN5750 : _GEN3709;
wire  _GEN5752 = io_x[10] ? _GEN5751 : _GEN5749;
wire  _GEN5753 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5754 = io_x[14] ? _GEN3709 : _GEN5753;
wire  _GEN5755 = io_x[10] ? _GEN3711 : _GEN5754;
wire  _GEN5756 = io_x[23] ? _GEN5755 : _GEN5752;
wire  _GEN5757 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5758 = io_x[14] ? _GEN5757 : _GEN3709;
wire  _GEN5759 = io_x[10] ? _GEN5758 : _GEN3711;
wire  _GEN5760 = io_x[23] ? _GEN3741 : _GEN5759;
wire  _GEN5761 = io_x[16] ? _GEN5760 : _GEN5756;
wire  _GEN5762 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5763 = io_x[10] ? _GEN3711 : _GEN5762;
wire  _GEN5764 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5765 = io_x[14] ? _GEN5764 : _GEN3708;
wire  _GEN5766 = io_x[10] ? _GEN5765 : _GEN3711;
wire  _GEN5767 = io_x[23] ? _GEN5766 : _GEN5763;
wire  _GEN5768 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5769 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5770 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5771 = io_x[14] ? _GEN5770 : _GEN5769;
wire  _GEN5772 = io_x[10] ? _GEN5771 : _GEN5768;
wire  _GEN5773 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN5774 = io_x[23] ? _GEN5773 : _GEN5772;
wire  _GEN5775 = io_x[16] ? _GEN5774 : _GEN5767;
wire  _GEN5776 = io_x[12] ? _GEN5775 : _GEN5761;
wire  _GEN5777 = io_x[2] ? _GEN5776 : _GEN5747;
wire  _GEN5778 = io_x[9] ? _GEN5777 : _GEN5732;
wire  _GEN5779 = io_x[13] ? _GEN5778 : _GEN5692;
wire  _GEN5780 = io_x[16] ? _GEN3727 : _GEN3707;
wire  _GEN5781 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN5782 = io_x[23] ? _GEN3741 : _GEN5781;
wire  _GEN5783 = io_x[16] ? _GEN3707 : _GEN5782;
wire  _GEN5784 = io_x[12] ? _GEN5783 : _GEN5780;
wire  _GEN5785 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN5786 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5787 = io_x[10] ? _GEN3716 : _GEN5786;
wire  _GEN5788 = io_x[23] ? _GEN5787 : _GEN5785;
wire  _GEN5789 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5790 = io_x[10] ? _GEN3711 : _GEN5789;
wire  _GEN5791 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5792 = io_x[14] ? _GEN5791 : _GEN3708;
wire  _GEN5793 = io_x[10] ? _GEN5792 : _GEN3711;
wire  _GEN5794 = io_x[23] ? _GEN5793 : _GEN5790;
wire  _GEN5795 = io_x[16] ? _GEN5794 : _GEN5788;
wire  _GEN5796 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5797 = io_x[14] ? _GEN5796 : _GEN3709;
wire  _GEN5798 = io_x[10] ? _GEN5797 : _GEN3711;
wire  _GEN5799 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5800 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5801 = io_x[14] ? _GEN5800 : _GEN5799;
wire  _GEN5802 = io_x[10] ? _GEN5801 : _GEN3716;
wire  _GEN5803 = io_x[23] ? _GEN5802 : _GEN5798;
wire  _GEN5804 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5805 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5806 = io_x[14] ? _GEN5805 : _GEN5804;
wire  _GEN5807 = io_x[10] ? _GEN5806 : _GEN3711;
wire  _GEN5808 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5809 = io_x[14] ? _GEN5808 : _GEN3708;
wire  _GEN5810 = io_x[10] ? _GEN5809 : _GEN3711;
wire  _GEN5811 = io_x[23] ? _GEN5810 : _GEN5807;
wire  _GEN5812 = io_x[16] ? _GEN5811 : _GEN5803;
wire  _GEN5813 = io_x[12] ? _GEN5812 : _GEN5795;
wire  _GEN5814 = io_x[2] ? _GEN5813 : _GEN5784;
wire  _GEN5815 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5816 = io_x[10] ? _GEN5815 : _GEN3716;
wire  _GEN5817 = io_x[23] ? _GEN3741 : _GEN5816;
wire  _GEN5818 = io_x[16] ? _GEN5817 : _GEN3727;
wire  _GEN5819 = io_x[12] ? _GEN5818 : _GEN3893;
wire  _GEN5820 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN5821 = io_x[23] ? _GEN3713 : _GEN5820;
wire  _GEN5822 = io_x[16] ? _GEN3707 : _GEN5821;
wire  _GEN5823 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5824 = io_x[10] ? _GEN5823 : _GEN3711;
wire  _GEN5825 = io_x[23] ? _GEN3713 : _GEN5824;
wire  _GEN5826 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5827 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5828 = io_x[14] ? _GEN5827 : _GEN5826;
wire  _GEN5829 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5830 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5831 = io_x[14] ? _GEN5830 : _GEN5829;
wire  _GEN5832 = io_x[10] ? _GEN5831 : _GEN5828;
wire  _GEN5833 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5834 = io_x[14] ? _GEN5833 : _GEN3709;
wire  _GEN5835 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5836 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5837 = io_x[14] ? _GEN5836 : _GEN5835;
wire  _GEN5838 = io_x[10] ? _GEN5837 : _GEN5834;
wire  _GEN5839 = io_x[23] ? _GEN5838 : _GEN5832;
wire  _GEN5840 = io_x[16] ? _GEN5839 : _GEN5825;
wire  _GEN5841 = io_x[12] ? _GEN5840 : _GEN5822;
wire  _GEN5842 = io_x[2] ? _GEN5841 : _GEN5819;
wire  _GEN5843 = io_x[9] ? _GEN5842 : _GEN5814;
wire  _GEN5844 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5845 = io_x[14] ? _GEN5844 : _GEN3708;
wire  _GEN5846 = io_x[10] ? _GEN5845 : _GEN3711;
wire  _GEN5847 = io_x[23] ? _GEN5846 : _GEN3713;
wire  _GEN5848 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5849 = io_x[14] ? _GEN5848 : _GEN3708;
wire  _GEN5850 = io_x[10] ? _GEN5849 : _GEN3711;
wire  _GEN5851 = io_x[23] ? _GEN3713 : _GEN5850;
wire  _GEN5852 = io_x[16] ? _GEN5851 : _GEN5847;
wire  _GEN5853 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5854 = io_x[10] ? _GEN5853 : _GEN3711;
wire  _GEN5855 = io_x[23] ? _GEN3713 : _GEN5854;
wire  _GEN5856 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5857 = io_x[14] ? _GEN3709 : _GEN5856;
wire  _GEN5858 = io_x[10] ? _GEN5857 : _GEN3711;
wire  _GEN5859 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5860 = io_x[14] ? _GEN3708 : _GEN5859;
wire  _GEN5861 = io_x[10] ? _GEN5860 : _GEN3716;
wire  _GEN5862 = io_x[23] ? _GEN5861 : _GEN5858;
wire  _GEN5863 = io_x[16] ? _GEN5862 : _GEN5855;
wire  _GEN5864 = io_x[12] ? _GEN5863 : _GEN5852;
wire  _GEN5865 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5866 = io_x[10] ? _GEN5865 : _GEN3711;
wire  _GEN5867 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN5868 = io_x[23] ? _GEN5867 : _GEN5866;
wire  _GEN5869 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5870 = io_x[14] ? _GEN5869 : _GEN3709;
wire  _GEN5871 = io_x[10] ? _GEN5870 : _GEN3716;
wire  _GEN5872 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5873 = io_x[14] ? _GEN5872 : _GEN3708;
wire  _GEN5874 = io_x[10] ? _GEN5873 : _GEN3711;
wire  _GEN5875 = io_x[23] ? _GEN5874 : _GEN5871;
wire  _GEN5876 = io_x[16] ? _GEN5875 : _GEN5868;
wire  _GEN5877 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5878 = io_x[14] ? _GEN3708 : _GEN5877;
wire  _GEN5879 = io_x[10] ? _GEN5878 : _GEN3711;
wire  _GEN5880 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5881 = io_x[14] ? _GEN3708 : _GEN5880;
wire  _GEN5882 = io_x[10] ? _GEN5881 : _GEN3711;
wire  _GEN5883 = io_x[23] ? _GEN5882 : _GEN5879;
wire  _GEN5884 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5885 = io_x[14] ? _GEN3709 : _GEN5884;
wire  _GEN5886 = io_x[10] ? _GEN5885 : _GEN3711;
wire  _GEN5887 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5888 = io_x[14] ? _GEN3709 : _GEN5887;
wire  _GEN5889 = io_x[10] ? _GEN5888 : _GEN3711;
wire  _GEN5890 = io_x[23] ? _GEN5889 : _GEN5886;
wire  _GEN5891 = io_x[16] ? _GEN5890 : _GEN5883;
wire  _GEN5892 = io_x[12] ? _GEN5891 : _GEN5876;
wire  _GEN5893 = io_x[2] ? _GEN5892 : _GEN5864;
wire  _GEN5894 = io_x[23] ? _GEN3741 : _GEN3713;
wire  _GEN5895 = io_x[23] ? _GEN3741 : _GEN3713;
wire  _GEN5896 = io_x[16] ? _GEN5895 : _GEN5894;
wire  _GEN5897 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5898 = io_x[14] ? _GEN5897 : _GEN3709;
wire  _GEN5899 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5900 = io_x[14] ? _GEN5899 : _GEN3709;
wire  _GEN5901 = io_x[10] ? _GEN5900 : _GEN5898;
wire  _GEN5902 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5903 = io_x[14] ? _GEN5902 : _GEN3709;
wire  _GEN5904 = io_x[10] ? _GEN5903 : _GEN3711;
wire  _GEN5905 = io_x[23] ? _GEN5904 : _GEN5901;
wire  _GEN5906 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5907 = io_x[14] ? _GEN5906 : _GEN3709;
wire  _GEN5908 = io_x[10] ? _GEN5907 : _GEN3711;
wire  _GEN5909 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5910 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5911 = io_x[14] ? _GEN5910 : _GEN3709;
wire  _GEN5912 = io_x[10] ? _GEN5911 : _GEN5909;
wire  _GEN5913 = io_x[23] ? _GEN5912 : _GEN5908;
wire  _GEN5914 = io_x[16] ? _GEN5913 : _GEN5905;
wire  _GEN5915 = io_x[12] ? _GEN5914 : _GEN5896;
wire  _GEN5916 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5917 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5918 = io_x[14] ? _GEN5917 : _GEN5916;
wire  _GEN5919 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5920 = io_x[10] ? _GEN5919 : _GEN5918;
wire  _GEN5921 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5922 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5923 = io_x[14] ? _GEN5922 : _GEN5921;
wire  _GEN5924 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5925 = io_x[10] ? _GEN5924 : _GEN5923;
wire  _GEN5926 = io_x[23] ? _GEN5925 : _GEN5920;
wire  _GEN5927 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5928 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5929 = io_x[14] ? _GEN5928 : _GEN5927;
wire  _GEN5930 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5931 = io_x[10] ? _GEN5930 : _GEN5929;
wire  _GEN5932 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5933 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5934 = io_x[14] ? _GEN5933 : _GEN5932;
wire  _GEN5935 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN5936 = io_x[10] ? _GEN5935 : _GEN5934;
wire  _GEN5937 = io_x[23] ? _GEN5936 : _GEN5931;
wire  _GEN5938 = io_x[16] ? _GEN5937 : _GEN5926;
wire  _GEN5939 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5940 = io_x[14] ? _GEN5939 : _GEN3708;
wire  _GEN5941 = io_x[10] ? _GEN5940 : _GEN3716;
wire  _GEN5942 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5943 = io_x[14] ? _GEN5942 : _GEN3709;
wire  _GEN5944 = io_x[10] ? _GEN5943 : _GEN3716;
wire  _GEN5945 = io_x[23] ? _GEN5944 : _GEN5941;
wire  _GEN5946 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5947 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5948 = io_x[14] ? _GEN5947 : _GEN5946;
wire  _GEN5949 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5950 = io_x[14] ? _GEN5949 : _GEN3709;
wire  _GEN5951 = io_x[10] ? _GEN5950 : _GEN5948;
wire  _GEN5952 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5953 = io_x[14] ? _GEN3708 : _GEN5952;
wire  _GEN5954 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5955 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5956 = io_x[14] ? _GEN5955 : _GEN5954;
wire  _GEN5957 = io_x[10] ? _GEN5956 : _GEN5953;
wire  _GEN5958 = io_x[23] ? _GEN5957 : _GEN5951;
wire  _GEN5959 = io_x[16] ? _GEN5958 : _GEN5945;
wire  _GEN5960 = io_x[12] ? _GEN5959 : _GEN5938;
wire  _GEN5961 = io_x[2] ? _GEN5960 : _GEN5915;
wire  _GEN5962 = io_x[9] ? _GEN5961 : _GEN5893;
wire  _GEN5963 = io_x[13] ? _GEN5962 : _GEN5843;
wire  _GEN5964 = io_x[7] ? _GEN5963 : _GEN5779;
wire  _GEN5965 = io_x[15] ? _GEN5964 : _GEN5622;
wire  _GEN5966 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN5967 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN5968 = io_x[23] ? _GEN5967 : _GEN5966;
wire  _GEN5969 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5970 = io_x[14] ? _GEN5969 : _GEN3708;
wire  _GEN5971 = io_x[10] ? _GEN3711 : _GEN5970;
wire  _GEN5972 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5973 = io_x[14] ? _GEN5972 : _GEN3709;
wire  _GEN5974 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN5975 = io_x[10] ? _GEN5974 : _GEN5973;
wire  _GEN5976 = io_x[23] ? _GEN5975 : _GEN5971;
wire  _GEN5977 = io_x[16] ? _GEN5976 : _GEN5968;
wire  _GEN5978 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN5979 = io_x[23] ? _GEN5978 : _GEN3741;
wire  _GEN5980 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5981 = io_x[14] ? _GEN5980 : _GEN3708;
wire  _GEN5982 = io_x[10] ? _GEN5981 : _GEN3711;
wire  _GEN5983 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN5984 = io_x[23] ? _GEN5983 : _GEN5982;
wire  _GEN5985 = io_x[16] ? _GEN5984 : _GEN5979;
wire  _GEN5986 = io_x[12] ? _GEN5985 : _GEN5977;
wire  _GEN5987 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5988 = io_x[14] ? _GEN5987 : _GEN3708;
wire  _GEN5989 = io_x[10] ? _GEN3711 : _GEN5988;
wire  _GEN5990 = io_x[23] ? _GEN3713 : _GEN5989;
wire  _GEN5991 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN5992 = io_x[14] ? _GEN5991 : _GEN3708;
wire  _GEN5993 = io_x[10] ? _GEN3711 : _GEN5992;
wire  _GEN5994 = io_x[23] ? _GEN3713 : _GEN5993;
wire  _GEN5995 = io_x[16] ? _GEN5994 : _GEN5990;
wire  _GEN5996 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN5997 = io_x[14] ? _GEN5996 : _GEN3709;
wire  _GEN5998 = io_x[10] ? _GEN5997 : _GEN3716;
wire  _GEN5999 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN6000 = io_x[23] ? _GEN5999 : _GEN5998;
wire  _GEN6001 = io_x[16] ? _GEN6000 : _GEN3707;
wire  _GEN6002 = io_x[12] ? _GEN6001 : _GEN5995;
wire  _GEN6003 = io_x[2] ? _GEN6002 : _GEN5986;
wire  _GEN6004 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6005 = io_x[10] ? _GEN6004 : _GEN3711;
wire  _GEN6006 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6007 = io_x[14] ? _GEN6006 : _GEN3709;
wire  _GEN6008 = io_x[10] ? _GEN6007 : _GEN3711;
wire  _GEN6009 = io_x[23] ? _GEN6008 : _GEN6005;
wire  _GEN6010 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6011 = io_x[10] ? _GEN6010 : _GEN3716;
wire  _GEN6012 = io_x[23] ? _GEN6011 : _GEN3741;
wire  _GEN6013 = io_x[16] ? _GEN6012 : _GEN6009;
wire  _GEN6014 = io_x[12] ? _GEN6013 : _GEN3893;
wire  _GEN6015 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6016 = io_x[14] ? _GEN6015 : _GEN3709;
wire  _GEN6017 = io_x[10] ? _GEN6016 : _GEN3711;
wire  _GEN6018 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6019 = io_x[10] ? _GEN6018 : _GEN3711;
wire  _GEN6020 = io_x[23] ? _GEN6019 : _GEN6017;
wire  _GEN6021 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6022 = io_x[14] ? _GEN6021 : _GEN3709;
wire  _GEN6023 = io_x[10] ? _GEN6022 : _GEN3716;
wire  _GEN6024 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6025 = io_x[14] ? _GEN6024 : _GEN3709;
wire  _GEN6026 = io_x[10] ? _GEN6025 : _GEN3716;
wire  _GEN6027 = io_x[23] ? _GEN6026 : _GEN6023;
wire  _GEN6028 = io_x[16] ? _GEN6027 : _GEN6020;
wire  _GEN6029 = io_x[12] ? _GEN6028 : _GEN4478;
wire  _GEN6030 = io_x[2] ? _GEN6029 : _GEN6014;
wire  _GEN6031 = io_x[9] ? _GEN6030 : _GEN6003;
wire  _GEN6032 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6033 = io_x[10] ? _GEN6032 : _GEN3711;
wire  _GEN6034 = io_x[23] ? _GEN6033 : _GEN3713;
wire  _GEN6035 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6036 = io_x[14] ? _GEN6035 : _GEN3709;
wire  _GEN6037 = io_x[10] ? _GEN6036 : _GEN3711;
wire  _GEN6038 = io_x[23] ? _GEN3713 : _GEN6037;
wire  _GEN6039 = io_x[16] ? _GEN6038 : _GEN6034;
wire  _GEN6040 = io_x[23] ? _GEN3741 : _GEN3713;
wire  _GEN6041 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6042 = io_x[14] ? _GEN6041 : _GEN3709;
wire  _GEN6043 = io_x[10] ? _GEN3716 : _GEN6042;
wire  _GEN6044 = io_x[23] ? _GEN6043 : _GEN3713;
wire  _GEN6045 = io_x[16] ? _GEN6044 : _GEN6040;
wire  _GEN6046 = io_x[12] ? _GEN6045 : _GEN6039;
wire  _GEN6047 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6048 = io_x[14] ? _GEN3709 : _GEN6047;
wire  _GEN6049 = io_x[10] ? _GEN6048 : _GEN3711;
wire  _GEN6050 = io_x[23] ? _GEN3741 : _GEN6049;
wire  _GEN6051 = io_x[16] ? _GEN6050 : _GEN3727;
wire  _GEN6052 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6053 = io_x[10] ? _GEN6052 : _GEN3711;
wire  _GEN6054 = io_x[23] ? _GEN3713 : _GEN6053;
wire  _GEN6055 = io_x[16] ? _GEN6054 : _GEN3707;
wire  _GEN6056 = io_x[12] ? _GEN6055 : _GEN6051;
wire  _GEN6057 = io_x[2] ? _GEN6056 : _GEN6046;
wire  _GEN6058 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6059 = io_x[10] ? _GEN6058 : _GEN3711;
wire  _GEN6060 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6061 = io_x[14] ? _GEN6060 : _GEN3709;
wire  _GEN6062 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6063 = io_x[10] ? _GEN6062 : _GEN6061;
wire  _GEN6064 = io_x[23] ? _GEN6063 : _GEN6059;
wire  _GEN6065 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6066 = io_x[14] ? _GEN6065 : _GEN3709;
wire  _GEN6067 = io_x[10] ? _GEN6066 : _GEN3711;
wire  _GEN6068 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6069 = io_x[14] ? _GEN6068 : _GEN3709;
wire  _GEN6070 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6071 = io_x[14] ? _GEN3708 : _GEN6070;
wire  _GEN6072 = io_x[10] ? _GEN6071 : _GEN6069;
wire  _GEN6073 = io_x[23] ? _GEN6072 : _GEN6067;
wire  _GEN6074 = io_x[16] ? _GEN6073 : _GEN6064;
wire  _GEN6075 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6076 = io_x[10] ? _GEN6075 : _GEN3711;
wire  _GEN6077 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6078 = io_x[14] ? _GEN6077 : _GEN3709;
wire  _GEN6079 = io_x[10] ? _GEN6078 : _GEN3711;
wire  _GEN6080 = io_x[23] ? _GEN6079 : _GEN6076;
wire  _GEN6081 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6082 = io_x[14] ? _GEN6081 : _GEN3709;
wire  _GEN6083 = io_x[10] ? _GEN6082 : _GEN3711;
wire  _GEN6084 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6085 = io_x[14] ? _GEN6084 : _GEN3709;
wire  _GEN6086 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6087 = io_x[14] ? _GEN6086 : _GEN3709;
wire  _GEN6088 = io_x[10] ? _GEN6087 : _GEN6085;
wire  _GEN6089 = io_x[23] ? _GEN6088 : _GEN6083;
wire  _GEN6090 = io_x[16] ? _GEN6089 : _GEN6080;
wire  _GEN6091 = io_x[12] ? _GEN6090 : _GEN6074;
wire  _GEN6092 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6093 = io_x[14] ? _GEN3709 : _GEN6092;
wire  _GEN6094 = io_x[10] ? _GEN6093 : _GEN3711;
wire  _GEN6095 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6096 = io_x[14] ? _GEN6095 : _GEN3708;
wire  _GEN6097 = io_x[10] ? _GEN3711 : _GEN6096;
wire  _GEN6098 = io_x[23] ? _GEN6097 : _GEN6094;
wire  _GEN6099 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6100 = io_x[10] ? _GEN6099 : _GEN3716;
wire  _GEN6101 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6102 = io_x[14] ? _GEN6101 : _GEN3709;
wire  _GEN6103 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6104 = io_x[14] ? _GEN3709 : _GEN6103;
wire  _GEN6105 = io_x[10] ? _GEN6104 : _GEN6102;
wire  _GEN6106 = io_x[23] ? _GEN6105 : _GEN6100;
wire  _GEN6107 = io_x[16] ? _GEN6106 : _GEN6098;
wire  _GEN6108 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN6109 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN6110 = io_x[23] ? _GEN6109 : _GEN6108;
wire  _GEN6111 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN6112 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6113 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6114 = io_x[14] ? _GEN6113 : _GEN3709;
wire  _GEN6115 = io_x[10] ? _GEN6114 : _GEN6112;
wire  _GEN6116 = io_x[23] ? _GEN6115 : _GEN6111;
wire  _GEN6117 = io_x[16] ? _GEN6116 : _GEN6110;
wire  _GEN6118 = io_x[12] ? _GEN6117 : _GEN6107;
wire  _GEN6119 = io_x[2] ? _GEN6118 : _GEN6091;
wire  _GEN6120 = io_x[9] ? _GEN6119 : _GEN6057;
wire  _GEN6121 = io_x[13] ? _GEN6120 : _GEN6031;
wire  _GEN6122 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6123 = io_x[14] ? _GEN6122 : _GEN3709;
wire  _GEN6124 = io_x[10] ? _GEN6123 : _GEN3711;
wire  _GEN6125 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6126 = io_x[14] ? _GEN6125 : _GEN3709;
wire  _GEN6127 = io_x[10] ? _GEN6126 : _GEN3716;
wire  _GEN6128 = io_x[23] ? _GEN6127 : _GEN6124;
wire  _GEN6129 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6130 = io_x[14] ? _GEN6129 : _GEN3709;
wire  _GEN6131 = io_x[10] ? _GEN6130 : _GEN3711;
wire  _GEN6132 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6133 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6134 = io_x[14] ? _GEN6133 : _GEN3709;
wire  _GEN6135 = io_x[10] ? _GEN6134 : _GEN6132;
wire  _GEN6136 = io_x[23] ? _GEN6135 : _GEN6131;
wire  _GEN6137 = io_x[16] ? _GEN6136 : _GEN6128;
wire  _GEN6138 = io_x[12] ? _GEN6137 : _GEN4478;
wire  _GEN6139 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6140 = io_x[14] ? _GEN6139 : _GEN3709;
wire  _GEN6141 = io_x[10] ? _GEN6140 : _GEN3716;
wire  _GEN6142 = io_x[23] ? _GEN3713 : _GEN6141;
wire  _GEN6143 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6144 = io_x[14] ? _GEN6143 : _GEN3708;
wire  _GEN6145 = io_x[10] ? _GEN6144 : _GEN3711;
wire  _GEN6146 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6147 = io_x[14] ? _GEN6146 : _GEN3709;
wire  _GEN6148 = io_x[10] ? _GEN6147 : _GEN3711;
wire  _GEN6149 = io_x[23] ? _GEN6148 : _GEN6145;
wire  _GEN6150 = io_x[16] ? _GEN6149 : _GEN6142;
wire  _GEN6151 = io_x[12] ? _GEN6150 : _GEN4478;
wire  _GEN6152 = io_x[2] ? _GEN6151 : _GEN6138;
wire  _GEN6153 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6154 = io_x[14] ? _GEN6153 : _GEN3709;
wire  _GEN6155 = io_x[10] ? _GEN3711 : _GEN6154;
wire  _GEN6156 = io_x[23] ? _GEN6155 : _GEN3713;
wire  _GEN6157 = io_x[16] ? _GEN6156 : _GEN3707;
wire  _GEN6158 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6159 = io_x[14] ? _GEN6158 : _GEN3709;
wire  _GEN6160 = io_x[10] ? _GEN3711 : _GEN6159;
wire  _GEN6161 = io_x[23] ? _GEN6160 : _GEN3741;
wire  _GEN6162 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6163 = io_x[14] ? _GEN6162 : _GEN3709;
wire  _GEN6164 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6165 = io_x[14] ? _GEN6164 : _GEN3709;
wire  _GEN6166 = io_x[10] ? _GEN6165 : _GEN6163;
wire  _GEN6167 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6168 = io_x[10] ? _GEN6167 : _GEN3716;
wire  _GEN6169 = io_x[23] ? _GEN6168 : _GEN6166;
wire  _GEN6170 = io_x[16] ? _GEN6169 : _GEN6161;
wire  _GEN6171 = io_x[12] ? _GEN6170 : _GEN6157;
wire  _GEN6172 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6173 = io_x[14] ? _GEN6172 : _GEN3709;
wire  _GEN6174 = io_x[10] ? _GEN6173 : _GEN3716;
wire  _GEN6175 = io_x[23] ? _GEN3713 : _GEN6174;
wire  _GEN6176 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6177 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6178 = io_x[14] ? _GEN6177 : _GEN3709;
wire  _GEN6179 = io_x[10] ? _GEN6178 : _GEN6176;
wire  _GEN6180 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6181 = io_x[14] ? _GEN6180 : _GEN3709;
wire  _GEN6182 = io_x[10] ? _GEN3711 : _GEN6181;
wire  _GEN6183 = io_x[23] ? _GEN6182 : _GEN6179;
wire  _GEN6184 = io_x[16] ? _GEN6183 : _GEN6175;
wire  _GEN6185 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6186 = io_x[14] ? _GEN6185 : _GEN3709;
wire  _GEN6187 = io_x[10] ? _GEN3711 : _GEN6186;
wire  _GEN6188 = io_x[23] ? _GEN3741 : _GEN6187;
wire  _GEN6189 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6190 = io_x[14] ? _GEN6189 : _GEN3709;
wire  _GEN6191 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6192 = io_x[10] ? _GEN6191 : _GEN6190;
wire  _GEN6193 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6194 = io_x[14] ? _GEN6193 : _GEN3709;
wire  _GEN6195 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6196 = io_x[14] ? _GEN6195 : _GEN3709;
wire  _GEN6197 = io_x[10] ? _GEN6196 : _GEN6194;
wire  _GEN6198 = io_x[23] ? _GEN6197 : _GEN6192;
wire  _GEN6199 = io_x[16] ? _GEN6198 : _GEN6188;
wire  _GEN6200 = io_x[12] ? _GEN6199 : _GEN6184;
wire  _GEN6201 = io_x[2] ? _GEN6200 : _GEN6171;
wire  _GEN6202 = io_x[9] ? _GEN6201 : _GEN6152;
wire  _GEN6203 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6204 = io_x[14] ? _GEN3709 : _GEN6203;
wire  _GEN6205 = io_x[10] ? _GEN6204 : _GEN3711;
wire  _GEN6206 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6207 = io_x[14] ? _GEN3709 : _GEN6206;
wire  _GEN6208 = io_x[10] ? _GEN6207 : _GEN3711;
wire  _GEN6209 = io_x[23] ? _GEN6208 : _GEN6205;
wire  _GEN6210 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6211 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6212 = io_x[14] ? _GEN6211 : _GEN6210;
wire  _GEN6213 = io_x[10] ? _GEN6212 : _GEN3711;
wire  _GEN6214 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6215 = io_x[14] ? _GEN3709 : _GEN6214;
wire  _GEN6216 = io_x[10] ? _GEN6215 : _GEN3711;
wire  _GEN6217 = io_x[23] ? _GEN6216 : _GEN6213;
wire  _GEN6218 = io_x[16] ? _GEN6217 : _GEN6209;
wire  _GEN6219 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN6220 = io_x[23] ? _GEN3741 : _GEN6219;
wire  _GEN6221 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6222 = io_x[14] ? _GEN6221 : _GEN3709;
wire  _GEN6223 = io_x[10] ? _GEN3716 : _GEN6222;
wire  _GEN6224 = io_x[23] ? _GEN3741 : _GEN6223;
wire  _GEN6225 = io_x[16] ? _GEN6224 : _GEN6220;
wire  _GEN6226 = io_x[12] ? _GEN6225 : _GEN6218;
wire  _GEN6227 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6228 = io_x[14] ? _GEN3709 : _GEN6227;
wire  _GEN6229 = io_x[10] ? _GEN6228 : _GEN3711;
wire  _GEN6230 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN6231 = io_x[23] ? _GEN6230 : _GEN6229;
wire  _GEN6232 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6233 = io_x[14] ? _GEN3709 : _GEN6232;
wire  _GEN6234 = io_x[10] ? _GEN6233 : _GEN3716;
wire  _GEN6235 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN6236 = io_x[23] ? _GEN6235 : _GEN6234;
wire  _GEN6237 = io_x[16] ? _GEN6236 : _GEN6231;
wire  _GEN6238 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN6239 = io_x[23] ? _GEN6238 : _GEN3713;
wire  _GEN6240 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6241 = io_x[10] ? _GEN3711 : _GEN6240;
wire  _GEN6242 = io_x[23] ? _GEN6241 : _GEN3713;
wire  _GEN6243 = io_x[16] ? _GEN6242 : _GEN6239;
wire  _GEN6244 = io_x[12] ? _GEN6243 : _GEN6237;
wire  _GEN6245 = io_x[2] ? _GEN6244 : _GEN6226;
wire  _GEN6246 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6247 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6248 = io_x[14] ? _GEN6247 : _GEN6246;
wire  _GEN6249 = io_x[10] ? _GEN3711 : _GEN6248;
wire  _GEN6250 = io_x[23] ? _GEN6249 : _GEN3713;
wire  _GEN6251 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6252 = io_x[14] ? _GEN6251 : _GEN3709;
wire  _GEN6253 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6254 = io_x[14] ? _GEN3708 : _GEN6253;
wire  _GEN6255 = io_x[10] ? _GEN6254 : _GEN6252;
wire  _GEN6256 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN6257 = io_x[23] ? _GEN6256 : _GEN6255;
wire  _GEN6258 = io_x[16] ? _GEN6257 : _GEN6250;
wire  _GEN6259 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6260 = io_x[14] ? _GEN6259 : _GEN3709;
wire  _GEN6261 = io_x[10] ? _GEN6260 : _GEN3711;
wire  _GEN6262 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6263 = io_x[14] ? _GEN6262 : _GEN3709;
wire  _GEN6264 = io_x[10] ? _GEN6263 : _GEN3711;
wire  _GEN6265 = io_x[23] ? _GEN6264 : _GEN6261;
wire  _GEN6266 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6267 = io_x[14] ? _GEN6266 : _GEN3709;
wire  _GEN6268 = io_x[10] ? _GEN3711 : _GEN6267;
wire  _GEN6269 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6270 = io_x[14] ? _GEN6269 : _GEN3709;
wire  _GEN6271 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6272 = io_x[14] ? _GEN6271 : _GEN3708;
wire  _GEN6273 = io_x[10] ? _GEN6272 : _GEN6270;
wire  _GEN6274 = io_x[23] ? _GEN6273 : _GEN6268;
wire  _GEN6275 = io_x[16] ? _GEN6274 : _GEN6265;
wire  _GEN6276 = io_x[12] ? _GEN6275 : _GEN6258;
wire  _GEN6277 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6278 = io_x[14] ? _GEN6277 : _GEN3709;
wire  _GEN6279 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6280 = io_x[14] ? _GEN3709 : _GEN6279;
wire  _GEN6281 = io_x[10] ? _GEN6280 : _GEN6278;
wire  _GEN6282 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6283 = io_x[10] ? _GEN3711 : _GEN6282;
wire  _GEN6284 = io_x[23] ? _GEN6283 : _GEN6281;
wire  _GEN6285 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6286 = io_x[14] ? _GEN6285 : _GEN3708;
wire  _GEN6287 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6288 = io_x[10] ? _GEN6287 : _GEN6286;
wire  _GEN6289 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6290 = io_x[14] ? _GEN6289 : _GEN3709;
wire  _GEN6291 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6292 = io_x[10] ? _GEN6291 : _GEN6290;
wire  _GEN6293 = io_x[23] ? _GEN6292 : _GEN6288;
wire  _GEN6294 = io_x[16] ? _GEN6293 : _GEN6284;
wire  _GEN6295 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6296 = io_x[14] ? _GEN3708 : _GEN6295;
wire  _GEN6297 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6298 = io_x[14] ? _GEN6297 : _GEN3709;
wire  _GEN6299 = io_x[10] ? _GEN6298 : _GEN6296;
wire  _GEN6300 = io_x[23] ? _GEN3741 : _GEN6299;
wire  _GEN6301 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6302 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6303 = io_x[14] ? _GEN6302 : _GEN6301;
wire  _GEN6304 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6305 = io_x[14] ? _GEN6304 : _GEN3708;
wire  _GEN6306 = io_x[10] ? _GEN6305 : _GEN6303;
wire  _GEN6307 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6308 = io_x[14] ? _GEN6307 : _GEN3709;
wire  _GEN6309 = io_x[10] ? _GEN6308 : _GEN3716;
wire  _GEN6310 = io_x[23] ? _GEN6309 : _GEN6306;
wire  _GEN6311 = io_x[16] ? _GEN6310 : _GEN6300;
wire  _GEN6312 = io_x[12] ? _GEN6311 : _GEN6294;
wire  _GEN6313 = io_x[2] ? _GEN6312 : _GEN6276;
wire  _GEN6314 = io_x[9] ? _GEN6313 : _GEN6245;
wire  _GEN6315 = io_x[13] ? _GEN6314 : _GEN6202;
wire  _GEN6316 = io_x[7] ? _GEN6315 : _GEN6121;
wire  _GEN6317 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6318 = io_x[14] ? _GEN6317 : _GEN3709;
wire  _GEN6319 = io_x[10] ? _GEN3711 : _GEN6318;
wire  _GEN6320 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6321 = io_x[14] ? _GEN6320 : _GEN3709;
wire  _GEN6322 = io_x[10] ? _GEN3711 : _GEN6321;
wire  _GEN6323 = io_x[23] ? _GEN6322 : _GEN6319;
wire  _GEN6324 = io_x[16] ? _GEN6323 : _GEN3707;
wire  _GEN6325 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6326 = io_x[14] ? _GEN3709 : _GEN6325;
wire  _GEN6327 = io_x[10] ? _GEN6326 : _GEN3711;
wire  _GEN6328 = io_x[23] ? _GEN3741 : _GEN6327;
wire  _GEN6329 = io_x[16] ? _GEN6328 : _GEN3727;
wire  _GEN6330 = io_x[12] ? _GEN6329 : _GEN6324;
wire  _GEN6331 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6332 = io_x[14] ? _GEN6331 : _GEN3709;
wire  _GEN6333 = io_x[10] ? _GEN3711 : _GEN6332;
wire  _GEN6334 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN6335 = io_x[23] ? _GEN6334 : _GEN6333;
wire  _GEN6336 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6337 = io_x[14] ? _GEN6336 : _GEN3709;
wire  _GEN6338 = io_x[10] ? _GEN3711 : _GEN6337;
wire  _GEN6339 = io_x[23] ? _GEN3713 : _GEN6338;
wire  _GEN6340 = io_x[16] ? _GEN6339 : _GEN6335;
wire  _GEN6341 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6342 = io_x[14] ? _GEN3709 : _GEN6341;
wire  _GEN6343 = io_x[10] ? _GEN6342 : _GEN3711;
wire  _GEN6344 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6345 = io_x[10] ? _GEN6344 : _GEN3711;
wire  _GEN6346 = io_x[23] ? _GEN6345 : _GEN6343;
wire  _GEN6347 = io_x[16] ? _GEN6346 : _GEN3707;
wire  _GEN6348 = io_x[12] ? _GEN6347 : _GEN6340;
wire  _GEN6349 = io_x[2] ? _GEN6348 : _GEN6330;
wire  _GEN6350 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6351 = io_x[10] ? _GEN3711 : _GEN6350;
wire  _GEN6352 = io_x[23] ? _GEN6351 : _GEN3713;
wire  _GEN6353 = io_x[16] ? _GEN6352 : _GEN3707;
wire  _GEN6354 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6355 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6356 = io_x[10] ? _GEN6355 : _GEN6354;
wire  _GEN6357 = io_x[23] ? _GEN6356 : _GEN3741;
wire  _GEN6358 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6359 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6360 = io_x[14] ? _GEN6359 : _GEN3709;
wire  _GEN6361 = io_x[10] ? _GEN6360 : _GEN6358;
wire  _GEN6362 = io_x[23] ? _GEN3741 : _GEN6361;
wire  _GEN6363 = io_x[16] ? _GEN6362 : _GEN6357;
wire  _GEN6364 = io_x[12] ? _GEN6363 : _GEN6353;
wire  _GEN6365 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6366 = io_x[14] ? _GEN6365 : _GEN3708;
wire  _GEN6367 = io_x[10] ? _GEN3711 : _GEN6366;
wire  _GEN6368 = io_x[23] ? _GEN6367 : _GEN3713;
wire  _GEN6369 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6370 = io_x[14] ? _GEN6369 : _GEN3708;
wire  _GEN6371 = io_x[10] ? _GEN3711 : _GEN6370;
wire  _GEN6372 = io_x[23] ? _GEN6371 : _GEN3741;
wire  _GEN6373 = io_x[16] ? _GEN6372 : _GEN6368;
wire  _GEN6374 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6375 = io_x[14] ? _GEN6374 : _GEN3708;
wire  _GEN6376 = io_x[10] ? _GEN6375 : _GEN3711;
wire  _GEN6377 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN6378 = io_x[23] ? _GEN6377 : _GEN6376;
wire  _GEN6379 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6380 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6381 = io_x[14] ? _GEN6380 : _GEN3709;
wire  _GEN6382 = io_x[10] ? _GEN6381 : _GEN6379;
wire  _GEN6383 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6384 = io_x[10] ? _GEN3711 : _GEN6383;
wire  _GEN6385 = io_x[23] ? _GEN6384 : _GEN6382;
wire  _GEN6386 = io_x[16] ? _GEN6385 : _GEN6378;
wire  _GEN6387 = io_x[12] ? _GEN6386 : _GEN6373;
wire  _GEN6388 = io_x[2] ? _GEN6387 : _GEN6364;
wire  _GEN6389 = io_x[9] ? _GEN6388 : _GEN6349;
wire  _GEN6390 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6391 = io_x[14] ? _GEN3709 : _GEN6390;
wire  _GEN6392 = io_x[10] ? _GEN6391 : _GEN3711;
wire  _GEN6393 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6394 = io_x[10] ? _GEN6393 : _GEN3716;
wire  _GEN6395 = io_x[23] ? _GEN6394 : _GEN6392;
wire  _GEN6396 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6397 = io_x[10] ? _GEN6396 : _GEN3711;
wire  _GEN6398 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6399 = io_x[10] ? _GEN6398 : _GEN3711;
wire  _GEN6400 = io_x[23] ? _GEN6399 : _GEN6397;
wire  _GEN6401 = io_x[16] ? _GEN6400 : _GEN6395;
wire  _GEN6402 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6403 = io_x[10] ? _GEN3711 : _GEN6402;
wire  _GEN6404 = io_x[23] ? _GEN6403 : _GEN3741;
wire  _GEN6405 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6406 = io_x[14] ? _GEN3709 : _GEN6405;
wire  _GEN6407 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6408 = io_x[10] ? _GEN6407 : _GEN6406;
wire  _GEN6409 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6410 = io_x[14] ? _GEN3708 : _GEN6409;
wire  _GEN6411 = io_x[10] ? _GEN3711 : _GEN6410;
wire  _GEN6412 = io_x[23] ? _GEN6411 : _GEN6408;
wire  _GEN6413 = io_x[16] ? _GEN6412 : _GEN6404;
wire  _GEN6414 = io_x[12] ? _GEN6413 : _GEN6401;
wire  _GEN6415 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6416 = io_x[10] ? _GEN6415 : _GEN3711;
wire  _GEN6417 = io_x[23] ? _GEN3713 : _GEN6416;
wire  _GEN6418 = io_x[16] ? _GEN6417 : _GEN3727;
wire  _GEN6419 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6420 = io_x[14] ? _GEN3708 : _GEN6419;
wire  _GEN6421 = io_x[10] ? _GEN3711 : _GEN6420;
wire  _GEN6422 = io_x[23] ? _GEN3741 : _GEN6421;
wire  _GEN6423 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6424 = io_x[14] ? _GEN3708 : _GEN6423;
wire  _GEN6425 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6426 = io_x[10] ? _GEN6425 : _GEN6424;
wire  _GEN6427 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6428 = io_x[14] ? _GEN6427 : _GEN3709;
wire  _GEN6429 = io_x[10] ? _GEN3716 : _GEN6428;
wire  _GEN6430 = io_x[23] ? _GEN6429 : _GEN6426;
wire  _GEN6431 = io_x[16] ? _GEN6430 : _GEN6422;
wire  _GEN6432 = io_x[12] ? _GEN6431 : _GEN6418;
wire  _GEN6433 = io_x[2] ? _GEN6432 : _GEN6414;
wire  _GEN6434 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6435 = io_x[14] ? _GEN6434 : _GEN3709;
wire  _GEN6436 = io_x[10] ? _GEN6435 : _GEN3711;
wire  _GEN6437 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6438 = io_x[14] ? _GEN3709 : _GEN6437;
wire  _GEN6439 = io_x[10] ? _GEN6438 : _GEN3716;
wire  _GEN6440 = io_x[23] ? _GEN6439 : _GEN6436;
wire  _GEN6441 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6442 = io_x[14] ? _GEN6441 : _GEN3709;
wire  _GEN6443 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6444 = io_x[14] ? _GEN6443 : _GEN3709;
wire  _GEN6445 = io_x[10] ? _GEN6444 : _GEN6442;
wire  _GEN6446 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6447 = io_x[10] ? _GEN6446 : _GEN3716;
wire  _GEN6448 = io_x[23] ? _GEN6447 : _GEN6445;
wire  _GEN6449 = io_x[16] ? _GEN6448 : _GEN6440;
wire  _GEN6450 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6451 = io_x[14] ? _GEN3709 : _GEN6450;
wire  _GEN6452 = io_x[10] ? _GEN6451 : _GEN3711;
wire  _GEN6453 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6454 = io_x[10] ? _GEN6453 : _GEN3711;
wire  _GEN6455 = io_x[23] ? _GEN6454 : _GEN6452;
wire  _GEN6456 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6457 = io_x[14] ? _GEN6456 : _GEN3708;
wire  _GEN6458 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6459 = io_x[14] ? _GEN6458 : _GEN3709;
wire  _GEN6460 = io_x[10] ? _GEN6459 : _GEN6457;
wire  _GEN6461 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6462 = io_x[10] ? _GEN6461 : _GEN3711;
wire  _GEN6463 = io_x[23] ? _GEN6462 : _GEN6460;
wire  _GEN6464 = io_x[16] ? _GEN6463 : _GEN6455;
wire  _GEN6465 = io_x[12] ? _GEN6464 : _GEN6449;
wire  _GEN6466 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6467 = io_x[14] ? _GEN6466 : _GEN3708;
wire  _GEN6468 = io_x[10] ? _GEN6467 : _GEN3711;
wire  _GEN6469 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6470 = io_x[14] ? _GEN3709 : _GEN6469;
wire  _GEN6471 = io_x[10] ? _GEN3711 : _GEN6470;
wire  _GEN6472 = io_x[23] ? _GEN6471 : _GEN6468;
wire  _GEN6473 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6474 = io_x[10] ? _GEN6473 : _GEN3716;
wire  _GEN6475 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6476 = io_x[14] ? _GEN6475 : _GEN3709;
wire  _GEN6477 = io_x[10] ? _GEN3716 : _GEN6476;
wire  _GEN6478 = io_x[23] ? _GEN6477 : _GEN6474;
wire  _GEN6479 = io_x[16] ? _GEN6478 : _GEN6472;
wire  _GEN6480 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6481 = io_x[14] ? _GEN3708 : _GEN6480;
wire  _GEN6482 = io_x[10] ? _GEN6481 : _GEN3716;
wire  _GEN6483 = io_x[23] ? _GEN3713 : _GEN6482;
wire  _GEN6484 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6485 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6486 = io_x[14] ? _GEN6485 : _GEN3709;
wire  _GEN6487 = io_x[10] ? _GEN6486 : _GEN6484;
wire  _GEN6488 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6489 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6490 = io_x[14] ? _GEN6489 : _GEN6488;
wire  _GEN6491 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6492 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6493 = io_x[14] ? _GEN6492 : _GEN6491;
wire  _GEN6494 = io_x[10] ? _GEN6493 : _GEN6490;
wire  _GEN6495 = io_x[23] ? _GEN6494 : _GEN6487;
wire  _GEN6496 = io_x[16] ? _GEN6495 : _GEN6483;
wire  _GEN6497 = io_x[12] ? _GEN6496 : _GEN6479;
wire  _GEN6498 = io_x[2] ? _GEN6497 : _GEN6465;
wire  _GEN6499 = io_x[9] ? _GEN6498 : _GEN6433;
wire  _GEN6500 = io_x[13] ? _GEN6499 : _GEN6389;
wire  _GEN6501 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6502 = io_x[14] ? _GEN6501 : _GEN3709;
wire  _GEN6503 = io_x[10] ? _GEN6502 : _GEN3716;
wire  _GEN6504 = io_x[23] ? _GEN6503 : _GEN3741;
wire  _GEN6505 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6506 = io_x[14] ? _GEN6505 : _GEN3709;
wire  _GEN6507 = io_x[10] ? _GEN6506 : _GEN3711;
wire  _GEN6508 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6509 = io_x[14] ? _GEN6508 : _GEN3709;
wire  _GEN6510 = io_x[10] ? _GEN6509 : _GEN3716;
wire  _GEN6511 = io_x[23] ? _GEN6510 : _GEN6507;
wire  _GEN6512 = io_x[16] ? _GEN6511 : _GEN6504;
wire  _GEN6513 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6514 = io_x[14] ? _GEN6513 : _GEN3708;
wire  _GEN6515 = io_x[10] ? _GEN6514 : _GEN3716;
wire  _GEN6516 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6517 = io_x[14] ? _GEN6516 : _GEN3709;
wire  _GEN6518 = io_x[10] ? _GEN6517 : _GEN3711;
wire  _GEN6519 = io_x[23] ? _GEN6518 : _GEN6515;
wire  _GEN6520 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6521 = io_x[14] ? _GEN6520 : _GEN3709;
wire  _GEN6522 = io_x[10] ? _GEN6521 : _GEN3711;
wire  _GEN6523 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6524 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6525 = io_x[14] ? _GEN6524 : _GEN6523;
wire  _GEN6526 = io_x[10] ? _GEN6525 : _GEN3711;
wire  _GEN6527 = io_x[23] ? _GEN6526 : _GEN6522;
wire  _GEN6528 = io_x[16] ? _GEN6527 : _GEN6519;
wire  _GEN6529 = io_x[12] ? _GEN6528 : _GEN6512;
wire  _GEN6530 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6531 = io_x[14] ? _GEN6530 : _GEN3709;
wire  _GEN6532 = io_x[10] ? _GEN6531 : _GEN3711;
wire  _GEN6533 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6534 = io_x[10] ? _GEN6533 : _GEN3711;
wire  _GEN6535 = io_x[23] ? _GEN6534 : _GEN6532;
wire  _GEN6536 = io_x[16] ? _GEN3727 : _GEN6535;
wire  _GEN6537 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6538 = io_x[14] ? _GEN6537 : _GEN3709;
wire  _GEN6539 = io_x[10] ? _GEN6538 : _GEN3711;
wire  _GEN6540 = io_x[10] ? _GEN3711 : _GEN3716;
wire  _GEN6541 = io_x[23] ? _GEN6540 : _GEN6539;
wire  _GEN6542 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6543 = io_x[14] ? _GEN3709 : _GEN6542;
wire  _GEN6544 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6545 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6546 = io_x[14] ? _GEN6545 : _GEN6544;
wire  _GEN6547 = io_x[10] ? _GEN6546 : _GEN6543;
wire  _GEN6548 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6549 = io_x[14] ? _GEN6548 : _GEN3708;
wire  _GEN6550 = io_x[10] ? _GEN6549 : _GEN3716;
wire  _GEN6551 = io_x[23] ? _GEN6550 : _GEN6547;
wire  _GEN6552 = io_x[16] ? _GEN6551 : _GEN6541;
wire  _GEN6553 = io_x[12] ? _GEN6552 : _GEN6536;
wire  _GEN6554 = io_x[2] ? _GEN6553 : _GEN6529;
wire  _GEN6555 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6556 = io_x[14] ? _GEN6555 : _GEN3709;
wire  _GEN6557 = io_x[10] ? _GEN3711 : _GEN6556;
wire  _GEN6558 = io_x[23] ? _GEN3713 : _GEN6557;
wire  _GEN6559 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6560 = io_x[14] ? _GEN6559 : _GEN3708;
wire  _GEN6561 = io_x[10] ? _GEN3711 : _GEN6560;
wire  _GEN6562 = io_x[23] ? _GEN3713 : _GEN6561;
wire  _GEN6563 = io_x[16] ? _GEN6562 : _GEN6558;
wire  _GEN6564 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN6565 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6566 = io_x[10] ? _GEN6565 : _GEN3716;
wire  _GEN6567 = io_x[23] ? _GEN6566 : _GEN6564;
wire  _GEN6568 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6569 = io_x[14] ? _GEN3708 : _GEN6568;
wire  _GEN6570 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6571 = io_x[14] ? _GEN3708 : _GEN6570;
wire  _GEN6572 = io_x[10] ? _GEN6571 : _GEN6569;
wire  _GEN6573 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6574 = io_x[14] ? _GEN6573 : _GEN3709;
wire  _GEN6575 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6576 = io_x[14] ? _GEN6575 : _GEN3708;
wire  _GEN6577 = io_x[10] ? _GEN6576 : _GEN6574;
wire  _GEN6578 = io_x[23] ? _GEN6577 : _GEN6572;
wire  _GEN6579 = io_x[16] ? _GEN6578 : _GEN6567;
wire  _GEN6580 = io_x[12] ? _GEN6579 : _GEN6563;
wire  _GEN6581 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6582 = io_x[14] ? _GEN6581 : _GEN3709;
wire  _GEN6583 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6584 = io_x[14] ? _GEN6583 : _GEN3708;
wire  _GEN6585 = io_x[10] ? _GEN6584 : _GEN6582;
wire  _GEN6586 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6587 = io_x[14] ? _GEN6586 : _GEN3709;
wire  _GEN6588 = io_x[10] ? _GEN3716 : _GEN6587;
wire  _GEN6589 = io_x[23] ? _GEN6588 : _GEN6585;
wire  _GEN6590 = io_x[16] ? _GEN6589 : _GEN3727;
wire  _GEN6591 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6592 = io_x[14] ? _GEN6591 : _GEN3708;
wire  _GEN6593 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6594 = io_x[14] ? _GEN3709 : _GEN6593;
wire  _GEN6595 = io_x[10] ? _GEN6594 : _GEN6592;
wire  _GEN6596 = io_x[23] ? _GEN3741 : _GEN6595;
wire  _GEN6597 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6598 = io_x[14] ? _GEN3708 : _GEN6597;
wire  _GEN6599 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6600 = io_x[14] ? _GEN3709 : _GEN6599;
wire  _GEN6601 = io_x[10] ? _GEN6600 : _GEN6598;
wire  _GEN6602 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6603 = io_x[14] ? _GEN3708 : _GEN6602;
wire  _GEN6604 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6605 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6606 = io_x[14] ? _GEN6605 : _GEN6604;
wire  _GEN6607 = io_x[10] ? _GEN6606 : _GEN6603;
wire  _GEN6608 = io_x[23] ? _GEN6607 : _GEN6601;
wire  _GEN6609 = io_x[16] ? _GEN6608 : _GEN6596;
wire  _GEN6610 = io_x[12] ? _GEN6609 : _GEN6590;
wire  _GEN6611 = io_x[2] ? _GEN6610 : _GEN6580;
wire  _GEN6612 = io_x[9] ? _GEN6611 : _GEN6554;
wire  _GEN6613 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6614 = io_x[14] ? _GEN6613 : _GEN3708;
wire  _GEN6615 = io_x[10] ? _GEN6614 : _GEN3716;
wire  _GEN6616 = io_x[23] ? _GEN6615 : _GEN3741;
wire  _GEN6617 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6618 = io_x[14] ? _GEN6617 : _GEN3708;
wire  _GEN6619 = io_x[10] ? _GEN6618 : _GEN3711;
wire  _GEN6620 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6621 = io_x[14] ? _GEN6620 : _GEN3709;
wire  _GEN6622 = io_x[10] ? _GEN6621 : _GEN3711;
wire  _GEN6623 = io_x[23] ? _GEN6622 : _GEN6619;
wire  _GEN6624 = io_x[16] ? _GEN6623 : _GEN6616;
wire  _GEN6625 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6626 = io_x[14] ? _GEN3709 : _GEN6625;
wire  _GEN6627 = io_x[10] ? _GEN6626 : _GEN3711;
wire  _GEN6628 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6629 = io_x[14] ? _GEN3709 : _GEN6628;
wire  _GEN6630 = io_x[10] ? _GEN6629 : _GEN3711;
wire  _GEN6631 = io_x[23] ? _GEN6630 : _GEN6627;
wire  _GEN6632 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6633 = io_x[14] ? _GEN3708 : _GEN6632;
wire  _GEN6634 = io_x[10] ? _GEN6633 : _GEN3711;
wire  _GEN6635 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6636 = io_x[14] ? _GEN3709 : _GEN6635;
wire  _GEN6637 = io_x[10] ? _GEN6636 : _GEN3711;
wire  _GEN6638 = io_x[23] ? _GEN6637 : _GEN6634;
wire  _GEN6639 = io_x[16] ? _GEN6638 : _GEN6631;
wire  _GEN6640 = io_x[12] ? _GEN6639 : _GEN6624;
wire  _GEN6641 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6642 = io_x[14] ? _GEN6641 : _GEN3709;
wire  _GEN6643 = io_x[10] ? _GEN6642 : _GEN3711;
wire  _GEN6644 = io_x[23] ? _GEN3713 : _GEN6643;
wire  _GEN6645 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6646 = io_x[14] ? _GEN3709 : _GEN6645;
wire  _GEN6647 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6648 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6649 = io_x[14] ? _GEN6648 : _GEN6647;
wire  _GEN6650 = io_x[10] ? _GEN6649 : _GEN6646;
wire  _GEN6651 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6652 = io_x[14] ? _GEN6651 : _GEN3709;
wire  _GEN6653 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6654 = io_x[14] ? _GEN6653 : _GEN3709;
wire  _GEN6655 = io_x[10] ? _GEN6654 : _GEN6652;
wire  _GEN6656 = io_x[23] ? _GEN6655 : _GEN6650;
wire  _GEN6657 = io_x[16] ? _GEN6656 : _GEN6644;
wire  _GEN6658 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6659 = io_x[14] ? _GEN6658 : _GEN3709;
wire  _GEN6660 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6661 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6662 = io_x[14] ? _GEN6661 : _GEN6660;
wire  _GEN6663 = io_x[10] ? _GEN6662 : _GEN6659;
wire  _GEN6664 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6665 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6666 = io_x[14] ? _GEN6665 : _GEN6664;
wire  _GEN6667 = io_x[10] ? _GEN6666 : _GEN3716;
wire  _GEN6668 = io_x[23] ? _GEN6667 : _GEN6663;
wire  _GEN6669 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6670 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6671 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6672 = io_x[14] ? _GEN6671 : _GEN6670;
wire  _GEN6673 = io_x[10] ? _GEN6672 : _GEN6669;
wire  _GEN6674 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6675 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6676 = io_x[14] ? _GEN6675 : _GEN6674;
wire  _GEN6677 = io_x[10] ? _GEN6676 : _GEN3711;
wire  _GEN6678 = io_x[23] ? _GEN6677 : _GEN6673;
wire  _GEN6679 = io_x[16] ? _GEN6678 : _GEN6668;
wire  _GEN6680 = io_x[12] ? _GEN6679 : _GEN6657;
wire  _GEN6681 = io_x[2] ? _GEN6680 : _GEN6640;
wire  _GEN6682 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6683 = io_x[10] ? _GEN3716 : _GEN6682;
wire  _GEN6684 = io_x[23] ? _GEN6683 : _GEN3741;
wire  _GEN6685 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6686 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6687 = io_x[14] ? _GEN6686 : _GEN6685;
wire  _GEN6688 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6689 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6690 = io_x[14] ? _GEN6689 : _GEN6688;
wire  _GEN6691 = io_x[10] ? _GEN6690 : _GEN6687;
wire  _GEN6692 = io_x[10] ? _GEN3716 : _GEN3711;
wire  _GEN6693 = io_x[23] ? _GEN6692 : _GEN6691;
wire  _GEN6694 = io_x[16] ? _GEN6693 : _GEN6684;
wire  _GEN6695 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6696 = io_x[14] ? _GEN3708 : _GEN6695;
wire  _GEN6697 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6698 = io_x[14] ? _GEN6697 : _GEN3709;
wire  _GEN6699 = io_x[10] ? _GEN6698 : _GEN6696;
wire  _GEN6700 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6701 = io_x[14] ? _GEN3709 : _GEN6700;
wire  _GEN6702 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6703 = io_x[14] ? _GEN6702 : _GEN3708;
wire  _GEN6704 = io_x[10] ? _GEN6703 : _GEN6701;
wire  _GEN6705 = io_x[23] ? _GEN6704 : _GEN6699;
wire  _GEN6706 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6707 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6708 = io_x[14] ? _GEN6707 : _GEN6706;
wire  _GEN6709 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6710 = io_x[14] ? _GEN6709 : _GEN3709;
wire  _GEN6711 = io_x[10] ? _GEN6710 : _GEN6708;
wire  _GEN6712 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6713 = io_x[14] ? _GEN3708 : _GEN6712;
wire  _GEN6714 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6715 = io_x[14] ? _GEN6714 : _GEN3708;
wire  _GEN6716 = io_x[10] ? _GEN6715 : _GEN6713;
wire  _GEN6717 = io_x[23] ? _GEN6716 : _GEN6711;
wire  _GEN6718 = io_x[16] ? _GEN6717 : _GEN6705;
wire  _GEN6719 = io_x[12] ? _GEN6718 : _GEN6694;
wire  _GEN6720 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6721 = io_x[14] ? _GEN6720 : _GEN3708;
wire  _GEN6722 = io_x[14] ? _GEN3709 : _GEN3708;
wire  _GEN6723 = io_x[10] ? _GEN6722 : _GEN6721;
wire  _GEN6724 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6725 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6726 = io_x[14] ? _GEN6725 : _GEN6724;
wire  _GEN6727 = io_x[14] ? _GEN3708 : _GEN3709;
wire  _GEN6728 = io_x[10] ? _GEN6727 : _GEN6726;
wire  _GEN6729 = io_x[23] ? _GEN6728 : _GEN6723;
wire  _GEN6730 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6731 = io_x[14] ? _GEN3708 : _GEN6730;
wire  _GEN6732 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6733 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6734 = io_x[14] ? _GEN6733 : _GEN6732;
wire  _GEN6735 = io_x[10] ? _GEN6734 : _GEN6731;
wire  _GEN6736 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6737 = io_x[14] ? _GEN3708 : _GEN6736;
wire  _GEN6738 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6739 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6740 = io_x[14] ? _GEN6739 : _GEN6738;
wire  _GEN6741 = io_x[10] ? _GEN6740 : _GEN6737;
wire  _GEN6742 = io_x[23] ? _GEN6741 : _GEN6735;
wire  _GEN6743 = io_x[16] ? _GEN6742 : _GEN6729;
wire  _GEN6744 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6745 = io_x[14] ? _GEN6744 : _GEN3708;
wire  _GEN6746 = io_x[10] ? _GEN6745 : _GEN3711;
wire  _GEN6747 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6748 = io_x[14] ? _GEN6747 : _GEN3708;
wire  _GEN6749 = io_x[10] ? _GEN6748 : _GEN3716;
wire  _GEN6750 = io_x[23] ? _GEN6749 : _GEN6746;
wire  _GEN6751 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6752 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6753 = io_x[14] ? _GEN6752 : _GEN6751;
wire  _GEN6754 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6755 = io_x[14] ? _GEN6754 : _GEN3708;
wire  _GEN6756 = io_x[10] ? _GEN6755 : _GEN6753;
wire  _GEN6757 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6758 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6759 = io_x[14] ? _GEN6758 : _GEN6757;
wire  _GEN6760 = io_x[6] ? _GEN3719 : _GEN3720;
wire  _GEN6761 = io_x[6] ? _GEN3720 : _GEN3719;
wire  _GEN6762 = io_x[14] ? _GEN6761 : _GEN6760;
wire  _GEN6763 = io_x[10] ? _GEN6762 : _GEN6759;
wire  _GEN6764 = io_x[23] ? _GEN6763 : _GEN6756;
wire  _GEN6765 = io_x[16] ? _GEN6764 : _GEN6750;
wire  _GEN6766 = io_x[12] ? _GEN6765 : _GEN6743;
wire  _GEN6767 = io_x[2] ? _GEN6766 : _GEN6719;
wire  _GEN6768 = io_x[9] ? _GEN6767 : _GEN6681;
wire  _GEN6769 = io_x[13] ? _GEN6768 : _GEN6612;
wire  _GEN6770 = io_x[7] ? _GEN6769 : _GEN6500;
wire  _GEN6771 = io_x[15] ? _GEN6770 : _GEN6316;
wire  _GEN6772 = io_x[3] ? _GEN6771 : _GEN5965;
wire  _GEN6773 = io_x[26] ? _GEN6772 : _GEN5365;
assign io_y[8] = _GEN6773;
wire  _GEN6774 = 1'b0;
wire  _GEN6775 = 1'b1;
wire  _GEN6776 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6777 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6778 = io_x[9] ? _GEN6777 : _GEN6776;
wire  _GEN6779 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6780 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6781 = io_x[9] ? _GEN6780 : _GEN6779;
wire  _GEN6782 = io_x[23] ? _GEN6781 : _GEN6778;
wire  _GEN6783 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6784 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6785 = io_x[9] ? _GEN6784 : _GEN6783;
wire  _GEN6786 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6787 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6788 = io_x[9] ? _GEN6787 : _GEN6786;
wire  _GEN6789 = io_x[23] ? _GEN6788 : _GEN6785;
wire  _GEN6790 = io_x[25] ? _GEN6789 : _GEN6782;
wire  _GEN6791 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6792 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6793 = io_x[9] ? _GEN6792 : _GEN6791;
wire  _GEN6794 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6795 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6796 = io_x[9] ? _GEN6795 : _GEN6794;
wire  _GEN6797 = io_x[23] ? _GEN6796 : _GEN6793;
wire  _GEN6798 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6799 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6800 = io_x[9] ? _GEN6799 : _GEN6798;
wire  _GEN6801 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6802 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6803 = io_x[9] ? _GEN6802 : _GEN6801;
wire  _GEN6804 = io_x[23] ? _GEN6803 : _GEN6800;
wire  _GEN6805 = io_x[25] ? _GEN6804 : _GEN6797;
wire  _GEN6806 = io_x[5] ? _GEN6805 : _GEN6790;
wire  _GEN6807 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6808 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6809 = io_x[9] ? _GEN6808 : _GEN6807;
wire  _GEN6810 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6811 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6812 = io_x[9] ? _GEN6811 : _GEN6810;
wire  _GEN6813 = io_x[23] ? _GEN6812 : _GEN6809;
wire  _GEN6814 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6815 = 1'b1;
wire  _GEN6816 = io_x[9] ? _GEN6815 : _GEN6814;
wire  _GEN6817 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6818 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6819 = io_x[9] ? _GEN6818 : _GEN6817;
wire  _GEN6820 = io_x[23] ? _GEN6819 : _GEN6816;
wire  _GEN6821 = io_x[25] ? _GEN6820 : _GEN6813;
wire  _GEN6822 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6823 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6824 = io_x[9] ? _GEN6823 : _GEN6822;
wire  _GEN6825 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6826 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6827 = io_x[9] ? _GEN6826 : _GEN6825;
wire  _GEN6828 = io_x[23] ? _GEN6827 : _GEN6824;
wire  _GEN6829 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6830 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6831 = io_x[9] ? _GEN6830 : _GEN6829;
wire  _GEN6832 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6833 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6834 = io_x[9] ? _GEN6833 : _GEN6832;
wire  _GEN6835 = io_x[23] ? _GEN6834 : _GEN6831;
wire  _GEN6836 = io_x[25] ? _GEN6835 : _GEN6828;
wire  _GEN6837 = io_x[5] ? _GEN6836 : _GEN6821;
wire  _GEN6838 = io_x[21] ? _GEN6837 : _GEN6806;
wire  _GEN6839 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6840 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6841 = io_x[9] ? _GEN6840 : _GEN6839;
wire  _GEN6842 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6843 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6844 = io_x[9] ? _GEN6843 : _GEN6842;
wire  _GEN6845 = io_x[23] ? _GEN6844 : _GEN6841;
wire  _GEN6846 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6847 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6848 = io_x[9] ? _GEN6847 : _GEN6846;
wire  _GEN6849 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6850 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6851 = io_x[9] ? _GEN6850 : _GEN6849;
wire  _GEN6852 = io_x[23] ? _GEN6851 : _GEN6848;
wire  _GEN6853 = io_x[25] ? _GEN6852 : _GEN6845;
wire  _GEN6854 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6855 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6856 = io_x[9] ? _GEN6855 : _GEN6854;
wire  _GEN6857 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6858 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6859 = io_x[9] ? _GEN6858 : _GEN6857;
wire  _GEN6860 = io_x[23] ? _GEN6859 : _GEN6856;
wire  _GEN6861 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6862 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6863 = io_x[9] ? _GEN6862 : _GEN6861;
wire  _GEN6864 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6865 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6866 = io_x[9] ? _GEN6865 : _GEN6864;
wire  _GEN6867 = io_x[23] ? _GEN6866 : _GEN6863;
wire  _GEN6868 = io_x[25] ? _GEN6867 : _GEN6860;
wire  _GEN6869 = io_x[5] ? _GEN6868 : _GEN6853;
wire  _GEN6870 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6871 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6872 = io_x[9] ? _GEN6871 : _GEN6870;
wire  _GEN6873 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6874 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6875 = io_x[9] ? _GEN6874 : _GEN6873;
wire  _GEN6876 = io_x[23] ? _GEN6875 : _GEN6872;
wire  _GEN6877 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6878 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6879 = io_x[9] ? _GEN6878 : _GEN6877;
wire  _GEN6880 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6881 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6882 = io_x[9] ? _GEN6881 : _GEN6880;
wire  _GEN6883 = io_x[23] ? _GEN6882 : _GEN6879;
wire  _GEN6884 = io_x[25] ? _GEN6883 : _GEN6876;
wire  _GEN6885 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6886 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6887 = io_x[9] ? _GEN6886 : _GEN6885;
wire  _GEN6888 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6889 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6890 = io_x[9] ? _GEN6889 : _GEN6888;
wire  _GEN6891 = io_x[23] ? _GEN6890 : _GEN6887;
wire  _GEN6892 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6893 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6894 = io_x[9] ? _GEN6893 : _GEN6892;
wire  _GEN6895 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6896 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6897 = io_x[9] ? _GEN6896 : _GEN6895;
wire  _GEN6898 = io_x[23] ? _GEN6897 : _GEN6894;
wire  _GEN6899 = io_x[25] ? _GEN6898 : _GEN6891;
wire  _GEN6900 = io_x[5] ? _GEN6899 : _GEN6884;
wire  _GEN6901 = io_x[21] ? _GEN6900 : _GEN6869;
wire  _GEN6902 = io_x[13] ? _GEN6901 : _GEN6838;
wire  _GEN6903 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6904 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6905 = io_x[9] ? _GEN6904 : _GEN6903;
wire  _GEN6906 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6907 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6908 = io_x[9] ? _GEN6907 : _GEN6906;
wire  _GEN6909 = io_x[23] ? _GEN6908 : _GEN6905;
wire  _GEN6910 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6911 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6912 = io_x[9] ? _GEN6911 : _GEN6910;
wire  _GEN6913 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6914 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6915 = io_x[9] ? _GEN6914 : _GEN6913;
wire  _GEN6916 = io_x[23] ? _GEN6915 : _GEN6912;
wire  _GEN6917 = io_x[25] ? _GEN6916 : _GEN6909;
wire  _GEN6918 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6919 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6920 = io_x[9] ? _GEN6919 : _GEN6918;
wire  _GEN6921 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6922 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6923 = io_x[9] ? _GEN6922 : _GEN6921;
wire  _GEN6924 = io_x[23] ? _GEN6923 : _GEN6920;
wire  _GEN6925 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6926 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6927 = io_x[9] ? _GEN6926 : _GEN6925;
wire  _GEN6928 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6929 = io_x[9] ? _GEN6928 : _GEN6815;
wire  _GEN6930 = io_x[23] ? _GEN6929 : _GEN6927;
wire  _GEN6931 = io_x[25] ? _GEN6930 : _GEN6924;
wire  _GEN6932 = io_x[5] ? _GEN6931 : _GEN6917;
wire  _GEN6933 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6934 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6935 = io_x[9] ? _GEN6934 : _GEN6933;
wire  _GEN6936 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6937 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6938 = io_x[9] ? _GEN6937 : _GEN6936;
wire  _GEN6939 = io_x[23] ? _GEN6938 : _GEN6935;
wire  _GEN6940 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6941 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6942 = io_x[9] ? _GEN6941 : _GEN6940;
wire  _GEN6943 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6944 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6945 = io_x[9] ? _GEN6944 : _GEN6943;
wire  _GEN6946 = io_x[23] ? _GEN6945 : _GEN6942;
wire  _GEN6947 = io_x[25] ? _GEN6946 : _GEN6939;
wire  _GEN6948 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6949 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6950 = io_x[9] ? _GEN6949 : _GEN6948;
wire  _GEN6951 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6952 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6953 = io_x[9] ? _GEN6952 : _GEN6951;
wire  _GEN6954 = io_x[23] ? _GEN6953 : _GEN6950;
wire  _GEN6955 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6956 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6957 = io_x[9] ? _GEN6956 : _GEN6955;
wire  _GEN6958 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6959 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6960 = io_x[9] ? _GEN6959 : _GEN6958;
wire  _GEN6961 = io_x[23] ? _GEN6960 : _GEN6957;
wire  _GEN6962 = io_x[25] ? _GEN6961 : _GEN6954;
wire  _GEN6963 = io_x[5] ? _GEN6962 : _GEN6947;
wire  _GEN6964 = io_x[21] ? _GEN6963 : _GEN6932;
wire  _GEN6965 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6966 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6967 = io_x[9] ? _GEN6966 : _GEN6965;
wire  _GEN6968 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6969 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6970 = io_x[9] ? _GEN6969 : _GEN6968;
wire  _GEN6971 = io_x[23] ? _GEN6970 : _GEN6967;
wire  _GEN6972 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6973 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6974 = io_x[9] ? _GEN6973 : _GEN6972;
wire  _GEN6975 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6976 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6977 = io_x[9] ? _GEN6976 : _GEN6975;
wire  _GEN6978 = io_x[23] ? _GEN6977 : _GEN6974;
wire  _GEN6979 = io_x[25] ? _GEN6978 : _GEN6971;
wire  _GEN6980 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6981 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6982 = io_x[9] ? _GEN6981 : _GEN6980;
wire  _GEN6983 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6984 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6985 = io_x[9] ? _GEN6984 : _GEN6983;
wire  _GEN6986 = io_x[23] ? _GEN6985 : _GEN6982;
wire  _GEN6987 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6988 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6989 = io_x[9] ? _GEN6988 : _GEN6987;
wire  _GEN6990 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6991 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6992 = io_x[9] ? _GEN6991 : _GEN6990;
wire  _GEN6993 = io_x[23] ? _GEN6992 : _GEN6989;
wire  _GEN6994 = io_x[25] ? _GEN6993 : _GEN6986;
wire  _GEN6995 = io_x[5] ? _GEN6994 : _GEN6979;
wire  _GEN6996 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN6997 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN6998 = io_x[9] ? _GEN6997 : _GEN6996;
wire  _GEN6999 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN7000 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN7001 = io_x[9] ? _GEN7000 : _GEN6999;
wire  _GEN7002 = io_x[23] ? _GEN7001 : _GEN6998;
wire  _GEN7003 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN7004 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN7005 = io_x[9] ? _GEN7004 : _GEN7003;
wire  _GEN7006 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN7007 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN7008 = io_x[9] ? _GEN7007 : _GEN7006;
wire  _GEN7009 = io_x[23] ? _GEN7008 : _GEN7005;
wire  _GEN7010 = io_x[25] ? _GEN7009 : _GEN7002;
wire  _GEN7011 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN7012 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN7013 = io_x[9] ? _GEN7012 : _GEN7011;
wire  _GEN7014 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN7015 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN7016 = io_x[9] ? _GEN7015 : _GEN7014;
wire  _GEN7017 = io_x[23] ? _GEN7016 : _GEN7013;
wire  _GEN7018 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN7019 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN7020 = io_x[9] ? _GEN7019 : _GEN7018;
wire  _GEN7021 = io_x[1] ? _GEN6774 : _GEN6775;
wire  _GEN7022 = io_x[1] ? _GEN6775 : _GEN6774;
wire  _GEN7023 = io_x[9] ? _GEN7022 : _GEN7021;
wire  _GEN7024 = io_x[23] ? _GEN7023 : _GEN7020;
wire  _GEN7025 = io_x[25] ? _GEN7024 : _GEN7017;
wire  _GEN7026 = io_x[5] ? _GEN7025 : _GEN7010;
wire  _GEN7027 = io_x[21] ? _GEN7026 : _GEN6995;
wire  _GEN7028 = io_x[13] ? _GEN7027 : _GEN6964;
wire  _GEN7029 = io_x[29] ? _GEN7028 : _GEN6902;
assign io_y[7] = _GEN7029;
wire  _GEN7030 = 1'b0;
wire  _GEN7031 = 1'b1;
wire  _GEN7032 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7033 = 1'b0;
wire  _GEN7034 = io_x[8] ? _GEN7033 : _GEN7032;
wire  _GEN7035 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7036 = io_x[8] ? _GEN7035 : _GEN7033;
wire  _GEN7037 = io_x[24] ? _GEN7036 : _GEN7034;
wire  _GEN7038 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7039 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7040 = io_x[8] ? _GEN7039 : _GEN7038;
wire  _GEN7041 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7042 = io_x[8] ? _GEN7041 : _GEN7033;
wire  _GEN7043 = io_x[24] ? _GEN7042 : _GEN7040;
wire  _GEN7044 = io_x[3] ? _GEN7043 : _GEN7037;
wire  _GEN7045 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7046 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7047 = io_x[8] ? _GEN7046 : _GEN7045;
wire  _GEN7048 = 1'b1;
wire  _GEN7049 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7050 = io_x[8] ? _GEN7049 : _GEN7048;
wire  _GEN7051 = io_x[24] ? _GEN7050 : _GEN7047;
wire  _GEN7052 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7053 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7054 = io_x[8] ? _GEN7053 : _GEN7052;
wire  _GEN7055 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7056 = io_x[8] ? _GEN7055 : _GEN7048;
wire  _GEN7057 = io_x[24] ? _GEN7056 : _GEN7054;
wire  _GEN7058 = io_x[3] ? _GEN7057 : _GEN7051;
wire  _GEN7059 = io_x[5] ? _GEN7058 : _GEN7044;
wire  _GEN7060 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7061 = io_x[8] ? _GEN7033 : _GEN7060;
wire  _GEN7062 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7063 = io_x[8] ? _GEN7048 : _GEN7062;
wire  _GEN7064 = io_x[24] ? _GEN7063 : _GEN7061;
wire  _GEN7065 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7066 = io_x[8] ? _GEN7065 : _GEN7033;
wire  _GEN7067 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7068 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7069 = io_x[8] ? _GEN7068 : _GEN7067;
wire  _GEN7070 = io_x[24] ? _GEN7069 : _GEN7066;
wire  _GEN7071 = io_x[3] ? _GEN7070 : _GEN7064;
wire  _GEN7072 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7073 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7074 = io_x[8] ? _GEN7073 : _GEN7072;
wire  _GEN7075 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7076 = io_x[8] ? _GEN7033 : _GEN7075;
wire  _GEN7077 = io_x[24] ? _GEN7076 : _GEN7074;
wire  _GEN7078 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7079 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7080 = io_x[8] ? _GEN7079 : _GEN7078;
wire  _GEN7081 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7082 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7083 = io_x[8] ? _GEN7082 : _GEN7081;
wire  _GEN7084 = io_x[24] ? _GEN7083 : _GEN7080;
wire  _GEN7085 = io_x[3] ? _GEN7084 : _GEN7077;
wire  _GEN7086 = io_x[5] ? _GEN7085 : _GEN7071;
wire  _GEN7087 = io_x[7] ? _GEN7086 : _GEN7059;
wire  _GEN7088 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7089 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7090 = io_x[8] ? _GEN7089 : _GEN7088;
wire  _GEN7091 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7092 = io_x[8] ? _GEN7048 : _GEN7091;
wire  _GEN7093 = io_x[24] ? _GEN7092 : _GEN7090;
wire  _GEN7094 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7095 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7096 = io_x[8] ? _GEN7095 : _GEN7094;
wire  _GEN7097 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7098 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7099 = io_x[8] ? _GEN7098 : _GEN7097;
wire  _GEN7100 = io_x[24] ? _GEN7099 : _GEN7096;
wire  _GEN7101 = io_x[3] ? _GEN7100 : _GEN7093;
wire  _GEN7102 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7103 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7104 = io_x[8] ? _GEN7103 : _GEN7102;
wire  _GEN7105 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7106 = io_x[8] ? _GEN7105 : _GEN7048;
wire  _GEN7107 = io_x[24] ? _GEN7106 : _GEN7104;
wire  _GEN7108 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7109 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7110 = io_x[8] ? _GEN7109 : _GEN7108;
wire  _GEN7111 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7112 = io_x[8] ? _GEN7111 : _GEN7048;
wire  _GEN7113 = io_x[24] ? _GEN7112 : _GEN7110;
wire  _GEN7114 = io_x[3] ? _GEN7113 : _GEN7107;
wire  _GEN7115 = io_x[5] ? _GEN7114 : _GEN7101;
wire  _GEN7116 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7117 = io_x[8] ? _GEN7116 : _GEN7033;
wire  _GEN7118 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7119 = io_x[8] ? _GEN7048 : _GEN7118;
wire  _GEN7120 = io_x[24] ? _GEN7119 : _GEN7117;
wire  _GEN7121 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7122 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7123 = io_x[8] ? _GEN7122 : _GEN7121;
wire  _GEN7124 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7125 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7126 = io_x[8] ? _GEN7125 : _GEN7124;
wire  _GEN7127 = io_x[24] ? _GEN7126 : _GEN7123;
wire  _GEN7128 = io_x[3] ? _GEN7127 : _GEN7120;
wire  _GEN7129 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7130 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7131 = io_x[8] ? _GEN7130 : _GEN7129;
wire  _GEN7132 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7133 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7134 = io_x[8] ? _GEN7133 : _GEN7132;
wire  _GEN7135 = io_x[24] ? _GEN7134 : _GEN7131;
wire  _GEN7136 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7137 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7138 = io_x[8] ? _GEN7137 : _GEN7136;
wire  _GEN7139 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7140 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7141 = io_x[8] ? _GEN7140 : _GEN7139;
wire  _GEN7142 = io_x[24] ? _GEN7141 : _GEN7138;
wire  _GEN7143 = io_x[3] ? _GEN7142 : _GEN7135;
wire  _GEN7144 = io_x[5] ? _GEN7143 : _GEN7128;
wire  _GEN7145 = io_x[7] ? _GEN7144 : _GEN7115;
wire  _GEN7146 = io_x[9] ? _GEN7145 : _GEN7087;
wire  _GEN7147 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7148 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7149 = io_x[8] ? _GEN7148 : _GEN7147;
wire  _GEN7150 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7151 = io_x[8] ? _GEN7033 : _GEN7150;
wire  _GEN7152 = io_x[24] ? _GEN7151 : _GEN7149;
wire  _GEN7153 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7154 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7155 = io_x[8] ? _GEN7154 : _GEN7153;
wire  _GEN7156 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7157 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7158 = io_x[8] ? _GEN7157 : _GEN7156;
wire  _GEN7159 = io_x[24] ? _GEN7158 : _GEN7155;
wire  _GEN7160 = io_x[3] ? _GEN7159 : _GEN7152;
wire  _GEN7161 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7162 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7163 = io_x[8] ? _GEN7162 : _GEN7161;
wire  _GEN7164 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7165 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7166 = io_x[8] ? _GEN7165 : _GEN7164;
wire  _GEN7167 = io_x[24] ? _GEN7166 : _GEN7163;
wire  _GEN7168 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7169 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7170 = io_x[8] ? _GEN7169 : _GEN7168;
wire  _GEN7171 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7172 = io_x[8] ? _GEN7171 : _GEN7048;
wire  _GEN7173 = io_x[24] ? _GEN7172 : _GEN7170;
wire  _GEN7174 = io_x[3] ? _GEN7173 : _GEN7167;
wire  _GEN7175 = io_x[5] ? _GEN7174 : _GEN7160;
wire  _GEN7176 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7177 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7178 = io_x[8] ? _GEN7177 : _GEN7176;
wire  _GEN7179 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7180 = io_x[8] ? _GEN7033 : _GEN7179;
wire  _GEN7181 = io_x[24] ? _GEN7180 : _GEN7178;
wire  _GEN7182 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7183 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7184 = io_x[8] ? _GEN7183 : _GEN7182;
wire  _GEN7185 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7186 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7187 = io_x[8] ? _GEN7186 : _GEN7185;
wire  _GEN7188 = io_x[24] ? _GEN7187 : _GEN7184;
wire  _GEN7189 = io_x[3] ? _GEN7188 : _GEN7181;
wire  _GEN7190 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7191 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7192 = io_x[8] ? _GEN7191 : _GEN7190;
wire  _GEN7193 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7194 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7195 = io_x[8] ? _GEN7194 : _GEN7193;
wire  _GEN7196 = io_x[24] ? _GEN7195 : _GEN7192;
wire  _GEN7197 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7198 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7199 = io_x[8] ? _GEN7198 : _GEN7197;
wire  _GEN7200 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7201 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7202 = io_x[8] ? _GEN7201 : _GEN7200;
wire  _GEN7203 = io_x[24] ? _GEN7202 : _GEN7199;
wire  _GEN7204 = io_x[3] ? _GEN7203 : _GEN7196;
wire  _GEN7205 = io_x[5] ? _GEN7204 : _GEN7189;
wire  _GEN7206 = io_x[7] ? _GEN7205 : _GEN7175;
wire  _GEN7207 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7208 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7209 = io_x[8] ? _GEN7208 : _GEN7207;
wire  _GEN7210 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7211 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7212 = io_x[8] ? _GEN7211 : _GEN7210;
wire  _GEN7213 = io_x[24] ? _GEN7212 : _GEN7209;
wire  _GEN7214 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7215 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7216 = io_x[8] ? _GEN7215 : _GEN7214;
wire  _GEN7217 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7218 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7219 = io_x[8] ? _GEN7218 : _GEN7217;
wire  _GEN7220 = io_x[24] ? _GEN7219 : _GEN7216;
wire  _GEN7221 = io_x[3] ? _GEN7220 : _GEN7213;
wire  _GEN7222 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7223 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7224 = io_x[8] ? _GEN7223 : _GEN7222;
wire  _GEN7225 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7226 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7227 = io_x[8] ? _GEN7226 : _GEN7225;
wire  _GEN7228 = io_x[24] ? _GEN7227 : _GEN7224;
wire  _GEN7229 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7230 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7231 = io_x[8] ? _GEN7230 : _GEN7229;
wire  _GEN7232 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7233 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7234 = io_x[8] ? _GEN7233 : _GEN7232;
wire  _GEN7235 = io_x[24] ? _GEN7234 : _GEN7231;
wire  _GEN7236 = io_x[3] ? _GEN7235 : _GEN7228;
wire  _GEN7237 = io_x[5] ? _GEN7236 : _GEN7221;
wire  _GEN7238 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7239 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7240 = io_x[8] ? _GEN7239 : _GEN7238;
wire  _GEN7241 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7242 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7243 = io_x[8] ? _GEN7242 : _GEN7241;
wire  _GEN7244 = io_x[24] ? _GEN7243 : _GEN7240;
wire  _GEN7245 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7246 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7247 = io_x[8] ? _GEN7246 : _GEN7245;
wire  _GEN7248 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7249 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7250 = io_x[8] ? _GEN7249 : _GEN7248;
wire  _GEN7251 = io_x[24] ? _GEN7250 : _GEN7247;
wire  _GEN7252 = io_x[3] ? _GEN7251 : _GEN7244;
wire  _GEN7253 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7254 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7255 = io_x[8] ? _GEN7254 : _GEN7253;
wire  _GEN7256 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7257 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7258 = io_x[8] ? _GEN7257 : _GEN7256;
wire  _GEN7259 = io_x[24] ? _GEN7258 : _GEN7255;
wire  _GEN7260 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7261 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7262 = io_x[8] ? _GEN7261 : _GEN7260;
wire  _GEN7263 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7264 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7265 = io_x[8] ? _GEN7264 : _GEN7263;
wire  _GEN7266 = io_x[24] ? _GEN7265 : _GEN7262;
wire  _GEN7267 = io_x[3] ? _GEN7266 : _GEN7259;
wire  _GEN7268 = io_x[5] ? _GEN7267 : _GEN7252;
wire  _GEN7269 = io_x[7] ? _GEN7268 : _GEN7237;
wire  _GEN7270 = io_x[9] ? _GEN7269 : _GEN7206;
wire  _GEN7271 = io_x[0] ? _GEN7270 : _GEN7146;
wire  _GEN7272 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7273 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7274 = io_x[8] ? _GEN7273 : _GEN7272;
wire  _GEN7275 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7276 = io_x[8] ? _GEN7275 : _GEN7048;
wire  _GEN7277 = io_x[24] ? _GEN7276 : _GEN7274;
wire  _GEN7278 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7279 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7280 = io_x[8] ? _GEN7279 : _GEN7278;
wire  _GEN7281 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7282 = io_x[8] ? _GEN7281 : _GEN7048;
wire  _GEN7283 = io_x[24] ? _GEN7282 : _GEN7280;
wire  _GEN7284 = io_x[3] ? _GEN7283 : _GEN7277;
wire  _GEN7285 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7286 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7287 = io_x[8] ? _GEN7286 : _GEN7285;
wire  _GEN7288 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7289 = io_x[8] ? _GEN7288 : _GEN7048;
wire  _GEN7290 = io_x[24] ? _GEN7289 : _GEN7287;
wire  _GEN7291 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7292 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7293 = io_x[8] ? _GEN7292 : _GEN7291;
wire  _GEN7294 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7295 = io_x[8] ? _GEN7294 : _GEN7048;
wire  _GEN7296 = io_x[24] ? _GEN7295 : _GEN7293;
wire  _GEN7297 = io_x[3] ? _GEN7296 : _GEN7290;
wire  _GEN7298 = io_x[5] ? _GEN7297 : _GEN7284;
wire  _GEN7299 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7300 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7301 = io_x[8] ? _GEN7300 : _GEN7299;
wire  _GEN7302 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7303 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7304 = io_x[8] ? _GEN7303 : _GEN7302;
wire  _GEN7305 = io_x[24] ? _GEN7304 : _GEN7301;
wire  _GEN7306 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7307 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7308 = io_x[8] ? _GEN7307 : _GEN7306;
wire  _GEN7309 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7310 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7311 = io_x[8] ? _GEN7310 : _GEN7309;
wire  _GEN7312 = io_x[24] ? _GEN7311 : _GEN7308;
wire  _GEN7313 = io_x[3] ? _GEN7312 : _GEN7305;
wire  _GEN7314 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7315 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7316 = io_x[8] ? _GEN7315 : _GEN7314;
wire  _GEN7317 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7318 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7319 = io_x[8] ? _GEN7318 : _GEN7317;
wire  _GEN7320 = io_x[24] ? _GEN7319 : _GEN7316;
wire  _GEN7321 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7322 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7323 = io_x[8] ? _GEN7322 : _GEN7321;
wire  _GEN7324 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7325 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7326 = io_x[8] ? _GEN7325 : _GEN7324;
wire  _GEN7327 = io_x[24] ? _GEN7326 : _GEN7323;
wire  _GEN7328 = io_x[3] ? _GEN7327 : _GEN7320;
wire  _GEN7329 = io_x[5] ? _GEN7328 : _GEN7313;
wire  _GEN7330 = io_x[7] ? _GEN7329 : _GEN7298;
wire  _GEN7331 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7332 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7333 = io_x[8] ? _GEN7332 : _GEN7331;
wire  _GEN7334 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7335 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7336 = io_x[8] ? _GEN7335 : _GEN7334;
wire  _GEN7337 = io_x[24] ? _GEN7336 : _GEN7333;
wire  _GEN7338 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7339 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7340 = io_x[8] ? _GEN7339 : _GEN7338;
wire  _GEN7341 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7342 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7343 = io_x[8] ? _GEN7342 : _GEN7341;
wire  _GEN7344 = io_x[24] ? _GEN7343 : _GEN7340;
wire  _GEN7345 = io_x[3] ? _GEN7344 : _GEN7337;
wire  _GEN7346 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7347 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7348 = io_x[8] ? _GEN7347 : _GEN7346;
wire  _GEN7349 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7350 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7351 = io_x[8] ? _GEN7350 : _GEN7349;
wire  _GEN7352 = io_x[24] ? _GEN7351 : _GEN7348;
wire  _GEN7353 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7354 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7355 = io_x[8] ? _GEN7354 : _GEN7353;
wire  _GEN7356 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7357 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7358 = io_x[8] ? _GEN7357 : _GEN7356;
wire  _GEN7359 = io_x[24] ? _GEN7358 : _GEN7355;
wire  _GEN7360 = io_x[3] ? _GEN7359 : _GEN7352;
wire  _GEN7361 = io_x[5] ? _GEN7360 : _GEN7345;
wire  _GEN7362 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7363 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7364 = io_x[8] ? _GEN7363 : _GEN7362;
wire  _GEN7365 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7366 = io_x[8] ? _GEN7365 : _GEN7048;
wire  _GEN7367 = io_x[24] ? _GEN7366 : _GEN7364;
wire  _GEN7368 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7369 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7370 = io_x[8] ? _GEN7369 : _GEN7368;
wire  _GEN7371 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7372 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7373 = io_x[8] ? _GEN7372 : _GEN7371;
wire  _GEN7374 = io_x[24] ? _GEN7373 : _GEN7370;
wire  _GEN7375 = io_x[3] ? _GEN7374 : _GEN7367;
wire  _GEN7376 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7377 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7378 = io_x[8] ? _GEN7377 : _GEN7376;
wire  _GEN7379 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7380 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7381 = io_x[8] ? _GEN7380 : _GEN7379;
wire  _GEN7382 = io_x[24] ? _GEN7381 : _GEN7378;
wire  _GEN7383 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7384 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7385 = io_x[8] ? _GEN7384 : _GEN7383;
wire  _GEN7386 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7387 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7388 = io_x[8] ? _GEN7387 : _GEN7386;
wire  _GEN7389 = io_x[24] ? _GEN7388 : _GEN7385;
wire  _GEN7390 = io_x[3] ? _GEN7389 : _GEN7382;
wire  _GEN7391 = io_x[5] ? _GEN7390 : _GEN7375;
wire  _GEN7392 = io_x[7] ? _GEN7391 : _GEN7361;
wire  _GEN7393 = io_x[9] ? _GEN7392 : _GEN7330;
wire  _GEN7394 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7395 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7396 = io_x[8] ? _GEN7395 : _GEN7394;
wire  _GEN7397 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7398 = io_x[8] ? _GEN7397 : _GEN7033;
wire  _GEN7399 = io_x[24] ? _GEN7398 : _GEN7396;
wire  _GEN7400 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7401 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7402 = io_x[8] ? _GEN7401 : _GEN7400;
wire  _GEN7403 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7404 = io_x[8] ? _GEN7403 : _GEN7048;
wire  _GEN7405 = io_x[24] ? _GEN7404 : _GEN7402;
wire  _GEN7406 = io_x[3] ? _GEN7405 : _GEN7399;
wire  _GEN7407 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7408 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7409 = io_x[8] ? _GEN7408 : _GEN7407;
wire  _GEN7410 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7411 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7412 = io_x[8] ? _GEN7411 : _GEN7410;
wire  _GEN7413 = io_x[24] ? _GEN7412 : _GEN7409;
wire  _GEN7414 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7415 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7416 = io_x[8] ? _GEN7415 : _GEN7414;
wire  _GEN7417 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7418 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7419 = io_x[8] ? _GEN7418 : _GEN7417;
wire  _GEN7420 = io_x[24] ? _GEN7419 : _GEN7416;
wire  _GEN7421 = io_x[3] ? _GEN7420 : _GEN7413;
wire  _GEN7422 = io_x[5] ? _GEN7421 : _GEN7406;
wire  _GEN7423 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7424 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7425 = io_x[8] ? _GEN7424 : _GEN7423;
wire  _GEN7426 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7427 = io_x[8] ? _GEN7048 : _GEN7426;
wire  _GEN7428 = io_x[24] ? _GEN7427 : _GEN7425;
wire  _GEN7429 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7430 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7431 = io_x[8] ? _GEN7430 : _GEN7429;
wire  _GEN7432 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7433 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7434 = io_x[8] ? _GEN7433 : _GEN7432;
wire  _GEN7435 = io_x[24] ? _GEN7434 : _GEN7431;
wire  _GEN7436 = io_x[3] ? _GEN7435 : _GEN7428;
wire  _GEN7437 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7438 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7439 = io_x[8] ? _GEN7438 : _GEN7437;
wire  _GEN7440 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7441 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7442 = io_x[8] ? _GEN7441 : _GEN7440;
wire  _GEN7443 = io_x[24] ? _GEN7442 : _GEN7439;
wire  _GEN7444 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7445 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7446 = io_x[8] ? _GEN7445 : _GEN7444;
wire  _GEN7447 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7448 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7449 = io_x[8] ? _GEN7448 : _GEN7447;
wire  _GEN7450 = io_x[24] ? _GEN7449 : _GEN7446;
wire  _GEN7451 = io_x[3] ? _GEN7450 : _GEN7443;
wire  _GEN7452 = io_x[5] ? _GEN7451 : _GEN7436;
wire  _GEN7453 = io_x[7] ? _GEN7452 : _GEN7422;
wire  _GEN7454 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7455 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7456 = io_x[8] ? _GEN7455 : _GEN7454;
wire  _GEN7457 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7458 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7459 = io_x[8] ? _GEN7458 : _GEN7457;
wire  _GEN7460 = io_x[24] ? _GEN7459 : _GEN7456;
wire  _GEN7461 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7462 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7463 = io_x[8] ? _GEN7462 : _GEN7461;
wire  _GEN7464 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7465 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7466 = io_x[8] ? _GEN7465 : _GEN7464;
wire  _GEN7467 = io_x[24] ? _GEN7466 : _GEN7463;
wire  _GEN7468 = io_x[3] ? _GEN7467 : _GEN7460;
wire  _GEN7469 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7470 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7471 = io_x[8] ? _GEN7470 : _GEN7469;
wire  _GEN7472 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7473 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7474 = io_x[8] ? _GEN7473 : _GEN7472;
wire  _GEN7475 = io_x[24] ? _GEN7474 : _GEN7471;
wire  _GEN7476 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7477 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7478 = io_x[8] ? _GEN7477 : _GEN7476;
wire  _GEN7479 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7480 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7481 = io_x[8] ? _GEN7480 : _GEN7479;
wire  _GEN7482 = io_x[24] ? _GEN7481 : _GEN7478;
wire  _GEN7483 = io_x[3] ? _GEN7482 : _GEN7475;
wire  _GEN7484 = io_x[5] ? _GEN7483 : _GEN7468;
wire  _GEN7485 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7486 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7487 = io_x[8] ? _GEN7486 : _GEN7485;
wire  _GEN7488 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7489 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7490 = io_x[8] ? _GEN7489 : _GEN7488;
wire  _GEN7491 = io_x[24] ? _GEN7490 : _GEN7487;
wire  _GEN7492 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7493 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7494 = io_x[8] ? _GEN7493 : _GEN7492;
wire  _GEN7495 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7496 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7497 = io_x[8] ? _GEN7496 : _GEN7495;
wire  _GEN7498 = io_x[24] ? _GEN7497 : _GEN7494;
wire  _GEN7499 = io_x[3] ? _GEN7498 : _GEN7491;
wire  _GEN7500 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7501 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7502 = io_x[8] ? _GEN7501 : _GEN7500;
wire  _GEN7503 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7504 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7505 = io_x[8] ? _GEN7504 : _GEN7503;
wire  _GEN7506 = io_x[24] ? _GEN7505 : _GEN7502;
wire  _GEN7507 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7508 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7509 = io_x[8] ? _GEN7508 : _GEN7507;
wire  _GEN7510 = io_x[4] ? _GEN7030 : _GEN7031;
wire  _GEN7511 = io_x[4] ? _GEN7031 : _GEN7030;
wire  _GEN7512 = io_x[8] ? _GEN7511 : _GEN7510;
wire  _GEN7513 = io_x[24] ? _GEN7512 : _GEN7509;
wire  _GEN7514 = io_x[3] ? _GEN7513 : _GEN7506;
wire  _GEN7515 = io_x[5] ? _GEN7514 : _GEN7499;
wire  _GEN7516 = io_x[7] ? _GEN7515 : _GEN7484;
wire  _GEN7517 = io_x[9] ? _GEN7516 : _GEN7453;
wire  _GEN7518 = io_x[0] ? _GEN7517 : _GEN7393;
wire  _GEN7519 = io_x[12] ? _GEN7518 : _GEN7271;
assign io_y[6] = _GEN7519;
wire  _GEN7520 = 1'b0;
wire  _GEN7521 = 1'b1;
wire  _GEN7522 = 1'b0;
wire  _GEN7523 = 1'b1;
wire  _GEN7524 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7525 = io_x[11] ? _GEN7524 : _GEN7521;
wire  _GEN7526 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7527 = io_x[11] ? _GEN7526 : _GEN7521;
wire  _GEN7528 = io_x[9] ? _GEN7527 : _GEN7525;
wire  _GEN7529 = io_x[21] ? _GEN7528 : _GEN7520;
wire  _GEN7530 = 1'b0;
wire  _GEN7531 = 1'b0;
wire  _GEN7532 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7533 = io_x[11] ? _GEN7532 : _GEN7531;
wire  _GEN7534 = io_x[9] ? _GEN7533 : _GEN7530;
wire  _GEN7535 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7536 = io_x[11] ? _GEN7535 : _GEN7521;
wire  _GEN7537 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7538 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7539 = io_x[11] ? _GEN7538 : _GEN7537;
wire  _GEN7540 = io_x[9] ? _GEN7539 : _GEN7536;
wire  _GEN7541 = io_x[21] ? _GEN7540 : _GEN7534;
wire  _GEN7542 = io_x[31] ? _GEN7541 : _GEN7529;
wire  _GEN7543 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7544 = io_x[11] ? _GEN7543 : _GEN7531;
wire  _GEN7545 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7546 = io_x[11] ? _GEN7531 : _GEN7545;
wire  _GEN7547 = io_x[9] ? _GEN7546 : _GEN7544;
wire  _GEN7548 = 1'b1;
wire  _GEN7549 = io_x[11] ? _GEN7521 : _GEN7531;
wire  _GEN7550 = io_x[9] ? _GEN7549 : _GEN7548;
wire  _GEN7551 = io_x[21] ? _GEN7550 : _GEN7547;
wire  _GEN7552 = 1'b1;
wire  _GEN7553 = io_x[31] ? _GEN7552 : _GEN7551;
wire  _GEN7554 = io_x[30] ? _GEN7553 : _GEN7542;
wire  _GEN7555 = io_x[11] ? _GEN7521 : _GEN7531;
wire  _GEN7556 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7557 = io_x[11] ? _GEN7556 : _GEN7521;
wire  _GEN7558 = io_x[9] ? _GEN7557 : _GEN7555;
wire  _GEN7559 = 1'b1;
wire  _GEN7560 = io_x[21] ? _GEN7559 : _GEN7558;
wire  _GEN7561 = 1'b0;
wire  _GEN7562 = io_x[31] ? _GEN7561 : _GEN7560;
wire  _GEN7563 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7564 = io_x[11] ? _GEN7563 : _GEN7521;
wire  _GEN7565 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7566 = io_x[11] ? _GEN7565 : _GEN7531;
wire  _GEN7567 = io_x[9] ? _GEN7566 : _GEN7564;
wire  _GEN7568 = io_x[21] ? _GEN7520 : _GEN7567;
wire  _GEN7569 = io_x[31] ? _GEN7552 : _GEN7568;
wire  _GEN7570 = io_x[30] ? _GEN7569 : _GEN7562;
wire  _GEN7571 = io_x[29] ? _GEN7570 : _GEN7554;
wire  _GEN7572 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7573 = io_x[11] ? _GEN7572 : _GEN7521;
wire  _GEN7574 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7575 = io_x[11] ? _GEN7574 : _GEN7521;
wire  _GEN7576 = io_x[9] ? _GEN7575 : _GEN7573;
wire  _GEN7577 = io_x[21] ? _GEN7576 : _GEN7520;
wire  _GEN7578 = io_x[31] ? _GEN7552 : _GEN7577;
wire  _GEN7579 = 1'b1;
wire  _GEN7580 = io_x[30] ? _GEN7579 : _GEN7578;
wire  _GEN7581 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7582 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7583 = io_x[11] ? _GEN7582 : _GEN7581;
wire  _GEN7584 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7585 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7586 = io_x[11] ? _GEN7585 : _GEN7584;
wire  _GEN7587 = io_x[9] ? _GEN7586 : _GEN7583;
wire  _GEN7588 = io_x[21] ? _GEN7520 : _GEN7587;
wire  _GEN7589 = io_x[31] ? _GEN7552 : _GEN7588;
wire  _GEN7590 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7591 = io_x[11] ? _GEN7531 : _GEN7590;
wire  _GEN7592 = io_x[9] ? _GEN7530 : _GEN7591;
wire  _GEN7593 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7594 = io_x[11] ? _GEN7521 : _GEN7593;
wire  _GEN7595 = io_x[9] ? _GEN7548 : _GEN7594;
wire  _GEN7596 = io_x[21] ? _GEN7595 : _GEN7592;
wire  _GEN7597 = io_x[31] ? _GEN7552 : _GEN7596;
wire  _GEN7598 = io_x[30] ? _GEN7597 : _GEN7589;
wire  _GEN7599 = io_x[29] ? _GEN7598 : _GEN7580;
wire  _GEN7600 = io_x[28] ? _GEN7599 : _GEN7571;
wire  _GEN7601 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7602 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7603 = io_x[11] ? _GEN7602 : _GEN7601;
wire  _GEN7604 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7605 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7606 = io_x[11] ? _GEN7605 : _GEN7604;
wire  _GEN7607 = io_x[9] ? _GEN7606 : _GEN7603;
wire  _GEN7608 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7609 = io_x[11] ? _GEN7521 : _GEN7608;
wire  _GEN7610 = io_x[9] ? _GEN7609 : _GEN7548;
wire  _GEN7611 = io_x[21] ? _GEN7610 : _GEN7607;
wire  _GEN7612 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7613 = io_x[11] ? _GEN7612 : _GEN7531;
wire  _GEN7614 = io_x[9] ? _GEN7613 : _GEN7530;
wire  _GEN7615 = io_x[21] ? _GEN7520 : _GEN7614;
wire  _GEN7616 = io_x[31] ? _GEN7615 : _GEN7611;
wire  _GEN7617 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7618 = io_x[11] ? _GEN7617 : _GEN7521;
wire  _GEN7619 = io_x[9] ? _GEN7618 : _GEN7548;
wire  _GEN7620 = io_x[21] ? _GEN7559 : _GEN7619;
wire  _GEN7621 = io_x[31] ? _GEN7552 : _GEN7620;
wire  _GEN7622 = io_x[30] ? _GEN7621 : _GEN7616;
wire  _GEN7623 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7624 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7625 = io_x[11] ? _GEN7624 : _GEN7623;
wire  _GEN7626 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7627 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7628 = io_x[11] ? _GEN7627 : _GEN7626;
wire  _GEN7629 = io_x[9] ? _GEN7628 : _GEN7625;
wire  _GEN7630 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7631 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7632 = io_x[11] ? _GEN7631 : _GEN7630;
wire  _GEN7633 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7634 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7635 = io_x[11] ? _GEN7634 : _GEN7633;
wire  _GEN7636 = io_x[9] ? _GEN7635 : _GEN7632;
wire  _GEN7637 = io_x[21] ? _GEN7636 : _GEN7629;
wire  _GEN7638 = io_x[31] ? _GEN7561 : _GEN7637;
wire  _GEN7639 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7640 = io_x[11] ? _GEN7639 : _GEN7521;
wire  _GEN7641 = io_x[9] ? _GEN7640 : _GEN7530;
wire  _GEN7642 = io_x[21] ? _GEN7641 : _GEN7520;
wire  _GEN7643 = io_x[31] ? _GEN7552 : _GEN7642;
wire  _GEN7644 = io_x[30] ? _GEN7643 : _GEN7638;
wire  _GEN7645 = io_x[29] ? _GEN7644 : _GEN7622;
wire  _GEN7646 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7647 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7648 = io_x[11] ? _GEN7647 : _GEN7646;
wire  _GEN7649 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7650 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7651 = io_x[11] ? _GEN7650 : _GEN7649;
wire  _GEN7652 = io_x[9] ? _GEN7651 : _GEN7648;
wire  _GEN7653 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7654 = io_x[11] ? _GEN7653 : _GEN7521;
wire  _GEN7655 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7656 = io_x[11] ? _GEN7655 : _GEN7531;
wire  _GEN7657 = io_x[9] ? _GEN7656 : _GEN7654;
wire  _GEN7658 = io_x[21] ? _GEN7657 : _GEN7652;
wire  _GEN7659 = io_x[11] ? _GEN7531 : _GEN7521;
wire  _GEN7660 = io_x[9] ? _GEN7548 : _GEN7659;
wire  _GEN7661 = io_x[21] ? _GEN7660 : _GEN7520;
wire  _GEN7662 = io_x[31] ? _GEN7661 : _GEN7658;
wire  _GEN7663 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7664 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7665 = io_x[11] ? _GEN7664 : _GEN7663;
wire  _GEN7666 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7667 = io_x[11] ? _GEN7531 : _GEN7666;
wire  _GEN7668 = io_x[9] ? _GEN7667 : _GEN7665;
wire  _GEN7669 = io_x[21] ? _GEN7559 : _GEN7668;
wire  _GEN7670 = io_x[31] ? _GEN7552 : _GEN7669;
wire  _GEN7671 = io_x[30] ? _GEN7670 : _GEN7662;
wire  _GEN7672 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7673 = io_x[11] ? _GEN7672 : _GEN7521;
wire  _GEN7674 = io_x[9] ? _GEN7673 : _GEN7548;
wire  _GEN7675 = io_x[21] ? _GEN7520 : _GEN7674;
wire  _GEN7676 = io_x[31] ? _GEN7552 : _GEN7675;
wire  _GEN7677 = io_x[11] ? _GEN7521 : _GEN7531;
wire  _GEN7678 = io_x[9] ? _GEN7677 : _GEN7548;
wire  _GEN7679 = io_x[21] ? _GEN7520 : _GEN7678;
wire  _GEN7680 = io_x[31] ? _GEN7552 : _GEN7679;
wire  _GEN7681 = io_x[30] ? _GEN7680 : _GEN7676;
wire  _GEN7682 = io_x[29] ? _GEN7681 : _GEN7671;
wire  _GEN7683 = io_x[28] ? _GEN7682 : _GEN7645;
wire  _GEN7684 = io_x[27] ? _GEN7683 : _GEN7600;
wire  _GEN7685 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7686 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7687 = io_x[11] ? _GEN7686 : _GEN7685;
wire  _GEN7688 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7689 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7690 = io_x[11] ? _GEN7689 : _GEN7688;
wire  _GEN7691 = io_x[9] ? _GEN7690 : _GEN7687;
wire  _GEN7692 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7693 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7694 = io_x[11] ? _GEN7693 : _GEN7692;
wire  _GEN7695 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7696 = io_x[11] ? _GEN7695 : _GEN7521;
wire  _GEN7697 = io_x[9] ? _GEN7696 : _GEN7694;
wire  _GEN7698 = io_x[21] ? _GEN7697 : _GEN7691;
wire  _GEN7699 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7700 = io_x[11] ? _GEN7531 : _GEN7699;
wire  _GEN7701 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7702 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7703 = io_x[11] ? _GEN7702 : _GEN7701;
wire  _GEN7704 = io_x[9] ? _GEN7703 : _GEN7700;
wire  _GEN7705 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7706 = io_x[11] ? _GEN7705 : _GEN7531;
wire  _GEN7707 = io_x[9] ? _GEN7706 : _GEN7530;
wire  _GEN7708 = io_x[21] ? _GEN7707 : _GEN7704;
wire  _GEN7709 = io_x[31] ? _GEN7708 : _GEN7698;
wire  _GEN7710 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7711 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7712 = io_x[11] ? _GEN7711 : _GEN7710;
wire  _GEN7713 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7714 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7715 = io_x[11] ? _GEN7714 : _GEN7713;
wire  _GEN7716 = io_x[9] ? _GEN7715 : _GEN7712;
wire  _GEN7717 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7718 = io_x[11] ? _GEN7717 : _GEN7521;
wire  _GEN7719 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7720 = io_x[11] ? _GEN7531 : _GEN7719;
wire  _GEN7721 = io_x[9] ? _GEN7720 : _GEN7718;
wire  _GEN7722 = io_x[21] ? _GEN7721 : _GEN7716;
wire  _GEN7723 = io_x[31] ? _GEN7552 : _GEN7722;
wire  _GEN7724 = io_x[30] ? _GEN7723 : _GEN7709;
wire  _GEN7725 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7726 = io_x[11] ? _GEN7725 : _GEN7531;
wire  _GEN7727 = io_x[9] ? _GEN7726 : _GEN7530;
wire  _GEN7728 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7729 = io_x[11] ? _GEN7728 : _GEN7521;
wire  _GEN7730 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7731 = io_x[11] ? _GEN7730 : _GEN7521;
wire  _GEN7732 = io_x[9] ? _GEN7731 : _GEN7729;
wire  _GEN7733 = io_x[21] ? _GEN7732 : _GEN7727;
wire  _GEN7734 = io_x[31] ? _GEN7561 : _GEN7733;
wire  _GEN7735 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7736 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7737 = io_x[11] ? _GEN7736 : _GEN7735;
wire  _GEN7738 = io_x[9] ? _GEN7530 : _GEN7737;
wire  _GEN7739 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7740 = io_x[11] ? _GEN7739 : _GEN7521;
wire  _GEN7741 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7742 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7743 = io_x[11] ? _GEN7742 : _GEN7741;
wire  _GEN7744 = io_x[9] ? _GEN7743 : _GEN7740;
wire  _GEN7745 = io_x[21] ? _GEN7744 : _GEN7738;
wire  _GEN7746 = io_x[31] ? _GEN7552 : _GEN7745;
wire  _GEN7747 = io_x[30] ? _GEN7746 : _GEN7734;
wire  _GEN7748 = io_x[29] ? _GEN7747 : _GEN7724;
wire  _GEN7749 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7750 = io_x[11] ? _GEN7749 : _GEN7521;
wire  _GEN7751 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7752 = io_x[11] ? _GEN7751 : _GEN7531;
wire  _GEN7753 = io_x[9] ? _GEN7752 : _GEN7750;
wire  _GEN7754 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7755 = io_x[11] ? _GEN7754 : _GEN7521;
wire  _GEN7756 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7757 = io_x[11] ? _GEN7756 : _GEN7521;
wire  _GEN7758 = io_x[9] ? _GEN7757 : _GEN7755;
wire  _GEN7759 = io_x[21] ? _GEN7758 : _GEN7753;
wire  _GEN7760 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7761 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7762 = io_x[11] ? _GEN7761 : _GEN7760;
wire  _GEN7763 = io_x[9] ? _GEN7762 : _GEN7530;
wire  _GEN7764 = io_x[21] ? _GEN7763 : _GEN7559;
wire  _GEN7765 = io_x[31] ? _GEN7764 : _GEN7759;
wire  _GEN7766 = io_x[30] ? _GEN7579 : _GEN7765;
wire  _GEN7767 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7768 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7769 = io_x[11] ? _GEN7768 : _GEN7767;
wire  _GEN7770 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7771 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7772 = io_x[11] ? _GEN7771 : _GEN7770;
wire  _GEN7773 = io_x[9] ? _GEN7772 : _GEN7769;
wire  _GEN7774 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7775 = io_x[11] ? _GEN7774 : _GEN7521;
wire  _GEN7776 = io_x[9] ? _GEN7548 : _GEN7775;
wire  _GEN7777 = io_x[21] ? _GEN7776 : _GEN7773;
wire  _GEN7778 = io_x[31] ? _GEN7552 : _GEN7777;
wire  _GEN7779 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7780 = io_x[11] ? _GEN7779 : _GEN7521;
wire  _GEN7781 = io_x[9] ? _GEN7780 : _GEN7548;
wire  _GEN7782 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7783 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7784 = io_x[11] ? _GEN7783 : _GEN7782;
wire  _GEN7785 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7786 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7787 = io_x[11] ? _GEN7786 : _GEN7785;
wire  _GEN7788 = io_x[9] ? _GEN7787 : _GEN7784;
wire  _GEN7789 = io_x[21] ? _GEN7788 : _GEN7781;
wire  _GEN7790 = io_x[31] ? _GEN7552 : _GEN7789;
wire  _GEN7791 = io_x[30] ? _GEN7790 : _GEN7778;
wire  _GEN7792 = io_x[29] ? _GEN7791 : _GEN7766;
wire  _GEN7793 = io_x[28] ? _GEN7792 : _GEN7748;
wire  _GEN7794 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7795 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7796 = io_x[11] ? _GEN7795 : _GEN7794;
wire  _GEN7797 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7798 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7799 = io_x[11] ? _GEN7798 : _GEN7797;
wire  _GEN7800 = io_x[9] ? _GEN7799 : _GEN7796;
wire  _GEN7801 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7802 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7803 = io_x[11] ? _GEN7802 : _GEN7801;
wire  _GEN7804 = io_x[9] ? _GEN7803 : _GEN7548;
wire  _GEN7805 = io_x[21] ? _GEN7804 : _GEN7800;
wire  _GEN7806 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7807 = io_x[11] ? _GEN7806 : _GEN7531;
wire  _GEN7808 = io_x[9] ? _GEN7807 : _GEN7530;
wire  _GEN7809 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7810 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7811 = io_x[11] ? _GEN7810 : _GEN7809;
wire  _GEN7812 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7813 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7814 = io_x[11] ? _GEN7813 : _GEN7812;
wire  _GEN7815 = io_x[9] ? _GEN7814 : _GEN7811;
wire  _GEN7816 = io_x[21] ? _GEN7815 : _GEN7808;
wire  _GEN7817 = io_x[31] ? _GEN7816 : _GEN7805;
wire  _GEN7818 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7819 = io_x[11] ? _GEN7818 : _GEN7521;
wire  _GEN7820 = io_x[9] ? _GEN7530 : _GEN7819;
wire  _GEN7821 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7822 = io_x[11] ? _GEN7821 : _GEN7521;
wire  _GEN7823 = io_x[9] ? _GEN7548 : _GEN7822;
wire  _GEN7824 = io_x[21] ? _GEN7823 : _GEN7820;
wire  _GEN7825 = io_x[31] ? _GEN7552 : _GEN7824;
wire  _GEN7826 = io_x[30] ? _GEN7825 : _GEN7817;
wire  _GEN7827 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7828 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7829 = io_x[11] ? _GEN7828 : _GEN7827;
wire  _GEN7830 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7831 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7832 = io_x[11] ? _GEN7831 : _GEN7830;
wire  _GEN7833 = io_x[9] ? _GEN7832 : _GEN7829;
wire  _GEN7834 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7835 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7836 = io_x[11] ? _GEN7835 : _GEN7834;
wire  _GEN7837 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7838 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7839 = io_x[11] ? _GEN7838 : _GEN7837;
wire  _GEN7840 = io_x[9] ? _GEN7839 : _GEN7836;
wire  _GEN7841 = io_x[21] ? _GEN7840 : _GEN7833;
wire  _GEN7842 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7843 = io_x[11] ? _GEN7842 : _GEN7531;
wire  _GEN7844 = io_x[9] ? _GEN7843 : _GEN7530;
wire  _GEN7845 = io_x[21] ? _GEN7559 : _GEN7844;
wire  _GEN7846 = io_x[31] ? _GEN7845 : _GEN7841;
wire  _GEN7847 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7848 = io_x[11] ? _GEN7531 : _GEN7847;
wire  _GEN7849 = io_x[9] ? _GEN7530 : _GEN7848;
wire  _GEN7850 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7851 = io_x[11] ? _GEN7850 : _GEN7521;
wire  _GEN7852 = io_x[9] ? _GEN7851 : _GEN7530;
wire  _GEN7853 = io_x[21] ? _GEN7852 : _GEN7849;
wire  _GEN7854 = io_x[31] ? _GEN7552 : _GEN7853;
wire  _GEN7855 = io_x[30] ? _GEN7854 : _GEN7846;
wire  _GEN7856 = io_x[29] ? _GEN7855 : _GEN7826;
wire  _GEN7857 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7858 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7859 = io_x[11] ? _GEN7858 : _GEN7857;
wire  _GEN7860 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7861 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7862 = io_x[11] ? _GEN7861 : _GEN7860;
wire  _GEN7863 = io_x[9] ? _GEN7862 : _GEN7859;
wire  _GEN7864 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7865 = io_x[11] ? _GEN7864 : _GEN7531;
wire  _GEN7866 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7867 = io_x[11] ? _GEN7866 : _GEN7531;
wire  _GEN7868 = io_x[9] ? _GEN7867 : _GEN7865;
wire  _GEN7869 = io_x[21] ? _GEN7868 : _GEN7863;
wire  _GEN7870 = io_x[11] ? _GEN7531 : _GEN7521;
wire  _GEN7871 = io_x[9] ? _GEN7870 : _GEN7548;
wire  _GEN7872 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7873 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7874 = io_x[11] ? _GEN7873 : _GEN7872;
wire  _GEN7875 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7876 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7877 = io_x[11] ? _GEN7876 : _GEN7875;
wire  _GEN7878 = io_x[9] ? _GEN7877 : _GEN7874;
wire  _GEN7879 = io_x[21] ? _GEN7878 : _GEN7871;
wire  _GEN7880 = io_x[31] ? _GEN7879 : _GEN7869;
wire  _GEN7881 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7882 = io_x[11] ? _GEN7881 : _GEN7521;
wire  _GEN7883 = io_x[9] ? _GEN7882 : _GEN7548;
wire  _GEN7884 = io_x[21] ? _GEN7883 : _GEN7520;
wire  _GEN7885 = io_x[31] ? _GEN7552 : _GEN7884;
wire  _GEN7886 = io_x[30] ? _GEN7885 : _GEN7880;
wire  _GEN7887 = io_x[11] ? _GEN7531 : _GEN7521;
wire  _GEN7888 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7889 = io_x[11] ? _GEN7888 : _GEN7531;
wire  _GEN7890 = io_x[9] ? _GEN7889 : _GEN7887;
wire  _GEN7891 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7892 = io_x[11] ? _GEN7891 : _GEN7521;
wire  _GEN7893 = io_x[9] ? _GEN7548 : _GEN7892;
wire  _GEN7894 = io_x[21] ? _GEN7893 : _GEN7890;
wire  _GEN7895 = io_x[31] ? _GEN7552 : _GEN7894;
wire  _GEN7896 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7897 = io_x[11] ? _GEN7896 : _GEN7521;
wire  _GEN7898 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7899 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7900 = io_x[11] ? _GEN7899 : _GEN7898;
wire  _GEN7901 = io_x[9] ? _GEN7900 : _GEN7897;
wire  _GEN7902 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7903 = io_x[11] ? _GEN7902 : _GEN7521;
wire  _GEN7904 = io_x[9] ? _GEN7548 : _GEN7903;
wire  _GEN7905 = io_x[21] ? _GEN7904 : _GEN7901;
wire  _GEN7906 = io_x[31] ? _GEN7552 : _GEN7905;
wire  _GEN7907 = io_x[30] ? _GEN7906 : _GEN7895;
wire  _GEN7908 = io_x[29] ? _GEN7907 : _GEN7886;
wire  _GEN7909 = io_x[28] ? _GEN7908 : _GEN7856;
wire  _GEN7910 = io_x[27] ? _GEN7909 : _GEN7793;
wire  _GEN7911 = io_x[16] ? _GEN7910 : _GEN7684;
wire  _GEN7912 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7913 = io_x[11] ? _GEN7912 : _GEN7531;
wire  _GEN7914 = io_x[9] ? _GEN7913 : _GEN7530;
wire  _GEN7915 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7916 = io_x[11] ? _GEN7915 : _GEN7531;
wire  _GEN7917 = io_x[9] ? _GEN7916 : _GEN7530;
wire  _GEN7918 = io_x[21] ? _GEN7917 : _GEN7914;
wire  _GEN7919 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7920 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7921 = io_x[11] ? _GEN7920 : _GEN7919;
wire  _GEN7922 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7923 = io_x[11] ? _GEN7922 : _GEN7521;
wire  _GEN7924 = io_x[9] ? _GEN7923 : _GEN7921;
wire  _GEN7925 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7926 = io_x[11] ? _GEN7925 : _GEN7531;
wire  _GEN7927 = io_x[9] ? _GEN7926 : _GEN7530;
wire  _GEN7928 = io_x[21] ? _GEN7927 : _GEN7924;
wire  _GEN7929 = io_x[31] ? _GEN7928 : _GEN7918;
wire  _GEN7930 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7931 = io_x[11] ? _GEN7521 : _GEN7930;
wire  _GEN7932 = io_x[9] ? _GEN7931 : _GEN7530;
wire  _GEN7933 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7934 = io_x[11] ? _GEN7933 : _GEN7521;
wire  _GEN7935 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7936 = io_x[11] ? _GEN7935 : _GEN7531;
wire  _GEN7937 = io_x[9] ? _GEN7936 : _GEN7934;
wire  _GEN7938 = io_x[21] ? _GEN7937 : _GEN7932;
wire  _GEN7939 = io_x[31] ? _GEN7552 : _GEN7938;
wire  _GEN7940 = io_x[30] ? _GEN7939 : _GEN7929;
wire  _GEN7941 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7942 = io_x[11] ? _GEN7941 : _GEN7521;
wire  _GEN7943 = io_x[9] ? _GEN7942 : _GEN7548;
wire  _GEN7944 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7945 = io_x[11] ? _GEN7944 : _GEN7521;
wire  _GEN7946 = io_x[9] ? _GEN7945 : _GEN7548;
wire  _GEN7947 = io_x[21] ? _GEN7946 : _GEN7943;
wire  _GEN7948 = io_x[31] ? _GEN7552 : _GEN7947;
wire  _GEN7949 = io_x[11] ? _GEN7531 : _GEN7521;
wire  _GEN7950 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7951 = io_x[11] ? _GEN7950 : _GEN7531;
wire  _GEN7952 = io_x[9] ? _GEN7951 : _GEN7949;
wire  _GEN7953 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7954 = io_x[11] ? _GEN7953 : _GEN7521;
wire  _GEN7955 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7956 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7957 = io_x[11] ? _GEN7956 : _GEN7955;
wire  _GEN7958 = io_x[9] ? _GEN7957 : _GEN7954;
wire  _GEN7959 = io_x[21] ? _GEN7958 : _GEN7952;
wire  _GEN7960 = io_x[31] ? _GEN7552 : _GEN7959;
wire  _GEN7961 = io_x[30] ? _GEN7960 : _GEN7948;
wire  _GEN7962 = io_x[29] ? _GEN7961 : _GEN7940;
wire  _GEN7963 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7964 = io_x[11] ? _GEN7963 : _GEN7521;
wire  _GEN7965 = io_x[9] ? _GEN7964 : _GEN7548;
wire  _GEN7966 = io_x[21] ? _GEN7965 : _GEN7520;
wire  _GEN7967 = io_x[31] ? _GEN7561 : _GEN7966;
wire  _GEN7968 = io_x[30] ? _GEN7579 : _GEN7967;
wire  _GEN7969 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7970 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7971 = io_x[11] ? _GEN7970 : _GEN7969;
wire  _GEN7972 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7973 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7974 = io_x[11] ? _GEN7973 : _GEN7972;
wire  _GEN7975 = io_x[9] ? _GEN7974 : _GEN7971;
wire  _GEN7976 = io_x[21] ? _GEN7520 : _GEN7975;
wire  _GEN7977 = io_x[31] ? _GEN7552 : _GEN7976;
wire  _GEN7978 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7979 = io_x[11] ? _GEN7521 : _GEN7978;
wire  _GEN7980 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7981 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7982 = io_x[11] ? _GEN7981 : _GEN7980;
wire  _GEN7983 = io_x[9] ? _GEN7982 : _GEN7979;
wire  _GEN7984 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7985 = io_x[11] ? _GEN7984 : _GEN7521;
wire  _GEN7986 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7987 = io_x[11] ? _GEN7521 : _GEN7986;
wire  _GEN7988 = io_x[9] ? _GEN7987 : _GEN7985;
wire  _GEN7989 = io_x[21] ? _GEN7988 : _GEN7983;
wire  _GEN7990 = io_x[31] ? _GEN7552 : _GEN7989;
wire  _GEN7991 = io_x[30] ? _GEN7990 : _GEN7977;
wire  _GEN7992 = io_x[29] ? _GEN7991 : _GEN7968;
wire  _GEN7993 = io_x[28] ? _GEN7992 : _GEN7962;
wire  _GEN7994 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7995 = io_x[11] ? _GEN7521 : _GEN7994;
wire  _GEN7996 = io_x[9] ? _GEN7995 : _GEN7548;
wire  _GEN7997 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN7998 = io_x[11] ? _GEN7997 : _GEN7531;
wire  _GEN7999 = io_x[9] ? _GEN7530 : _GEN7998;
wire  _GEN8000 = io_x[21] ? _GEN7999 : _GEN7996;
wire  _GEN8001 = io_x[21] ? _GEN7559 : _GEN7520;
wire  _GEN8002 = io_x[31] ? _GEN8001 : _GEN8000;
wire  _GEN8003 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8004 = io_x[11] ? _GEN8003 : _GEN7521;
wire  _GEN8005 = io_x[9] ? _GEN8004 : _GEN7548;
wire  _GEN8006 = io_x[21] ? _GEN8005 : _GEN7559;
wire  _GEN8007 = io_x[31] ? _GEN7552 : _GEN8006;
wire  _GEN8008 = io_x[30] ? _GEN8007 : _GEN8002;
wire  _GEN8009 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8010 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8011 = io_x[11] ? _GEN8010 : _GEN8009;
wire  _GEN8012 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8013 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8014 = io_x[11] ? _GEN8013 : _GEN8012;
wire  _GEN8015 = io_x[9] ? _GEN8014 : _GEN8011;
wire  _GEN8016 = io_x[21] ? _GEN7559 : _GEN8015;
wire  _GEN8017 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8018 = io_x[11] ? _GEN8017 : _GEN7531;
wire  _GEN8019 = io_x[9] ? _GEN7530 : _GEN8018;
wire  _GEN8020 = io_x[21] ? _GEN7520 : _GEN8019;
wire  _GEN8021 = io_x[31] ? _GEN8020 : _GEN8016;
wire  _GEN8022 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8023 = io_x[11] ? _GEN8022 : _GEN7531;
wire  _GEN8024 = io_x[9] ? _GEN7548 : _GEN8023;
wire  _GEN8025 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8026 = io_x[11] ? _GEN7531 : _GEN8025;
wire  _GEN8027 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8028 = io_x[11] ? _GEN7531 : _GEN8027;
wire  _GEN8029 = io_x[9] ? _GEN8028 : _GEN8026;
wire  _GEN8030 = io_x[21] ? _GEN8029 : _GEN8024;
wire  _GEN8031 = io_x[31] ? _GEN7552 : _GEN8030;
wire  _GEN8032 = io_x[30] ? _GEN8031 : _GEN8021;
wire  _GEN8033 = io_x[29] ? _GEN8032 : _GEN8008;
wire  _GEN8034 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8035 = io_x[11] ? _GEN8034 : _GEN7521;
wire  _GEN8036 = io_x[9] ? _GEN8035 : _GEN7530;
wire  _GEN8037 = io_x[21] ? _GEN7559 : _GEN8036;
wire  _GEN8038 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8039 = io_x[11] ? _GEN7521 : _GEN8038;
wire  _GEN8040 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8041 = io_x[11] ? _GEN8040 : _GEN7521;
wire  _GEN8042 = io_x[9] ? _GEN8041 : _GEN8039;
wire  _GEN8043 = io_x[11] ? _GEN7531 : _GEN7521;
wire  _GEN8044 = io_x[9] ? _GEN7548 : _GEN8043;
wire  _GEN8045 = io_x[21] ? _GEN8044 : _GEN8042;
wire  _GEN8046 = io_x[31] ? _GEN8045 : _GEN8037;
wire  _GEN8047 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8048 = io_x[11] ? _GEN8047 : _GEN7531;
wire  _GEN8049 = io_x[9] ? _GEN8048 : _GEN7530;
wire  _GEN8050 = io_x[21] ? _GEN7520 : _GEN8049;
wire  _GEN8051 = io_x[31] ? _GEN7552 : _GEN8050;
wire  _GEN8052 = io_x[30] ? _GEN8051 : _GEN8046;
wire  _GEN8053 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8054 = io_x[11] ? _GEN8053 : _GEN7521;
wire  _GEN8055 = io_x[9] ? _GEN8054 : _GEN7548;
wire  _GEN8056 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8057 = io_x[11] ? _GEN8056 : _GEN7521;
wire  _GEN8058 = io_x[9] ? _GEN8057 : _GEN7530;
wire  _GEN8059 = io_x[21] ? _GEN8058 : _GEN8055;
wire  _GEN8060 = io_x[31] ? _GEN7552 : _GEN8059;
wire  _GEN8061 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8062 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8063 = io_x[11] ? _GEN8062 : _GEN8061;
wire  _GEN8064 = io_x[9] ? _GEN8063 : _GEN7548;
wire  _GEN8065 = io_x[21] ? _GEN8064 : _GEN7559;
wire  _GEN8066 = io_x[31] ? _GEN7552 : _GEN8065;
wire  _GEN8067 = io_x[30] ? _GEN8066 : _GEN8060;
wire  _GEN8068 = io_x[29] ? _GEN8067 : _GEN8052;
wire  _GEN8069 = io_x[28] ? _GEN8068 : _GEN8033;
wire  _GEN8070 = io_x[27] ? _GEN8069 : _GEN7993;
wire  _GEN8071 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8072 = io_x[11] ? _GEN8071 : _GEN7531;
wire  _GEN8073 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8074 = io_x[11] ? _GEN8073 : _GEN7531;
wire  _GEN8075 = io_x[9] ? _GEN8074 : _GEN8072;
wire  _GEN8076 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8077 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8078 = io_x[11] ? _GEN8077 : _GEN8076;
wire  _GEN8079 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8080 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8081 = io_x[11] ? _GEN8080 : _GEN8079;
wire  _GEN8082 = io_x[9] ? _GEN8081 : _GEN8078;
wire  _GEN8083 = io_x[21] ? _GEN8082 : _GEN8075;
wire  _GEN8084 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8085 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8086 = io_x[11] ? _GEN8085 : _GEN8084;
wire  _GEN8087 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8088 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8089 = io_x[11] ? _GEN8088 : _GEN8087;
wire  _GEN8090 = io_x[9] ? _GEN8089 : _GEN8086;
wire  _GEN8091 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8092 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8093 = io_x[11] ? _GEN8092 : _GEN8091;
wire  _GEN8094 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8095 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8096 = io_x[11] ? _GEN8095 : _GEN8094;
wire  _GEN8097 = io_x[9] ? _GEN8096 : _GEN8093;
wire  _GEN8098 = io_x[21] ? _GEN8097 : _GEN8090;
wire  _GEN8099 = io_x[31] ? _GEN8098 : _GEN8083;
wire  _GEN8100 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8101 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8102 = io_x[11] ? _GEN8101 : _GEN8100;
wire  _GEN8103 = io_x[9] ? _GEN8102 : _GEN7530;
wire  _GEN8104 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8105 = io_x[11] ? _GEN8104 : _GEN7531;
wire  _GEN8106 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8107 = io_x[11] ? _GEN7521 : _GEN8106;
wire  _GEN8108 = io_x[9] ? _GEN8107 : _GEN8105;
wire  _GEN8109 = io_x[21] ? _GEN8108 : _GEN8103;
wire  _GEN8110 = io_x[31] ? _GEN7552 : _GEN8109;
wire  _GEN8111 = io_x[30] ? _GEN8110 : _GEN8099;
wire  _GEN8112 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8113 = io_x[11] ? _GEN8112 : _GEN7521;
wire  _GEN8114 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8115 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8116 = io_x[11] ? _GEN8115 : _GEN8114;
wire  _GEN8117 = io_x[9] ? _GEN8116 : _GEN8113;
wire  _GEN8118 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8119 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8120 = io_x[11] ? _GEN8119 : _GEN8118;
wire  _GEN8121 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8122 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8123 = io_x[11] ? _GEN8122 : _GEN8121;
wire  _GEN8124 = io_x[9] ? _GEN8123 : _GEN8120;
wire  _GEN8125 = io_x[21] ? _GEN8124 : _GEN8117;
wire  _GEN8126 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8127 = io_x[11] ? _GEN8126 : _GEN7521;
wire  _GEN8128 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8129 = io_x[11] ? _GEN7531 : _GEN8128;
wire  _GEN8130 = io_x[9] ? _GEN8129 : _GEN8127;
wire  _GEN8131 = io_x[21] ? _GEN7559 : _GEN8130;
wire  _GEN8132 = io_x[31] ? _GEN8131 : _GEN8125;
wire  _GEN8133 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8134 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8135 = io_x[11] ? _GEN8134 : _GEN8133;
wire  _GEN8136 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8137 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8138 = io_x[11] ? _GEN8137 : _GEN8136;
wire  _GEN8139 = io_x[9] ? _GEN8138 : _GEN8135;
wire  _GEN8140 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8141 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8142 = io_x[11] ? _GEN8141 : _GEN8140;
wire  _GEN8143 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8144 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8145 = io_x[11] ? _GEN8144 : _GEN8143;
wire  _GEN8146 = io_x[9] ? _GEN8145 : _GEN8142;
wire  _GEN8147 = io_x[21] ? _GEN8146 : _GEN8139;
wire  _GEN8148 = io_x[31] ? _GEN7552 : _GEN8147;
wire  _GEN8149 = io_x[30] ? _GEN8148 : _GEN8132;
wire  _GEN8150 = io_x[29] ? _GEN8149 : _GEN8111;
wire  _GEN8151 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8152 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8153 = io_x[11] ? _GEN8152 : _GEN8151;
wire  _GEN8154 = io_x[9] ? _GEN8153 : _GEN7530;
wire  _GEN8155 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8156 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8157 = io_x[11] ? _GEN8156 : _GEN8155;
wire  _GEN8158 = io_x[9] ? _GEN8157 : _GEN7530;
wire  _GEN8159 = io_x[21] ? _GEN8158 : _GEN8154;
wire  _GEN8160 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8161 = io_x[11] ? _GEN8160 : _GEN7531;
wire  _GEN8162 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8163 = io_x[11] ? _GEN8162 : _GEN7521;
wire  _GEN8164 = io_x[9] ? _GEN8163 : _GEN8161;
wire  _GEN8165 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8166 = io_x[11] ? _GEN7521 : _GEN8165;
wire  _GEN8167 = io_x[9] ? _GEN7548 : _GEN8166;
wire  _GEN8168 = io_x[21] ? _GEN8167 : _GEN8164;
wire  _GEN8169 = io_x[31] ? _GEN8168 : _GEN8159;
wire  _GEN8170 = io_x[21] ? _GEN7520 : _GEN7559;
wire  _GEN8171 = io_x[31] ? _GEN7552 : _GEN8170;
wire  _GEN8172 = io_x[30] ? _GEN8171 : _GEN8169;
wire  _GEN8173 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8174 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8175 = io_x[11] ? _GEN8174 : _GEN8173;
wire  _GEN8176 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8177 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8178 = io_x[11] ? _GEN8177 : _GEN8176;
wire  _GEN8179 = io_x[9] ? _GEN8178 : _GEN8175;
wire  _GEN8180 = io_x[21] ? _GEN7520 : _GEN8179;
wire  _GEN8181 = io_x[31] ? _GEN7552 : _GEN8180;
wire  _GEN8182 = io_x[11] ? _GEN7521 : _GEN7531;
wire  _GEN8183 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8184 = io_x[11] ? _GEN8183 : _GEN7521;
wire  _GEN8185 = io_x[9] ? _GEN8184 : _GEN8182;
wire  _GEN8186 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8187 = io_x[11] ? _GEN8186 : _GEN7521;
wire  _GEN8188 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8189 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8190 = io_x[11] ? _GEN8189 : _GEN8188;
wire  _GEN8191 = io_x[9] ? _GEN8190 : _GEN8187;
wire  _GEN8192 = io_x[21] ? _GEN8191 : _GEN8185;
wire  _GEN8193 = io_x[31] ? _GEN7552 : _GEN8192;
wire  _GEN8194 = io_x[30] ? _GEN8193 : _GEN8181;
wire  _GEN8195 = io_x[29] ? _GEN8194 : _GEN8172;
wire  _GEN8196 = io_x[28] ? _GEN8195 : _GEN8150;
wire  _GEN8197 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8198 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8199 = io_x[11] ? _GEN8198 : _GEN8197;
wire  _GEN8200 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8201 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8202 = io_x[11] ? _GEN8201 : _GEN8200;
wire  _GEN8203 = io_x[9] ? _GEN8202 : _GEN8199;
wire  _GEN8204 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8205 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8206 = io_x[11] ? _GEN8205 : _GEN8204;
wire  _GEN8207 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8208 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8209 = io_x[11] ? _GEN8208 : _GEN8207;
wire  _GEN8210 = io_x[9] ? _GEN8209 : _GEN8206;
wire  _GEN8211 = io_x[21] ? _GEN8210 : _GEN8203;
wire  _GEN8212 = io_x[11] ? _GEN7531 : _GEN7521;
wire  _GEN8213 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8214 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8215 = io_x[11] ? _GEN8214 : _GEN8213;
wire  _GEN8216 = io_x[9] ? _GEN8215 : _GEN8212;
wire  _GEN8217 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8218 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8219 = io_x[11] ? _GEN8218 : _GEN8217;
wire  _GEN8220 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8221 = io_x[11] ? _GEN8220 : _GEN7531;
wire  _GEN8222 = io_x[9] ? _GEN8221 : _GEN8219;
wire  _GEN8223 = io_x[21] ? _GEN8222 : _GEN8216;
wire  _GEN8224 = io_x[31] ? _GEN8223 : _GEN8211;
wire  _GEN8225 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8226 = io_x[11] ? _GEN8225 : _GEN7521;
wire  _GEN8227 = io_x[9] ? _GEN8226 : _GEN7548;
wire  _GEN8228 = io_x[21] ? _GEN8227 : _GEN7559;
wire  _GEN8229 = io_x[31] ? _GEN7552 : _GEN8228;
wire  _GEN8230 = io_x[30] ? _GEN8229 : _GEN8224;
wire  _GEN8231 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8232 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8233 = io_x[11] ? _GEN8232 : _GEN8231;
wire  _GEN8234 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8235 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8236 = io_x[11] ? _GEN8235 : _GEN8234;
wire  _GEN8237 = io_x[9] ? _GEN8236 : _GEN8233;
wire  _GEN8238 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8239 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8240 = io_x[11] ? _GEN8239 : _GEN8238;
wire  _GEN8241 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8242 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8243 = io_x[11] ? _GEN8242 : _GEN8241;
wire  _GEN8244 = io_x[9] ? _GEN8243 : _GEN8240;
wire  _GEN8245 = io_x[21] ? _GEN8244 : _GEN8237;
wire  _GEN8246 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8247 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8248 = io_x[11] ? _GEN8247 : _GEN8246;
wire  _GEN8249 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8250 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8251 = io_x[11] ? _GEN8250 : _GEN8249;
wire  _GEN8252 = io_x[9] ? _GEN8251 : _GEN8248;
wire  _GEN8253 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8254 = io_x[11] ? _GEN7531 : _GEN8253;
wire  _GEN8255 = io_x[9] ? _GEN8254 : _GEN7530;
wire  _GEN8256 = io_x[21] ? _GEN8255 : _GEN8252;
wire  _GEN8257 = io_x[31] ? _GEN8256 : _GEN8245;
wire  _GEN8258 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8259 = io_x[11] ? _GEN8258 : _GEN7521;
wire  _GEN8260 = io_x[9] ? _GEN8259 : _GEN7548;
wire  _GEN8261 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8262 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8263 = io_x[11] ? _GEN8262 : _GEN8261;
wire  _GEN8264 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8265 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8266 = io_x[11] ? _GEN8265 : _GEN8264;
wire  _GEN8267 = io_x[9] ? _GEN8266 : _GEN8263;
wire  _GEN8268 = io_x[21] ? _GEN8267 : _GEN8260;
wire  _GEN8269 = io_x[31] ? _GEN7552 : _GEN8268;
wire  _GEN8270 = io_x[30] ? _GEN8269 : _GEN8257;
wire  _GEN8271 = io_x[29] ? _GEN8270 : _GEN8230;
wire  _GEN8272 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8273 = io_x[11] ? _GEN8272 : _GEN7531;
wire  _GEN8274 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8275 = io_x[11] ? _GEN8274 : _GEN7521;
wire  _GEN8276 = io_x[9] ? _GEN8275 : _GEN8273;
wire  _GEN8277 = io_x[21] ? _GEN7520 : _GEN8276;
wire  _GEN8278 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8279 = io_x[11] ? _GEN8278 : _GEN7521;
wire  _GEN8280 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8281 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8282 = io_x[11] ? _GEN8281 : _GEN8280;
wire  _GEN8283 = io_x[9] ? _GEN8282 : _GEN8279;
wire  _GEN8284 = io_x[21] ? _GEN8283 : _GEN7559;
wire  _GEN8285 = io_x[31] ? _GEN8284 : _GEN8277;
wire  _GEN8286 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8287 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8288 = io_x[11] ? _GEN8287 : _GEN8286;
wire  _GEN8289 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8290 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8291 = io_x[11] ? _GEN8290 : _GEN8289;
wire  _GEN8292 = io_x[9] ? _GEN8291 : _GEN8288;
wire  _GEN8293 = io_x[21] ? _GEN7520 : _GEN8292;
wire  _GEN8294 = io_x[31] ? _GEN7552 : _GEN8293;
wire  _GEN8295 = io_x[30] ? _GEN8294 : _GEN8285;
wire  _GEN8296 = io_x[11] ? _GEN7531 : _GEN7521;
wire  _GEN8297 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8298 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8299 = io_x[11] ? _GEN8298 : _GEN8297;
wire  _GEN8300 = io_x[9] ? _GEN8299 : _GEN8296;
wire  _GEN8301 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8302 = io_x[11] ? _GEN8301 : _GEN7531;
wire  _GEN8303 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8304 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8305 = io_x[11] ? _GEN8304 : _GEN8303;
wire  _GEN8306 = io_x[9] ? _GEN8305 : _GEN8302;
wire  _GEN8307 = io_x[21] ? _GEN8306 : _GEN8300;
wire  _GEN8308 = io_x[31] ? _GEN7552 : _GEN8307;
wire  _GEN8309 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8310 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8311 = io_x[11] ? _GEN8310 : _GEN8309;
wire  _GEN8312 = io_x[9] ? _GEN8311 : _GEN7548;
wire  _GEN8313 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8314 = io_x[23] ? _GEN7523 : _GEN7522;
wire  _GEN8315 = io_x[11] ? _GEN8314 : _GEN8313;
wire  _GEN8316 = io_x[9] ? _GEN8315 : _GEN7548;
wire  _GEN8317 = io_x[21] ? _GEN8316 : _GEN8312;
wire  _GEN8318 = io_x[31] ? _GEN7552 : _GEN8317;
wire  _GEN8319 = io_x[30] ? _GEN8318 : _GEN8308;
wire  _GEN8320 = io_x[29] ? _GEN8319 : _GEN8295;
wire  _GEN8321 = io_x[28] ? _GEN8320 : _GEN8271;
wire  _GEN8322 = io_x[27] ? _GEN8321 : _GEN8196;
wire  _GEN8323 = io_x[16] ? _GEN8322 : _GEN8070;
wire  _GEN8324 = io_x[22] ? _GEN8323 : _GEN7911;
assign io_y[5] = _GEN8324;
wire  _GEN8325 = 1'b0;
wire  _GEN8326 = 1'b1;
wire  _GEN8327 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8328 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8329 = io_x[19] ? _GEN8328 : _GEN8327;
wire  _GEN8330 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8331 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8332 = io_x[19] ? _GEN8331 : _GEN8330;
wire  _GEN8333 = io_x[31] ? _GEN8332 : _GEN8329;
wire  _GEN8334 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8335 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8336 = io_x[19] ? _GEN8335 : _GEN8334;
wire  _GEN8337 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8338 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8339 = io_x[19] ? _GEN8338 : _GEN8337;
wire  _GEN8340 = io_x[31] ? _GEN8339 : _GEN8336;
wire  _GEN8341 = io_x[1] ? _GEN8340 : _GEN8333;
wire  _GEN8342 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8343 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8344 = io_x[19] ? _GEN8343 : _GEN8342;
wire  _GEN8345 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8346 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8347 = io_x[19] ? _GEN8346 : _GEN8345;
wire  _GEN8348 = io_x[31] ? _GEN8347 : _GEN8344;
wire  _GEN8349 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8350 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8351 = io_x[19] ? _GEN8350 : _GEN8349;
wire  _GEN8352 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8353 = io_x[22] ? _GEN8326 : _GEN8325;
wire  _GEN8354 = io_x[19] ? _GEN8353 : _GEN8352;
wire  _GEN8355 = io_x[31] ? _GEN8354 : _GEN8351;
wire  _GEN8356 = io_x[1] ? _GEN8355 : _GEN8348;
wire  _GEN8357 = io_x[3] ? _GEN8356 : _GEN8341;
assign io_y[4] = _GEN8357;
wire  _GEN8358 = 1'b0;
wire  _GEN8359 = 1'b1;
wire  _GEN8360 = io_x[21] ? _GEN8359 : _GEN8358;
assign io_y[3] = _GEN8360;
wire  _GEN8361 = 1'b0;
wire  _GEN8362 = 1'b1;
wire  _GEN8363 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8364 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8365 = io_x[21] ? _GEN8364 : _GEN8363;
wire  _GEN8366 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8367 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8368 = io_x[21] ? _GEN8367 : _GEN8366;
wire  _GEN8369 = io_x[5] ? _GEN8368 : _GEN8365;
wire  _GEN8370 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8371 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8372 = io_x[21] ? _GEN8371 : _GEN8370;
wire  _GEN8373 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8374 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8375 = io_x[21] ? _GEN8374 : _GEN8373;
wire  _GEN8376 = io_x[5] ? _GEN8375 : _GEN8372;
wire  _GEN8377 = io_x[3] ? _GEN8376 : _GEN8369;
wire  _GEN8378 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8379 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8380 = io_x[21] ? _GEN8379 : _GEN8378;
wire  _GEN8381 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8382 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8383 = io_x[21] ? _GEN8382 : _GEN8381;
wire  _GEN8384 = io_x[5] ? _GEN8383 : _GEN8380;
wire  _GEN8385 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8386 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8387 = io_x[21] ? _GEN8386 : _GEN8385;
wire  _GEN8388 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8389 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8390 = io_x[21] ? _GEN8389 : _GEN8388;
wire  _GEN8391 = io_x[5] ? _GEN8390 : _GEN8387;
wire  _GEN8392 = io_x[3] ? _GEN8391 : _GEN8384;
wire  _GEN8393 = io_x[29] ? _GEN8392 : _GEN8377;
wire  _GEN8394 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8395 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8396 = io_x[21] ? _GEN8395 : _GEN8394;
wire  _GEN8397 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8398 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8399 = io_x[21] ? _GEN8398 : _GEN8397;
wire  _GEN8400 = io_x[5] ? _GEN8399 : _GEN8396;
wire  _GEN8401 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8402 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8403 = io_x[21] ? _GEN8402 : _GEN8401;
wire  _GEN8404 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8405 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8406 = io_x[21] ? _GEN8405 : _GEN8404;
wire  _GEN8407 = io_x[5] ? _GEN8406 : _GEN8403;
wire  _GEN8408 = io_x[3] ? _GEN8407 : _GEN8400;
wire  _GEN8409 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8410 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8411 = io_x[21] ? _GEN8410 : _GEN8409;
wire  _GEN8412 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8413 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8414 = io_x[21] ? _GEN8413 : _GEN8412;
wire  _GEN8415 = io_x[5] ? _GEN8414 : _GEN8411;
wire  _GEN8416 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8417 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8418 = io_x[21] ? _GEN8417 : _GEN8416;
wire  _GEN8419 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8420 = io_x[20] ? _GEN8362 : _GEN8361;
wire  _GEN8421 = io_x[21] ? _GEN8420 : _GEN8419;
wire  _GEN8422 = io_x[5] ? _GEN8421 : _GEN8418;
wire  _GEN8423 = io_x[3] ? _GEN8422 : _GEN8415;
wire  _GEN8424 = io_x[29] ? _GEN8423 : _GEN8408;
wire  _GEN8425 = io_x[16] ? _GEN8424 : _GEN8393;
assign io_y[2] = _GEN8425;
wire  _GEN8426 = 1'b0;
wire  _GEN8427 = 1'b1;
wire  _GEN8428 = io_x[19] ? _GEN8427 : _GEN8426;
wire  _GEN8429 = io_x[19] ? _GEN8427 : _GEN8426;
wire  _GEN8430 = io_x[1] ? _GEN8429 : _GEN8428;
wire  _GEN8431 = io_x[19] ? _GEN8427 : _GEN8426;
wire  _GEN8432 = io_x[19] ? _GEN8427 : _GEN8426;
wire  _GEN8433 = io_x[1] ? _GEN8432 : _GEN8431;
wire  _GEN8434 = io_x[21] ? _GEN8433 : _GEN8430;
wire  _GEN8435 = io_x[19] ? _GEN8427 : _GEN8426;
wire  _GEN8436 = io_x[19] ? _GEN8427 : _GEN8426;
wire  _GEN8437 = io_x[1] ? _GEN8436 : _GEN8435;
wire  _GEN8438 = io_x[19] ? _GEN8427 : _GEN8426;
wire  _GEN8439 = io_x[19] ? _GEN8427 : _GEN8426;
wire  _GEN8440 = io_x[1] ? _GEN8439 : _GEN8438;
wire  _GEN8441 = io_x[21] ? _GEN8440 : _GEN8437;
wire  _GEN8442 = io_x[29] ? _GEN8441 : _GEN8434;
assign io_y[1] = _GEN8442;
wire  _GEN8443 = 1'b0;
wire  _GEN8444 = 1'b1;
wire  _GEN8445 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8446 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8447 = io_x[6] ? _GEN8446 : _GEN8445;
wire  _GEN8448 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8449 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8450 = io_x[6] ? _GEN8449 : _GEN8448;
wire  _GEN8451 = io_x[2] ? _GEN8450 : _GEN8447;
wire  _GEN8452 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8453 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8454 = io_x[6] ? _GEN8453 : _GEN8452;
wire  _GEN8455 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8456 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8457 = io_x[6] ? _GEN8456 : _GEN8455;
wire  _GEN8458 = io_x[2] ? _GEN8457 : _GEN8454;
wire  _GEN8459 = io_x[30] ? _GEN8458 : _GEN8451;
wire  _GEN8460 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8461 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8462 = io_x[6] ? _GEN8461 : _GEN8460;
wire  _GEN8463 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8464 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8465 = io_x[6] ? _GEN8464 : _GEN8463;
wire  _GEN8466 = io_x[2] ? _GEN8465 : _GEN8462;
wire  _GEN8467 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8468 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8469 = io_x[6] ? _GEN8468 : _GEN8467;
wire  _GEN8470 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8471 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8472 = io_x[6] ? _GEN8471 : _GEN8470;
wire  _GEN8473 = io_x[2] ? _GEN8472 : _GEN8469;
wire  _GEN8474 = io_x[30] ? _GEN8473 : _GEN8466;
wire  _GEN8475 = io_x[4] ? _GEN8474 : _GEN8459;
wire  _GEN8476 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8477 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8478 = io_x[6] ? _GEN8477 : _GEN8476;
wire  _GEN8479 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8480 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8481 = io_x[6] ? _GEN8480 : _GEN8479;
wire  _GEN8482 = io_x[2] ? _GEN8481 : _GEN8478;
wire  _GEN8483 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8484 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8485 = io_x[6] ? _GEN8484 : _GEN8483;
wire  _GEN8486 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8487 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8488 = io_x[6] ? _GEN8487 : _GEN8486;
wire  _GEN8489 = io_x[2] ? _GEN8488 : _GEN8485;
wire  _GEN8490 = io_x[30] ? _GEN8489 : _GEN8482;
wire  _GEN8491 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8492 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8493 = io_x[6] ? _GEN8492 : _GEN8491;
wire  _GEN8494 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8495 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8496 = io_x[6] ? _GEN8495 : _GEN8494;
wire  _GEN8497 = io_x[2] ? _GEN8496 : _GEN8493;
wire  _GEN8498 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8499 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8500 = io_x[6] ? _GEN8499 : _GEN8498;
wire  _GEN8501 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8502 = io_x[16] ? _GEN8444 : _GEN8443;
wire  _GEN8503 = io_x[6] ? _GEN8502 : _GEN8501;
wire  _GEN8504 = io_x[2] ? _GEN8503 : _GEN8500;
wire  _GEN8505 = io_x[30] ? _GEN8504 : _GEN8497;
wire  _GEN8506 = io_x[4] ? _GEN8505 : _GEN8490;
wire  _GEN8507 = io_x[0] ? _GEN8506 : _GEN8475;
assign io_y[0] = _GEN8507;
endmodule