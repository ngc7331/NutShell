module BBGSharePredictorImp_BSD_sim(
    input [31:0] pc,
    input [31:0] train_pc,
    input  train_taken,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    input [15:0] train_ghr_rdata,
    output  taken,
    output  pht_wdata,
    output [8:0] pht_raddr,
    output [8:0] pht_waddr,
    output  ghr_wdata
);
wire [98:0] io_x;
wire [20:0] io_y;
assign io_x = { pc, train_pc, train_taken, pht_rdata, ghr_rdata, train_ghr_rdata };
assign { taken, pht_wdata, pht_raddr, pht_waddr, ghr_wdata } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN3 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN4 = io_x[22] ? _GEN3 : _GEN2;
wire  _GEN5 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN6 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN7 = io_x[22] ? _GEN6 : _GEN5;
wire  _GEN8 = io_x[28] ? _GEN7 : _GEN4;
wire  _GEN9 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN10 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN11 = io_x[22] ? _GEN10 : _GEN9;
wire  _GEN12 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN13 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN14 = io_x[22] ? _GEN13 : _GEN12;
wire  _GEN15 = io_x[28] ? _GEN14 : _GEN11;
wire  _GEN16 = io_x[81] ? _GEN15 : _GEN8;
wire  _GEN17 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN18 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN19 = io_x[22] ? _GEN18 : _GEN17;
wire  _GEN20 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN21 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN22 = io_x[22] ? _GEN21 : _GEN20;
wire  _GEN23 = io_x[28] ? _GEN22 : _GEN19;
wire  _GEN24 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN25 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN26 = io_x[22] ? _GEN25 : _GEN24;
wire  _GEN27 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN28 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN29 = io_x[22] ? _GEN28 : _GEN27;
wire  _GEN30 = io_x[28] ? _GEN29 : _GEN26;
wire  _GEN31 = io_x[81] ? _GEN30 : _GEN23;
wire  _GEN32 = io_x[18] ? _GEN31 : _GEN16;
wire  _GEN33 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN34 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN35 = io_x[22] ? _GEN34 : _GEN33;
wire  _GEN36 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN37 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN38 = io_x[22] ? _GEN37 : _GEN36;
wire  _GEN39 = io_x[28] ? _GEN38 : _GEN35;
wire  _GEN40 = 1'b1;
wire  _GEN41 = io_x[81] ? _GEN40 : _GEN39;
wire  _GEN42 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN43 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN44 = io_x[22] ? _GEN43 : _GEN42;
wire  _GEN45 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN46 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN47 = io_x[22] ? _GEN46 : _GEN45;
wire  _GEN48 = io_x[28] ? _GEN47 : _GEN44;
wire  _GEN49 = io_x[81] ? _GEN40 : _GEN48;
wire  _GEN50 = io_x[18] ? _GEN49 : _GEN41;
wire  _GEN51 = io_x[80] ? _GEN50 : _GEN32;
wire  _GEN52 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN53 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN54 = io_x[22] ? _GEN53 : _GEN52;
wire  _GEN55 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN56 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN57 = io_x[22] ? _GEN56 : _GEN55;
wire  _GEN58 = io_x[28] ? _GEN57 : _GEN54;
wire  _GEN59 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN60 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN61 = io_x[22] ? _GEN60 : _GEN59;
wire  _GEN62 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN63 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN64 = io_x[22] ? _GEN63 : _GEN62;
wire  _GEN65 = io_x[28] ? _GEN64 : _GEN61;
wire  _GEN66 = io_x[81] ? _GEN65 : _GEN58;
wire  _GEN67 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN68 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN69 = io_x[22] ? _GEN68 : _GEN67;
wire  _GEN70 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN71 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN72 = io_x[22] ? _GEN71 : _GEN70;
wire  _GEN73 = io_x[28] ? _GEN72 : _GEN69;
wire  _GEN74 = 1'b0;
wire  _GEN75 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN76 = io_x[22] ? _GEN75 : _GEN74;
wire  _GEN77 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN78 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN79 = io_x[22] ? _GEN78 : _GEN77;
wire  _GEN80 = io_x[28] ? _GEN79 : _GEN76;
wire  _GEN81 = io_x[81] ? _GEN80 : _GEN73;
wire  _GEN82 = io_x[18] ? _GEN81 : _GEN66;
wire  _GEN83 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN84 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN85 = io_x[22] ? _GEN84 : _GEN83;
wire  _GEN86 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN87 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN88 = io_x[22] ? _GEN87 : _GEN86;
wire  _GEN89 = io_x[28] ? _GEN88 : _GEN85;
wire  _GEN90 = io_x[81] ? _GEN40 : _GEN89;
wire  _GEN91 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN92 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN93 = io_x[22] ? _GEN92 : _GEN91;
wire  _GEN94 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN95 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN96 = io_x[22] ? _GEN95 : _GEN94;
wire  _GEN97 = io_x[28] ? _GEN96 : _GEN93;
wire  _GEN98 = io_x[81] ? _GEN40 : _GEN97;
wire  _GEN99 = io_x[18] ? _GEN98 : _GEN90;
wire  _GEN100 = io_x[80] ? _GEN99 : _GEN82;
wire  _GEN101 = io_x[20] ? _GEN100 : _GEN51;
wire  _GEN102 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN103 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN104 = io_x[22] ? _GEN103 : _GEN102;
wire  _GEN105 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN106 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN107 = io_x[22] ? _GEN106 : _GEN105;
wire  _GEN108 = io_x[28] ? _GEN107 : _GEN104;
wire  _GEN109 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN110 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN111 = io_x[22] ? _GEN110 : _GEN109;
wire  _GEN112 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN113 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN114 = io_x[22] ? _GEN113 : _GEN112;
wire  _GEN115 = io_x[28] ? _GEN114 : _GEN111;
wire  _GEN116 = io_x[81] ? _GEN115 : _GEN108;
wire  _GEN117 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN118 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN119 = io_x[22] ? _GEN118 : _GEN117;
wire  _GEN120 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN121 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN122 = io_x[22] ? _GEN121 : _GEN120;
wire  _GEN123 = io_x[28] ? _GEN122 : _GEN119;
wire  _GEN124 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN125 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN126 = io_x[22] ? _GEN125 : _GEN124;
wire  _GEN127 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN128 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN129 = io_x[22] ? _GEN128 : _GEN127;
wire  _GEN130 = io_x[28] ? _GEN129 : _GEN126;
wire  _GEN131 = io_x[81] ? _GEN130 : _GEN123;
wire  _GEN132 = io_x[18] ? _GEN131 : _GEN116;
wire  _GEN133 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN134 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN135 = io_x[22] ? _GEN134 : _GEN133;
wire  _GEN136 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN137 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN138 = io_x[22] ? _GEN137 : _GEN136;
wire  _GEN139 = io_x[28] ? _GEN138 : _GEN135;
wire  _GEN140 = io_x[81] ? _GEN40 : _GEN139;
wire  _GEN141 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN142 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN143 = io_x[22] ? _GEN142 : _GEN141;
wire  _GEN144 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN145 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN146 = io_x[22] ? _GEN145 : _GEN144;
wire  _GEN147 = io_x[28] ? _GEN146 : _GEN143;
wire  _GEN148 = io_x[81] ? _GEN40 : _GEN147;
wire  _GEN149 = io_x[18] ? _GEN148 : _GEN140;
wire  _GEN150 = io_x[80] ? _GEN149 : _GEN132;
wire  _GEN151 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN152 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN153 = io_x[22] ? _GEN152 : _GEN151;
wire  _GEN154 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN155 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN156 = io_x[22] ? _GEN155 : _GEN154;
wire  _GEN157 = io_x[28] ? _GEN156 : _GEN153;
wire  _GEN158 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN159 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN160 = io_x[22] ? _GEN159 : _GEN158;
wire  _GEN161 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN162 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN163 = io_x[22] ? _GEN162 : _GEN161;
wire  _GEN164 = io_x[28] ? _GEN163 : _GEN160;
wire  _GEN165 = io_x[81] ? _GEN164 : _GEN157;
wire  _GEN166 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN167 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN168 = io_x[22] ? _GEN167 : _GEN166;
wire  _GEN169 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN170 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN171 = io_x[22] ? _GEN170 : _GEN169;
wire  _GEN172 = io_x[28] ? _GEN171 : _GEN168;
wire  _GEN173 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN174 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN175 = io_x[22] ? _GEN174 : _GEN173;
wire  _GEN176 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN177 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN178 = io_x[22] ? _GEN177 : _GEN176;
wire  _GEN179 = io_x[28] ? _GEN178 : _GEN175;
wire  _GEN180 = io_x[81] ? _GEN179 : _GEN172;
wire  _GEN181 = io_x[18] ? _GEN180 : _GEN165;
wire  _GEN182 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN183 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN184 = io_x[22] ? _GEN183 : _GEN182;
wire  _GEN185 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN186 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN187 = io_x[22] ? _GEN186 : _GEN185;
wire  _GEN188 = io_x[28] ? _GEN187 : _GEN184;
wire  _GEN189 = io_x[81] ? _GEN40 : _GEN188;
wire  _GEN190 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN191 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN192 = io_x[22] ? _GEN191 : _GEN190;
wire  _GEN193 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN194 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN195 = io_x[22] ? _GEN194 : _GEN193;
wire  _GEN196 = io_x[28] ? _GEN195 : _GEN192;
wire  _GEN197 = io_x[81] ? _GEN40 : _GEN196;
wire  _GEN198 = io_x[18] ? _GEN197 : _GEN189;
wire  _GEN199 = io_x[80] ? _GEN198 : _GEN181;
wire  _GEN200 = io_x[20] ? _GEN199 : _GEN150;
wire  _GEN201 = io_x[16] ? _GEN200 : _GEN101;
assign io_y[20] = _GEN201;
wire  _GEN202 = 1'b0;
wire  _GEN203 = 1'b1;
wire  _GEN204 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN205 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN206 = io_x[33] ? _GEN205 : _GEN204;
wire  _GEN207 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN208 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN209 = io_x[33] ? _GEN208 : _GEN207;
wire  _GEN210 = io_x[22] ? _GEN209 : _GEN206;
wire  _GEN211 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN212 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN213 = io_x[33] ? _GEN212 : _GEN211;
wire  _GEN214 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN215 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN216 = io_x[33] ? _GEN215 : _GEN214;
wire  _GEN217 = io_x[22] ? _GEN216 : _GEN213;
wire  _GEN218 = io_x[18] ? _GEN217 : _GEN210;
wire  _GEN219 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN220 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN221 = io_x[33] ? _GEN220 : _GEN219;
wire  _GEN222 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN223 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN224 = io_x[33] ? _GEN223 : _GEN222;
wire  _GEN225 = io_x[22] ? _GEN224 : _GEN221;
wire  _GEN226 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN227 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN228 = io_x[33] ? _GEN227 : _GEN226;
wire  _GEN229 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN230 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN231 = io_x[33] ? _GEN230 : _GEN229;
wire  _GEN232 = io_x[22] ? _GEN231 : _GEN228;
wire  _GEN233 = io_x[18] ? _GEN232 : _GEN225;
wire  _GEN234 = io_x[80] ? _GEN233 : _GEN218;
wire  _GEN235 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN236 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN237 = io_x[33] ? _GEN236 : _GEN235;
wire  _GEN238 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN239 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN240 = io_x[33] ? _GEN239 : _GEN238;
wire  _GEN241 = io_x[22] ? _GEN240 : _GEN237;
wire  _GEN242 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN243 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN244 = io_x[33] ? _GEN243 : _GEN242;
wire  _GEN245 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN246 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN247 = io_x[33] ? _GEN246 : _GEN245;
wire  _GEN248 = io_x[22] ? _GEN247 : _GEN244;
wire  _GEN249 = io_x[18] ? _GEN248 : _GEN241;
wire  _GEN250 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN251 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN252 = io_x[33] ? _GEN251 : _GEN250;
wire  _GEN253 = 1'b1;
wire  _GEN254 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN255 = io_x[33] ? _GEN254 : _GEN253;
wire  _GEN256 = io_x[22] ? _GEN255 : _GEN252;
wire  _GEN257 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN258 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN259 = io_x[33] ? _GEN258 : _GEN257;
wire  _GEN260 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN261 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN262 = io_x[33] ? _GEN261 : _GEN260;
wire  _GEN263 = io_x[22] ? _GEN262 : _GEN259;
wire  _GEN264 = io_x[18] ? _GEN263 : _GEN256;
wire  _GEN265 = io_x[80] ? _GEN264 : _GEN249;
wire  _GEN266 = io_x[20] ? _GEN265 : _GEN234;
wire  _GEN267 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN268 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN269 = io_x[33] ? _GEN268 : _GEN267;
wire  _GEN270 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN271 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN272 = io_x[33] ? _GEN271 : _GEN270;
wire  _GEN273 = io_x[22] ? _GEN272 : _GEN269;
wire  _GEN274 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN275 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN276 = io_x[33] ? _GEN275 : _GEN274;
wire  _GEN277 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN278 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN279 = io_x[33] ? _GEN278 : _GEN277;
wire  _GEN280 = io_x[22] ? _GEN279 : _GEN276;
wire  _GEN281 = io_x[18] ? _GEN280 : _GEN273;
wire  _GEN282 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN283 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN284 = io_x[33] ? _GEN283 : _GEN282;
wire  _GEN285 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN286 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN287 = io_x[33] ? _GEN286 : _GEN285;
wire  _GEN288 = io_x[22] ? _GEN287 : _GEN284;
wire  _GEN289 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN290 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN291 = io_x[33] ? _GEN290 : _GEN289;
wire  _GEN292 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN293 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN294 = io_x[33] ? _GEN293 : _GEN292;
wire  _GEN295 = io_x[22] ? _GEN294 : _GEN291;
wire  _GEN296 = io_x[18] ? _GEN295 : _GEN288;
wire  _GEN297 = io_x[80] ? _GEN296 : _GEN281;
wire  _GEN298 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN299 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN300 = io_x[33] ? _GEN299 : _GEN298;
wire  _GEN301 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN302 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN303 = io_x[33] ? _GEN302 : _GEN301;
wire  _GEN304 = io_x[22] ? _GEN303 : _GEN300;
wire  _GEN305 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN306 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN307 = io_x[33] ? _GEN306 : _GEN305;
wire  _GEN308 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN309 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN310 = io_x[33] ? _GEN309 : _GEN308;
wire  _GEN311 = io_x[22] ? _GEN310 : _GEN307;
wire  _GEN312 = io_x[18] ? _GEN311 : _GEN304;
wire  _GEN313 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN314 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN315 = io_x[33] ? _GEN314 : _GEN313;
wire  _GEN316 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN317 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN318 = io_x[33] ? _GEN317 : _GEN316;
wire  _GEN319 = io_x[22] ? _GEN318 : _GEN315;
wire  _GEN320 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN321 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN322 = io_x[33] ? _GEN321 : _GEN320;
wire  _GEN323 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN324 = io_x[34] ? _GEN203 : _GEN202;
wire  _GEN325 = io_x[33] ? _GEN324 : _GEN323;
wire  _GEN326 = io_x[22] ? _GEN325 : _GEN322;
wire  _GEN327 = io_x[18] ? _GEN326 : _GEN319;
wire  _GEN328 = io_x[80] ? _GEN327 : _GEN312;
wire  _GEN329 = io_x[20] ? _GEN328 : _GEN297;
wire  _GEN330 = io_x[16] ? _GEN329 : _GEN266;
assign io_y[19] = _GEN330;
wire  _GEN331 = 1'b0;
wire  _GEN332 = 1'b1;
wire  _GEN333 = 1'b1;
wire  _GEN334 = 1'b0;
wire  _GEN335 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN336 = 1'b0;
wire  _GEN337 = io_x[27] ? _GEN336 : _GEN335;
wire  _GEN338 = 1'b0;
wire  _GEN339 = io_x[19] ? _GEN338 : _GEN337;
wire  _GEN340 = io_x[23] ? _GEN339 : _GEN332;
wire  _GEN341 = io_x[18] ? _GEN340 : _GEN331;
wire  _GEN342 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN343 = 1'b1;
wire  _GEN344 = io_x[27] ? _GEN343 : _GEN342;
wire  _GEN345 = 1'b1;
wire  _GEN346 = io_x[19] ? _GEN345 : _GEN344;
wire  _GEN347 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN348 = io_x[27] ? _GEN347 : _GEN336;
wire  _GEN349 = io_x[19] ? _GEN348 : _GEN345;
wire  _GEN350 = io_x[23] ? _GEN349 : _GEN346;
wire  _GEN351 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN352 = io_x[27] ? _GEN351 : _GEN343;
wire  _GEN353 = io_x[19] ? _GEN352 : _GEN345;
wire  _GEN354 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN355 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN356 = io_x[27] ? _GEN355 : _GEN354;
wire  _GEN357 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN358 = io_x[19] ? _GEN357 : _GEN356;
wire  _GEN359 = io_x[23] ? _GEN358 : _GEN353;
wire  _GEN360 = io_x[18] ? _GEN359 : _GEN350;
wire  _GEN361 = io_x[33] ? _GEN360 : _GEN341;
wire  _GEN362 = 1'b1;
wire  _GEN363 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN364 = io_x[27] ? _GEN363 : _GEN343;
wire  _GEN365 = io_x[19] ? _GEN345 : _GEN364;
wire  _GEN366 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN367 = io_x[19] ? _GEN345 : _GEN366;
wire  _GEN368 = io_x[23] ? _GEN367 : _GEN365;
wire  _GEN369 = io_x[18] ? _GEN368 : _GEN362;
wire  _GEN370 = 1'b0;
wire  _GEN371 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN372 = io_x[27] ? _GEN371 : _GEN343;
wire  _GEN373 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN374 = io_x[27] ? _GEN373 : _GEN343;
wire  _GEN375 = io_x[19] ? _GEN374 : _GEN372;
wire  _GEN376 = io_x[23] ? _GEN375 : _GEN370;
wire  _GEN377 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN378 = io_x[27] ? _GEN377 : _GEN336;
wire  _GEN379 = io_x[19] ? _GEN345 : _GEN378;
wire  _GEN380 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN381 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN382 = io_x[27] ? _GEN381 : _GEN380;
wire  _GEN383 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN384 = io_x[27] ? _GEN383 : _GEN336;
wire  _GEN385 = io_x[19] ? _GEN384 : _GEN382;
wire  _GEN386 = io_x[23] ? _GEN385 : _GEN379;
wire  _GEN387 = io_x[18] ? _GEN386 : _GEN376;
wire  _GEN388 = io_x[33] ? _GEN387 : _GEN369;
wire  _GEN389 = io_x[31] ? _GEN388 : _GEN361;
wire  _GEN390 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN391 = io_x[27] ? _GEN390 : _GEN343;
wire  _GEN392 = io_x[19] ? _GEN338 : _GEN391;
wire  _GEN393 = io_x[23] ? _GEN392 : _GEN370;
wire  _GEN394 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN395 = io_x[19] ? _GEN338 : _GEN394;
wire  _GEN396 = io_x[23] ? _GEN395 : _GEN332;
wire  _GEN397 = io_x[18] ? _GEN396 : _GEN393;
wire  _GEN398 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN399 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN400 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN401 = io_x[27] ? _GEN400 : _GEN343;
wire  _GEN402 = io_x[19] ? _GEN401 : _GEN399;
wire  _GEN403 = io_x[23] ? _GEN402 : _GEN370;
wire  _GEN404 = io_x[18] ? _GEN403 : _GEN398;
wire  _GEN405 = io_x[33] ? _GEN404 : _GEN397;
wire  _GEN406 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN407 = io_x[27] ? _GEN343 : _GEN406;
wire  _GEN408 = io_x[19] ? _GEN407 : _GEN345;
wire  _GEN409 = io_x[23] ? _GEN408 : _GEN332;
wire  _GEN410 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN411 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN412 = io_x[19] ? _GEN411 : _GEN345;
wire  _GEN413 = io_x[23] ? _GEN412 : _GEN410;
wire  _GEN414 = io_x[18] ? _GEN413 : _GEN409;
wire  _GEN415 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN416 = io_x[19] ? _GEN415 : _GEN345;
wire  _GEN417 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN418 = io_x[27] ? _GEN343 : _GEN417;
wire  _GEN419 = io_x[19] ? _GEN418 : _GEN345;
wire  _GEN420 = io_x[23] ? _GEN419 : _GEN416;
wire  _GEN421 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN422 = io_x[19] ? _GEN345 : _GEN421;
wire  _GEN423 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN424 = io_x[27] ? _GEN423 : _GEN343;
wire  _GEN425 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN426 = io_x[27] ? _GEN425 : _GEN336;
wire  _GEN427 = io_x[19] ? _GEN426 : _GEN424;
wire  _GEN428 = io_x[23] ? _GEN427 : _GEN422;
wire  _GEN429 = io_x[18] ? _GEN428 : _GEN420;
wire  _GEN430 = io_x[33] ? _GEN429 : _GEN414;
wire  _GEN431 = io_x[31] ? _GEN430 : _GEN405;
wire  _GEN432 = io_x[28] ? _GEN431 : _GEN389;
wire  _GEN433 = io_x[23] ? _GEN332 : _GEN370;
wire  _GEN434 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN435 = io_x[19] ? _GEN434 : _GEN338;
wire  _GEN436 = io_x[23] ? _GEN435 : _GEN332;
wire  _GEN437 = io_x[18] ? _GEN436 : _GEN433;
wire  _GEN438 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN439 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN440 = io_x[19] ? _GEN439 : _GEN345;
wire  _GEN441 = io_x[23] ? _GEN440 : _GEN438;
wire  _GEN442 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN443 = io_x[27] ? _GEN442 : _GEN343;
wire  _GEN444 = io_x[19] ? _GEN443 : _GEN345;
wire  _GEN445 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN446 = io_x[27] ? _GEN445 : _GEN343;
wire  _GEN447 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN448 = io_x[19] ? _GEN447 : _GEN446;
wire  _GEN449 = io_x[23] ? _GEN448 : _GEN444;
wire  _GEN450 = io_x[18] ? _GEN449 : _GEN441;
wire  _GEN451 = io_x[33] ? _GEN450 : _GEN437;
wire  _GEN452 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN453 = io_x[19] ? _GEN345 : _GEN452;
wire  _GEN454 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN455 = io_x[27] ? _GEN454 : _GEN336;
wire  _GEN456 = io_x[19] ? _GEN455 : _GEN338;
wire  _GEN457 = io_x[23] ? _GEN456 : _GEN453;
wire  _GEN458 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN459 = io_x[27] ? _GEN343 : _GEN458;
wire  _GEN460 = io_x[19] ? _GEN459 : _GEN345;
wire  _GEN461 = io_x[23] ? _GEN460 : _GEN370;
wire  _GEN462 = io_x[18] ? _GEN461 : _GEN457;
wire  _GEN463 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN464 = io_x[27] ? _GEN343 : _GEN463;
wire  _GEN465 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN466 = io_x[27] ? _GEN465 : _GEN343;
wire  _GEN467 = io_x[19] ? _GEN466 : _GEN464;
wire  _GEN468 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN469 = io_x[19] ? _GEN468 : _GEN345;
wire  _GEN470 = io_x[23] ? _GEN469 : _GEN467;
wire  _GEN471 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN472 = io_x[27] ? _GEN471 : _GEN343;
wire  _GEN473 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN474 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN475 = io_x[27] ? _GEN474 : _GEN473;
wire  _GEN476 = io_x[19] ? _GEN475 : _GEN472;
wire  _GEN477 = io_x[23] ? _GEN476 : _GEN332;
wire  _GEN478 = io_x[18] ? _GEN477 : _GEN470;
wire  _GEN479 = io_x[33] ? _GEN478 : _GEN462;
wire  _GEN480 = io_x[31] ? _GEN479 : _GEN451;
wire  _GEN481 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN482 = io_x[27] ? _GEN343 : _GEN481;
wire  _GEN483 = io_x[19] ? _GEN482 : _GEN345;
wire  _GEN484 = io_x[23] ? _GEN483 : _GEN332;
wire  _GEN485 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN486 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN487 = io_x[27] ? _GEN486 : _GEN336;
wire  _GEN488 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN489 = io_x[27] ? _GEN488 : _GEN343;
wire  _GEN490 = io_x[19] ? _GEN489 : _GEN487;
wire  _GEN491 = io_x[23] ? _GEN490 : _GEN485;
wire  _GEN492 = io_x[18] ? _GEN491 : _GEN484;
wire  _GEN493 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN494 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN495 = io_x[27] ? _GEN336 : _GEN494;
wire  _GEN496 = io_x[19] ? _GEN495 : _GEN345;
wire  _GEN497 = io_x[23] ? _GEN496 : _GEN493;
wire  _GEN498 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN499 = io_x[27] ? _GEN336 : _GEN498;
wire  _GEN500 = io_x[19] ? _GEN499 : _GEN338;
wire  _GEN501 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN502 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN503 = io_x[19] ? _GEN502 : _GEN501;
wire  _GEN504 = io_x[23] ? _GEN503 : _GEN500;
wire  _GEN505 = io_x[18] ? _GEN504 : _GEN497;
wire  _GEN506 = io_x[33] ? _GEN505 : _GEN492;
wire  _GEN507 = io_x[23] ? _GEN332 : _GEN370;
wire  _GEN508 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN509 = io_x[27] ? _GEN508 : _GEN336;
wire  _GEN510 = io_x[19] ? _GEN509 : _GEN345;
wire  _GEN511 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN512 = io_x[27] ? _GEN511 : _GEN343;
wire  _GEN513 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN514 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN515 = io_x[27] ? _GEN514 : _GEN513;
wire  _GEN516 = io_x[19] ? _GEN515 : _GEN512;
wire  _GEN517 = io_x[23] ? _GEN516 : _GEN510;
wire  _GEN518 = io_x[18] ? _GEN517 : _GEN507;
wire  _GEN519 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN520 = io_x[19] ? _GEN519 : _GEN345;
wire  _GEN521 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN522 = io_x[27] ? _GEN521 : _GEN343;
wire  _GEN523 = io_x[19] ? _GEN522 : _GEN345;
wire  _GEN524 = io_x[23] ? _GEN523 : _GEN520;
wire  _GEN525 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN526 = io_x[27] ? _GEN525 : _GEN343;
wire  _GEN527 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN528 = io_x[27] ? _GEN336 : _GEN527;
wire  _GEN529 = io_x[19] ? _GEN528 : _GEN526;
wire  _GEN530 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN531 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN532 = io_x[27] ? _GEN531 : _GEN530;
wire  _GEN533 = io_x[19] ? _GEN532 : _GEN338;
wire  _GEN534 = io_x[23] ? _GEN533 : _GEN529;
wire  _GEN535 = io_x[18] ? _GEN534 : _GEN524;
wire  _GEN536 = io_x[33] ? _GEN535 : _GEN518;
wire  _GEN537 = io_x[31] ? _GEN536 : _GEN506;
wire  _GEN538 = io_x[28] ? _GEN537 : _GEN480;
wire  _GEN539 = io_x[26] ? _GEN538 : _GEN432;
wire  _GEN540 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN541 = io_x[27] ? _GEN540 : _GEN343;
wire  _GEN542 = io_x[19] ? _GEN345 : _GEN541;
wire  _GEN543 = io_x[23] ? _GEN542 : _GEN332;
wire  _GEN544 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN545 = io_x[27] ? _GEN544 : _GEN343;
wire  _GEN546 = io_x[19] ? _GEN338 : _GEN545;
wire  _GEN547 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN548 = io_x[27] ? _GEN547 : _GEN343;
wire  _GEN549 = io_x[19] ? _GEN338 : _GEN548;
wire  _GEN550 = io_x[23] ? _GEN549 : _GEN546;
wire  _GEN551 = io_x[18] ? _GEN550 : _GEN543;
wire  _GEN552 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN553 = io_x[27] ? _GEN552 : _GEN343;
wire  _GEN554 = io_x[19] ? _GEN345 : _GEN553;
wire  _GEN555 = io_x[23] ? _GEN554 : _GEN332;
wire  _GEN556 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN557 = io_x[19] ? _GEN338 : _GEN556;
wire  _GEN558 = io_x[23] ? _GEN557 : _GEN370;
wire  _GEN559 = io_x[18] ? _GEN558 : _GEN555;
wire  _GEN560 = io_x[33] ? _GEN559 : _GEN551;
wire  _GEN561 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN562 = io_x[19] ? _GEN345 : _GEN561;
wire  _GEN563 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN564 = io_x[27] ? _GEN563 : _GEN343;
wire  _GEN565 = io_x[19] ? _GEN345 : _GEN564;
wire  _GEN566 = io_x[23] ? _GEN565 : _GEN562;
wire  _GEN567 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN568 = io_x[27] ? _GEN567 : _GEN336;
wire  _GEN569 = io_x[19] ? _GEN345 : _GEN568;
wire  _GEN570 = io_x[23] ? _GEN569 : _GEN370;
wire  _GEN571 = io_x[18] ? _GEN570 : _GEN566;
wire  _GEN572 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN573 = io_x[27] ? _GEN572 : _GEN336;
wire  _GEN574 = io_x[19] ? _GEN345 : _GEN573;
wire  _GEN575 = io_x[23] ? _GEN574 : _GEN332;
wire  _GEN576 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN577 = io_x[27] ? _GEN576 : _GEN336;
wire  _GEN578 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN579 = io_x[27] ? _GEN336 : _GEN578;
wire  _GEN580 = io_x[19] ? _GEN579 : _GEN577;
wire  _GEN581 = io_x[23] ? _GEN332 : _GEN580;
wire  _GEN582 = io_x[18] ? _GEN581 : _GEN575;
wire  _GEN583 = io_x[33] ? _GEN582 : _GEN571;
wire  _GEN584 = io_x[31] ? _GEN583 : _GEN560;
wire  _GEN585 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN586 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN587 = io_x[27] ? _GEN586 : _GEN343;
wire  _GEN588 = io_x[19] ? _GEN587 : _GEN585;
wire  _GEN589 = io_x[23] ? _GEN588 : _GEN332;
wire  _GEN590 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN591 = io_x[27] ? _GEN590 : _GEN336;
wire  _GEN592 = io_x[19] ? _GEN345 : _GEN591;
wire  _GEN593 = io_x[23] ? _GEN332 : _GEN592;
wire  _GEN594 = io_x[18] ? _GEN593 : _GEN589;
wire  _GEN595 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN596 = io_x[27] ? _GEN595 : _GEN343;
wire  _GEN597 = io_x[19] ? _GEN596 : _GEN345;
wire  _GEN598 = io_x[23] ? _GEN597 : _GEN370;
wire  _GEN599 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN600 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN601 = io_x[27] ? _GEN600 : _GEN599;
wire  _GEN602 = io_x[19] ? _GEN345 : _GEN601;
wire  _GEN603 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN604 = io_x[27] ? _GEN603 : _GEN343;
wire  _GEN605 = io_x[19] ? _GEN604 : _GEN345;
wire  _GEN606 = io_x[23] ? _GEN605 : _GEN602;
wire  _GEN607 = io_x[18] ? _GEN606 : _GEN598;
wire  _GEN608 = io_x[33] ? _GEN607 : _GEN594;
wire  _GEN609 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN610 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN611 = io_x[19] ? _GEN610 : _GEN609;
wire  _GEN612 = io_x[23] ? _GEN611 : _GEN332;
wire  _GEN613 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN614 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN615 = io_x[27] ? _GEN614 : _GEN613;
wire  _GEN616 = io_x[19] ? _GEN615 : _GEN338;
wire  _GEN617 = io_x[23] ? _GEN616 : _GEN332;
wire  _GEN618 = io_x[18] ? _GEN617 : _GEN612;
wire  _GEN619 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN620 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN621 = io_x[27] ? _GEN620 : _GEN336;
wire  _GEN622 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN623 = io_x[27] ? _GEN622 : _GEN336;
wire  _GEN624 = io_x[19] ? _GEN623 : _GEN621;
wire  _GEN625 = io_x[23] ? _GEN624 : _GEN619;
wire  _GEN626 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN627 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN628 = io_x[27] ? _GEN627 : _GEN626;
wire  _GEN629 = io_x[19] ? _GEN628 : _GEN338;
wire  _GEN630 = io_x[23] ? _GEN629 : _GEN370;
wire  _GEN631 = io_x[18] ? _GEN630 : _GEN625;
wire  _GEN632 = io_x[33] ? _GEN631 : _GEN618;
wire  _GEN633 = io_x[31] ? _GEN632 : _GEN608;
wire  _GEN634 = io_x[28] ? _GEN633 : _GEN584;
wire  _GEN635 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN636 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN637 = io_x[27] ? _GEN636 : _GEN343;
wire  _GEN638 = io_x[19] ? _GEN637 : _GEN635;
wire  _GEN639 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN640 = io_x[19] ? _GEN345 : _GEN639;
wire  _GEN641 = io_x[23] ? _GEN640 : _GEN638;
wire  _GEN642 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN643 = io_x[19] ? _GEN345 : _GEN642;
wire  _GEN644 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN645 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN646 = io_x[27] ? _GEN645 : _GEN644;
wire  _GEN647 = io_x[19] ? _GEN345 : _GEN646;
wire  _GEN648 = io_x[23] ? _GEN647 : _GEN643;
wire  _GEN649 = io_x[18] ? _GEN648 : _GEN641;
wire  _GEN650 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN651 = io_x[27] ? _GEN343 : _GEN650;
wire  _GEN652 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN653 = io_x[19] ? _GEN652 : _GEN651;
wire  _GEN654 = io_x[23] ? _GEN653 : _GEN370;
wire  _GEN655 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN656 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN657 = io_x[27] ? _GEN656 : _GEN343;
wire  _GEN658 = io_x[19] ? _GEN657 : _GEN338;
wire  _GEN659 = io_x[23] ? _GEN658 : _GEN655;
wire  _GEN660 = io_x[18] ? _GEN659 : _GEN654;
wire  _GEN661 = io_x[33] ? _GEN660 : _GEN649;
wire  _GEN662 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN663 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN664 = io_x[27] ? _GEN343 : _GEN663;
wire  _GEN665 = io_x[19] ? _GEN664 : _GEN345;
wire  _GEN666 = io_x[23] ? _GEN665 : _GEN662;
wire  _GEN667 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN668 = io_x[27] ? _GEN336 : _GEN667;
wire  _GEN669 = io_x[19] ? _GEN668 : _GEN345;
wire  _GEN670 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN671 = io_x[27] ? _GEN336 : _GEN670;
wire  _GEN672 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN673 = io_x[19] ? _GEN672 : _GEN671;
wire  _GEN674 = io_x[23] ? _GEN673 : _GEN669;
wire  _GEN675 = io_x[18] ? _GEN674 : _GEN666;
wire  _GEN676 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN677 = io_x[27] ? _GEN676 : _GEN336;
wire  _GEN678 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN679 = io_x[27] ? _GEN678 : _GEN336;
wire  _GEN680 = io_x[19] ? _GEN679 : _GEN677;
wire  _GEN681 = io_x[23] ? _GEN680 : _GEN332;
wire  _GEN682 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN683 = io_x[27] ? _GEN343 : _GEN682;
wire  _GEN684 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN685 = io_x[27] ? _GEN343 : _GEN684;
wire  _GEN686 = io_x[19] ? _GEN685 : _GEN683;
wire  _GEN687 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN688 = io_x[27] ? _GEN687 : _GEN336;
wire  _GEN689 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN690 = io_x[27] ? _GEN689 : _GEN343;
wire  _GEN691 = io_x[19] ? _GEN690 : _GEN688;
wire  _GEN692 = io_x[23] ? _GEN691 : _GEN686;
wire  _GEN693 = io_x[18] ? _GEN692 : _GEN681;
wire  _GEN694 = io_x[33] ? _GEN693 : _GEN675;
wire  _GEN695 = io_x[31] ? _GEN694 : _GEN661;
wire  _GEN696 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN697 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN698 = io_x[19] ? _GEN345 : _GEN697;
wire  _GEN699 = io_x[23] ? _GEN698 : _GEN696;
wire  _GEN700 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN701 = io_x[27] ? _GEN700 : _GEN336;
wire  _GEN702 = io_x[19] ? _GEN701 : _GEN338;
wire  _GEN703 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN704 = io_x[23] ? _GEN703 : _GEN702;
wire  _GEN705 = io_x[18] ? _GEN704 : _GEN699;
wire  _GEN706 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN707 = io_x[27] ? _GEN706 : _GEN336;
wire  _GEN708 = io_x[19] ? _GEN345 : _GEN707;
wire  _GEN709 = io_x[23] ? _GEN708 : _GEN370;
wire  _GEN710 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN711 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN712 = io_x[27] ? _GEN343 : _GEN711;
wire  _GEN713 = io_x[19] ? _GEN712 : _GEN710;
wire  _GEN714 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN715 = io_x[23] ? _GEN714 : _GEN713;
wire  _GEN716 = io_x[18] ? _GEN715 : _GEN709;
wire  _GEN717 = io_x[33] ? _GEN716 : _GEN705;
wire  _GEN718 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN719 = io_x[27] ? _GEN343 : _GEN718;
wire  _GEN720 = io_x[19] ? _GEN719 : _GEN338;
wire  _GEN721 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN722 = io_x[27] ? _GEN721 : _GEN343;
wire  _GEN723 = io_x[19] ? _GEN338 : _GEN722;
wire  _GEN724 = io_x[23] ? _GEN723 : _GEN720;
wire  _GEN725 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN726 = io_x[19] ? _GEN338 : _GEN725;
wire  _GEN727 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN728 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN729 = io_x[27] ? _GEN728 : _GEN727;
wire  _GEN730 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN731 = io_x[19] ? _GEN730 : _GEN729;
wire  _GEN732 = io_x[23] ? _GEN731 : _GEN726;
wire  _GEN733 = io_x[18] ? _GEN732 : _GEN724;
wire  _GEN734 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN735 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN736 = io_x[27] ? _GEN735 : _GEN343;
wire  _GEN737 = io_x[19] ? _GEN736 : _GEN734;
wire  _GEN738 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN739 = io_x[27] ? _GEN738 : _GEN343;
wire  _GEN740 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN741 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN742 = io_x[27] ? _GEN741 : _GEN740;
wire  _GEN743 = io_x[19] ? _GEN742 : _GEN739;
wire  _GEN744 = io_x[23] ? _GEN743 : _GEN737;
wire  _GEN745 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN746 = io_x[27] ? _GEN343 : _GEN745;
wire  _GEN747 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN748 = io_x[27] ? _GEN747 : _GEN343;
wire  _GEN749 = io_x[19] ? _GEN748 : _GEN746;
wire  _GEN750 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN751 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN752 = io_x[27] ? _GEN751 : _GEN750;
wire  _GEN753 = io_x[19] ? _GEN752 : _GEN345;
wire  _GEN754 = io_x[23] ? _GEN753 : _GEN749;
wire  _GEN755 = io_x[18] ? _GEN754 : _GEN744;
wire  _GEN756 = io_x[33] ? _GEN755 : _GEN733;
wire  _GEN757 = io_x[31] ? _GEN756 : _GEN717;
wire  _GEN758 = io_x[28] ? _GEN757 : _GEN695;
wire  _GEN759 = io_x[26] ? _GEN758 : _GEN634;
wire  _GEN760 = io_x[20] ? _GEN759 : _GEN539;
wire  _GEN761 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN762 = io_x[19] ? _GEN761 : _GEN345;
wire  _GEN763 = io_x[23] ? _GEN762 : _GEN332;
wire  _GEN764 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN765 = io_x[19] ? _GEN764 : _GEN345;
wire  _GEN766 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN767 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN768 = io_x[19] ? _GEN767 : _GEN766;
wire  _GEN769 = io_x[23] ? _GEN768 : _GEN765;
wire  _GEN770 = io_x[18] ? _GEN769 : _GEN763;
wire  _GEN771 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN772 = io_x[27] ? _GEN771 : _GEN343;
wire  _GEN773 = io_x[19] ? _GEN345 : _GEN772;
wire  _GEN774 = io_x[23] ? _GEN370 : _GEN773;
wire  _GEN775 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN776 = io_x[27] ? _GEN775 : _GEN336;
wire  _GEN777 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN778 = io_x[19] ? _GEN777 : _GEN776;
wire  _GEN779 = io_x[23] ? _GEN778 : _GEN370;
wire  _GEN780 = io_x[18] ? _GEN779 : _GEN774;
wire  _GEN781 = io_x[33] ? _GEN780 : _GEN770;
wire  _GEN782 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN783 = io_x[23] ? _GEN332 : _GEN782;
wire  _GEN784 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN785 = io_x[23] ? _GEN784 : _GEN332;
wire  _GEN786 = io_x[18] ? _GEN785 : _GEN783;
wire  _GEN787 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN788 = io_x[27] ? _GEN787 : _GEN343;
wire  _GEN789 = io_x[19] ? _GEN788 : _GEN345;
wire  _GEN790 = io_x[23] ? _GEN789 : _GEN332;
wire  _GEN791 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN792 = io_x[27] ? _GEN791 : _GEN343;
wire  _GEN793 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN794 = io_x[27] ? _GEN793 : _GEN343;
wire  _GEN795 = io_x[19] ? _GEN794 : _GEN792;
wire  _GEN796 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN797 = io_x[27] ? _GEN796 : _GEN343;
wire  _GEN798 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN799 = io_x[19] ? _GEN798 : _GEN797;
wire  _GEN800 = io_x[23] ? _GEN799 : _GEN795;
wire  _GEN801 = io_x[18] ? _GEN800 : _GEN790;
wire  _GEN802 = io_x[33] ? _GEN801 : _GEN786;
wire  _GEN803 = io_x[31] ? _GEN802 : _GEN781;
wire  _GEN804 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN805 = io_x[27] ? _GEN804 : _GEN343;
wire  _GEN806 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN807 = io_x[27] ? _GEN806 : _GEN336;
wire  _GEN808 = io_x[19] ? _GEN807 : _GEN805;
wire  _GEN809 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN810 = io_x[27] ? _GEN809 : _GEN343;
wire  _GEN811 = io_x[19] ? _GEN338 : _GEN810;
wire  _GEN812 = io_x[23] ? _GEN811 : _GEN808;
wire  _GEN813 = io_x[18] ? _GEN812 : _GEN331;
wire  _GEN814 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN815 = io_x[23] ? _GEN332 : _GEN814;
wire  _GEN816 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN817 = io_x[27] ? _GEN816 : _GEN336;
wire  _GEN818 = io_x[19] ? _GEN817 : _GEN345;
wire  _GEN819 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN820 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN821 = io_x[27] ? _GEN820 : _GEN343;
wire  _GEN822 = io_x[19] ? _GEN821 : _GEN819;
wire  _GEN823 = io_x[23] ? _GEN822 : _GEN818;
wire  _GEN824 = io_x[18] ? _GEN823 : _GEN815;
wire  _GEN825 = io_x[33] ? _GEN824 : _GEN813;
wire  _GEN826 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN827 = io_x[27] ? _GEN343 : _GEN826;
wire  _GEN828 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN829 = io_x[19] ? _GEN828 : _GEN827;
wire  _GEN830 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN831 = io_x[23] ? _GEN830 : _GEN829;
wire  _GEN832 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN833 = io_x[27] ? _GEN336 : _GEN832;
wire  _GEN834 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN835 = io_x[27] ? _GEN343 : _GEN834;
wire  _GEN836 = io_x[19] ? _GEN835 : _GEN833;
wire  _GEN837 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN838 = io_x[27] ? _GEN837 : _GEN343;
wire  _GEN839 = io_x[19] ? _GEN338 : _GEN838;
wire  _GEN840 = io_x[23] ? _GEN839 : _GEN836;
wire  _GEN841 = io_x[18] ? _GEN840 : _GEN831;
wire  _GEN842 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN843 = io_x[27] ? _GEN343 : _GEN842;
wire  _GEN844 = io_x[19] ? _GEN843 : _GEN345;
wire  _GEN845 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN846 = io_x[27] ? _GEN343 : _GEN845;
wire  _GEN847 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN848 = io_x[19] ? _GEN847 : _GEN846;
wire  _GEN849 = io_x[23] ? _GEN848 : _GEN844;
wire  _GEN850 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN851 = io_x[27] ? _GEN343 : _GEN850;
wire  _GEN852 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN853 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN854 = io_x[27] ? _GEN853 : _GEN852;
wire  _GEN855 = io_x[19] ? _GEN854 : _GEN851;
wire  _GEN856 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN857 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN858 = io_x[27] ? _GEN857 : _GEN856;
wire  _GEN859 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN860 = io_x[27] ? _GEN859 : _GEN343;
wire  _GEN861 = io_x[19] ? _GEN860 : _GEN858;
wire  _GEN862 = io_x[23] ? _GEN861 : _GEN855;
wire  _GEN863 = io_x[18] ? _GEN862 : _GEN849;
wire  _GEN864 = io_x[33] ? _GEN863 : _GEN841;
wire  _GEN865 = io_x[31] ? _GEN864 : _GEN825;
wire  _GEN866 = io_x[28] ? _GEN865 : _GEN803;
wire  _GEN867 = io_x[23] ? _GEN332 : _GEN370;
wire  _GEN868 = io_x[18] ? _GEN362 : _GEN867;
wire  _GEN869 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN870 = io_x[19] ? _GEN338 : _GEN869;
wire  _GEN871 = io_x[23] ? _GEN332 : _GEN870;
wire  _GEN872 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN873 = io_x[27] ? _GEN336 : _GEN872;
wire  _GEN874 = io_x[19] ? _GEN338 : _GEN873;
wire  _GEN875 = io_x[23] ? _GEN332 : _GEN874;
wire  _GEN876 = io_x[18] ? _GEN875 : _GEN871;
wire  _GEN877 = io_x[33] ? _GEN876 : _GEN868;
wire  _GEN878 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN879 = io_x[27] ? _GEN336 : _GEN878;
wire  _GEN880 = io_x[19] ? _GEN879 : _GEN345;
wire  _GEN881 = io_x[23] ? _GEN370 : _GEN880;
wire  _GEN882 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN883 = io_x[27] ? _GEN882 : _GEN343;
wire  _GEN884 = io_x[19] ? _GEN345 : _GEN883;
wire  _GEN885 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN886 = io_x[27] ? _GEN885 : _GEN336;
wire  _GEN887 = io_x[19] ? _GEN886 : _GEN345;
wire  _GEN888 = io_x[23] ? _GEN887 : _GEN884;
wire  _GEN889 = io_x[18] ? _GEN888 : _GEN881;
wire  _GEN890 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN891 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN892 = io_x[27] ? _GEN891 : _GEN890;
wire  _GEN893 = io_x[19] ? _GEN892 : _GEN338;
wire  _GEN894 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN895 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN896 = io_x[27] ? _GEN895 : _GEN894;
wire  _GEN897 = io_x[19] ? _GEN896 : _GEN338;
wire  _GEN898 = io_x[23] ? _GEN897 : _GEN893;
wire  _GEN899 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN900 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN901 = io_x[27] ? _GEN900 : _GEN899;
wire  _GEN902 = io_x[19] ? _GEN901 : _GEN345;
wire  _GEN903 = io_x[23] ? _GEN902 : _GEN370;
wire  _GEN904 = io_x[18] ? _GEN903 : _GEN898;
wire  _GEN905 = io_x[33] ? _GEN904 : _GEN889;
wire  _GEN906 = io_x[31] ? _GEN905 : _GEN877;
wire  _GEN907 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN908 = io_x[27] ? _GEN343 : _GEN907;
wire  _GEN909 = io_x[19] ? _GEN908 : _GEN345;
wire  _GEN910 = io_x[23] ? _GEN370 : _GEN909;
wire  _GEN911 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN912 = io_x[27] ? _GEN911 : _GEN343;
wire  _GEN913 = io_x[19] ? _GEN338 : _GEN912;
wire  _GEN914 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN915 = io_x[27] ? _GEN914 : _GEN343;
wire  _GEN916 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN917 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN918 = io_x[27] ? _GEN917 : _GEN916;
wire  _GEN919 = io_x[19] ? _GEN918 : _GEN915;
wire  _GEN920 = io_x[23] ? _GEN919 : _GEN913;
wire  _GEN921 = io_x[18] ? _GEN920 : _GEN910;
wire  _GEN922 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN923 = io_x[27] ? _GEN343 : _GEN922;
wire  _GEN924 = io_x[19] ? _GEN923 : _GEN345;
wire  _GEN925 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN926 = io_x[27] ? _GEN925 : _GEN343;
wire  _GEN927 = io_x[19] ? _GEN926 : _GEN345;
wire  _GEN928 = io_x[23] ? _GEN927 : _GEN924;
wire  _GEN929 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN930 = io_x[19] ? _GEN338 : _GEN929;
wire  _GEN931 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN932 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN933 = io_x[27] ? _GEN932 : _GEN931;
wire  _GEN934 = io_x[19] ? _GEN933 : _GEN338;
wire  _GEN935 = io_x[23] ? _GEN934 : _GEN930;
wire  _GEN936 = io_x[18] ? _GEN935 : _GEN928;
wire  _GEN937 = io_x[33] ? _GEN936 : _GEN921;
wire  _GEN938 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN939 = io_x[27] ? _GEN938 : _GEN343;
wire  _GEN940 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN941 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN942 = io_x[27] ? _GEN941 : _GEN940;
wire  _GEN943 = io_x[19] ? _GEN942 : _GEN939;
wire  _GEN944 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN945 = io_x[27] ? _GEN944 : _GEN343;
wire  _GEN946 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN947 = io_x[19] ? _GEN946 : _GEN945;
wire  _GEN948 = io_x[23] ? _GEN947 : _GEN943;
wire  _GEN949 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN950 = io_x[19] ? _GEN345 : _GEN949;
wire  _GEN951 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN952 = io_x[27] ? _GEN951 : _GEN336;
wire  _GEN953 = io_x[19] ? _GEN952 : _GEN345;
wire  _GEN954 = io_x[23] ? _GEN953 : _GEN950;
wire  _GEN955 = io_x[18] ? _GEN954 : _GEN948;
wire  _GEN956 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN957 = io_x[27] ? _GEN956 : _GEN940;
wire  _GEN958 = io_x[19] ? _GEN957 : _GEN338;
wire  _GEN959 = io_x[27] ? _GEN944 : _GEN343;
wire  _GEN960 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN961 = io_x[27] ? _GEN960 : _GEN336;
wire  _GEN962 = io_x[19] ? _GEN961 : _GEN959;
wire  _GEN963 = io_x[23] ? _GEN962 : _GEN958;
wire  _GEN964 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN965 = io_x[27] ? _GEN336 : _GEN964;
wire  _GEN966 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN967 = io_x[27] ? _GEN966 : _GEN343;
wire  _GEN968 = io_x[19] ? _GEN967 : _GEN965;
wire  _GEN969 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN970 = io_x[27] ? _GEN969 : _GEN343;
wire  _GEN971 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN972 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN973 = io_x[27] ? _GEN972 : _GEN971;
wire  _GEN974 = io_x[19] ? _GEN973 : _GEN970;
wire  _GEN975 = io_x[23] ? _GEN974 : _GEN968;
wire  _GEN976 = io_x[18] ? _GEN975 : _GEN963;
wire  _GEN977 = io_x[33] ? _GEN976 : _GEN955;
wire  _GEN978 = io_x[31] ? _GEN977 : _GEN937;
wire  _GEN979 = io_x[28] ? _GEN978 : _GEN906;
wire  _GEN980 = io_x[26] ? _GEN979 : _GEN866;
wire  _GEN981 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN982 = io_x[27] ? _GEN981 : _GEN343;
wire  _GEN983 = io_x[19] ? _GEN982 : _GEN345;
wire  _GEN984 = io_x[23] ? _GEN983 : _GEN370;
wire  _GEN985 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN986 = io_x[27] ? _GEN985 : _GEN343;
wire  _GEN987 = io_x[19] ? _GEN345 : _GEN986;
wire  _GEN988 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN989 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN990 = io_x[27] ? _GEN989 : _GEN343;
wire  _GEN991 = io_x[19] ? _GEN990 : _GEN988;
wire  _GEN992 = io_x[23] ? _GEN991 : _GEN987;
wire  _GEN993 = io_x[18] ? _GEN992 : _GEN984;
wire  _GEN994 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN995 = io_x[27] ? _GEN994 : _GEN336;
wire  _GEN996 = io_x[19] ? _GEN345 : _GEN995;
wire  _GEN997 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN998 = io_x[27] ? _GEN997 : _GEN343;
wire  _GEN999 = io_x[19] ? _GEN998 : _GEN345;
wire  _GEN1000 = io_x[23] ? _GEN999 : _GEN996;
wire  _GEN1001 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1002 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1003 = io_x[27] ? _GEN1002 : _GEN343;
wire  _GEN1004 = io_x[19] ? _GEN1003 : _GEN338;
wire  _GEN1005 = io_x[23] ? _GEN1004 : _GEN1001;
wire  _GEN1006 = io_x[18] ? _GEN1005 : _GEN1000;
wire  _GEN1007 = io_x[33] ? _GEN1006 : _GEN993;
wire  _GEN1008 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1009 = io_x[19] ? _GEN338 : _GEN1008;
wire  _GEN1010 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1011 = io_x[19] ? _GEN345 : _GEN1010;
wire  _GEN1012 = io_x[23] ? _GEN1011 : _GEN1009;
wire  _GEN1013 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1014 = io_x[27] ? _GEN1013 : _GEN343;
wire  _GEN1015 = io_x[19] ? _GEN345 : _GEN1014;
wire  _GEN1016 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN1017 = io_x[23] ? _GEN1016 : _GEN1015;
wire  _GEN1018 = io_x[18] ? _GEN1017 : _GEN1012;
wire  _GEN1019 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1020 = io_x[27] ? _GEN1019 : _GEN343;
wire  _GEN1021 = io_x[19] ? _GEN338 : _GEN1020;
wire  _GEN1022 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1023 = io_x[27] ? _GEN1022 : _GEN343;
wire  _GEN1024 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1025 = io_x[27] ? _GEN1024 : _GEN343;
wire  _GEN1026 = io_x[19] ? _GEN1025 : _GEN1023;
wire  _GEN1027 = io_x[23] ? _GEN1026 : _GEN1021;
wire  _GEN1028 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1029 = io_x[27] ? _GEN1028 : _GEN343;
wire  _GEN1030 = io_x[19] ? _GEN345 : _GEN1029;
wire  _GEN1031 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1032 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1033 = io_x[27] ? _GEN1032 : _GEN1031;
wire  _GEN1034 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1035 = io_x[27] ? _GEN1034 : _GEN343;
wire  _GEN1036 = io_x[19] ? _GEN1035 : _GEN1033;
wire  _GEN1037 = io_x[23] ? _GEN1036 : _GEN1030;
wire  _GEN1038 = io_x[18] ? _GEN1037 : _GEN1027;
wire  _GEN1039 = io_x[33] ? _GEN1038 : _GEN1018;
wire  _GEN1040 = io_x[31] ? _GEN1039 : _GEN1007;
wire  _GEN1041 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1042 = io_x[19] ? _GEN1041 : _GEN345;
wire  _GEN1043 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1044 = io_x[27] ? _GEN1043 : _GEN343;
wire  _GEN1045 = io_x[19] ? _GEN345 : _GEN1044;
wire  _GEN1046 = io_x[23] ? _GEN1045 : _GEN1042;
wire  _GEN1047 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1048 = io_x[27] ? _GEN1047 : _GEN343;
wire  _GEN1049 = io_x[19] ? _GEN1048 : _GEN345;
wire  _GEN1050 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1051 = io_x[19] ? _GEN1050 : _GEN338;
wire  _GEN1052 = io_x[23] ? _GEN1051 : _GEN1049;
wire  _GEN1053 = io_x[18] ? _GEN1052 : _GEN1046;
wire  _GEN1054 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1055 = io_x[19] ? _GEN1054 : _GEN345;
wire  _GEN1056 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1057 = io_x[27] ? _GEN1056 : _GEN343;
wire  _GEN1058 = io_x[19] ? _GEN1057 : _GEN338;
wire  _GEN1059 = io_x[23] ? _GEN1058 : _GEN1055;
wire  _GEN1060 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1061 = io_x[27] ? _GEN1060 : _GEN336;
wire  _GEN1062 = io_x[19] ? _GEN1061 : _GEN345;
wire  _GEN1063 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1064 = io_x[27] ? _GEN1063 : _GEN343;
wire  _GEN1065 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1066 = io_x[27] ? _GEN1065 : _GEN336;
wire  _GEN1067 = io_x[19] ? _GEN1066 : _GEN1064;
wire  _GEN1068 = io_x[23] ? _GEN1067 : _GEN1062;
wire  _GEN1069 = io_x[18] ? _GEN1068 : _GEN1059;
wire  _GEN1070 = io_x[33] ? _GEN1069 : _GEN1053;
wire  _GEN1071 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1072 = io_x[27] ? _GEN343 : _GEN1071;
wire  _GEN1073 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1074 = io_x[19] ? _GEN1073 : _GEN1072;
wire  _GEN1075 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1076 = io_x[27] ? _GEN1075 : _GEN343;
wire  _GEN1077 = io_x[19] ? _GEN338 : _GEN1076;
wire  _GEN1078 = io_x[23] ? _GEN1077 : _GEN1074;
wire  _GEN1079 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1080 = io_x[27] ? _GEN336 : _GEN1079;
wire  _GEN1081 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1082 = io_x[27] ? _GEN1081 : _GEN343;
wire  _GEN1083 = io_x[19] ? _GEN1082 : _GEN1080;
wire  _GEN1084 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1085 = io_x[27] ? _GEN336 : _GEN1084;
wire  _GEN1086 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1087 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1088 = io_x[27] ? _GEN1087 : _GEN1086;
wire  _GEN1089 = io_x[19] ? _GEN1088 : _GEN1085;
wire  _GEN1090 = io_x[23] ? _GEN1089 : _GEN1083;
wire  _GEN1091 = io_x[18] ? _GEN1090 : _GEN1078;
wire  _GEN1092 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1093 = io_x[27] ? _GEN343 : _GEN1092;
wire  _GEN1094 = io_x[19] ? _GEN1093 : _GEN345;
wire  _GEN1095 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1096 = io_x[27] ? _GEN1095 : _GEN343;
wire  _GEN1097 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1098 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1099 = io_x[27] ? _GEN1098 : _GEN1097;
wire  _GEN1100 = io_x[19] ? _GEN1099 : _GEN1096;
wire  _GEN1101 = io_x[23] ? _GEN1100 : _GEN1094;
wire  _GEN1102 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1103 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1104 = io_x[27] ? _GEN1103 : _GEN1102;
wire  _GEN1105 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1106 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1107 = io_x[27] ? _GEN1106 : _GEN1105;
wire  _GEN1108 = io_x[19] ? _GEN1107 : _GEN1104;
wire  _GEN1109 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1110 = io_x[27] ? _GEN1109 : _GEN343;
wire  _GEN1111 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1112 = io_x[27] ? _GEN1111 : _GEN343;
wire  _GEN1113 = io_x[19] ? _GEN1112 : _GEN1110;
wire  _GEN1114 = io_x[23] ? _GEN1113 : _GEN1108;
wire  _GEN1115 = io_x[18] ? _GEN1114 : _GEN1101;
wire  _GEN1116 = io_x[33] ? _GEN1115 : _GEN1091;
wire  _GEN1117 = io_x[31] ? _GEN1116 : _GEN1070;
wire  _GEN1118 = io_x[28] ? _GEN1117 : _GEN1040;
wire  _GEN1119 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1120 = io_x[27] ? _GEN1119 : _GEN343;
wire  _GEN1121 = io_x[19] ? _GEN1120 : _GEN345;
wire  _GEN1122 = io_x[23] ? _GEN1121 : _GEN332;
wire  _GEN1123 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1124 = io_x[27] ? _GEN1123 : _GEN343;
wire  _GEN1125 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1126 = io_x[27] ? _GEN1125 : _GEN343;
wire  _GEN1127 = io_x[19] ? _GEN1126 : _GEN1124;
wire  _GEN1128 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1129 = io_x[27] ? _GEN336 : _GEN1128;
wire  _GEN1130 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1131 = io_x[19] ? _GEN1130 : _GEN1129;
wire  _GEN1132 = io_x[23] ? _GEN1131 : _GEN1127;
wire  _GEN1133 = io_x[18] ? _GEN1132 : _GEN1122;
wire  _GEN1134 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1135 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1136 = io_x[27] ? _GEN1135 : _GEN1134;
wire  _GEN1137 = io_x[19] ? _GEN1136 : _GEN338;
wire  _GEN1138 = io_x[23] ? _GEN370 : _GEN1137;
wire  _GEN1139 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1140 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1141 = io_x[27] ? _GEN1140 : _GEN1139;
wire  _GEN1142 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1143 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1144 = io_x[27] ? _GEN1143 : _GEN1142;
wire  _GEN1145 = io_x[19] ? _GEN1144 : _GEN1141;
wire  _GEN1146 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1147 = io_x[27] ? _GEN336 : _GEN1146;
wire  _GEN1148 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1149 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1150 = io_x[27] ? _GEN1149 : _GEN1148;
wire  _GEN1151 = io_x[19] ? _GEN1150 : _GEN1147;
wire  _GEN1152 = io_x[23] ? _GEN1151 : _GEN1145;
wire  _GEN1153 = io_x[18] ? _GEN1152 : _GEN1138;
wire  _GEN1154 = io_x[33] ? _GEN1153 : _GEN1133;
wire  _GEN1155 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1156 = io_x[27] ? _GEN336 : _GEN1155;
wire  _GEN1157 = io_x[19] ? _GEN1156 : _GEN345;
wire  _GEN1158 = io_x[23] ? _GEN332 : _GEN1157;
wire  _GEN1159 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1160 = io_x[27] ? _GEN1159 : _GEN343;
wire  _GEN1161 = io_x[19] ? _GEN1160 : _GEN345;
wire  _GEN1162 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1163 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1164 = io_x[27] ? _GEN1163 : _GEN336;
wire  _GEN1165 = io_x[19] ? _GEN1164 : _GEN1162;
wire  _GEN1166 = io_x[23] ? _GEN1165 : _GEN1161;
wire  _GEN1167 = io_x[18] ? _GEN1166 : _GEN1158;
wire  _GEN1168 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1169 = io_x[27] ? _GEN1168 : _GEN343;
wire  _GEN1170 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1171 = io_x[27] ? _GEN336 : _GEN1170;
wire  _GEN1172 = io_x[19] ? _GEN1171 : _GEN1169;
wire  _GEN1173 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1174 = io_x[27] ? _GEN1173 : _GEN343;
wire  _GEN1175 = io_x[19] ? _GEN1174 : _GEN338;
wire  _GEN1176 = io_x[23] ? _GEN1175 : _GEN1172;
wire  _GEN1177 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1178 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1179 = io_x[27] ? _GEN1178 : _GEN1177;
wire  _GEN1180 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1181 = io_x[27] ? _GEN1180 : _GEN343;
wire  _GEN1182 = io_x[19] ? _GEN1181 : _GEN1179;
wire  _GEN1183 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1184 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1185 = io_x[27] ? _GEN1184 : _GEN1183;
wire  _GEN1186 = io_x[19] ? _GEN1185 : _GEN345;
wire  _GEN1187 = io_x[23] ? _GEN1186 : _GEN1182;
wire  _GEN1188 = io_x[18] ? _GEN1187 : _GEN1176;
wire  _GEN1189 = io_x[33] ? _GEN1188 : _GEN1167;
wire  _GEN1190 = io_x[31] ? _GEN1189 : _GEN1154;
wire  _GEN1191 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1192 = io_x[27] ? _GEN1191 : _GEN336;
wire  _GEN1193 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1194 = io_x[27] ? _GEN343 : _GEN1193;
wire  _GEN1195 = io_x[19] ? _GEN1194 : _GEN1192;
wire  _GEN1196 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1197 = io_x[27] ? _GEN1196 : _GEN343;
wire  _GEN1198 = io_x[19] ? _GEN345 : _GEN1197;
wire  _GEN1199 = io_x[23] ? _GEN1198 : _GEN1195;
wire  _GEN1200 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1201 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1202 = io_x[27] ? _GEN1201 : _GEN1200;
wire  _GEN1203 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1204 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1205 = io_x[27] ? _GEN1204 : _GEN1203;
wire  _GEN1206 = io_x[19] ? _GEN1205 : _GEN1202;
wire  _GEN1207 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1208 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1209 = io_x[27] ? _GEN1208 : _GEN1207;
wire  _GEN1210 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1211 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1212 = io_x[27] ? _GEN1211 : _GEN1210;
wire  _GEN1213 = io_x[19] ? _GEN1212 : _GEN1209;
wire  _GEN1214 = io_x[23] ? _GEN1213 : _GEN1206;
wire  _GEN1215 = io_x[18] ? _GEN1214 : _GEN1199;
wire  _GEN1216 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1217 = io_x[27] ? _GEN1216 : _GEN336;
wire  _GEN1218 = io_x[19] ? _GEN1217 : _GEN338;
wire  _GEN1219 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1220 = io_x[19] ? _GEN1219 : _GEN345;
wire  _GEN1221 = io_x[23] ? _GEN1220 : _GEN1218;
wire  _GEN1222 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1223 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1224 = io_x[27] ? _GEN1223 : _GEN1222;
wire  _GEN1225 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1226 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1227 = io_x[27] ? _GEN1226 : _GEN1225;
wire  _GEN1228 = io_x[19] ? _GEN1227 : _GEN1224;
wire  _GEN1229 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1230 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1231 = io_x[27] ? _GEN1230 : _GEN1229;
wire  _GEN1232 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1233 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1234 = io_x[27] ? _GEN1233 : _GEN1232;
wire  _GEN1235 = io_x[19] ? _GEN1234 : _GEN1231;
wire  _GEN1236 = io_x[23] ? _GEN1235 : _GEN1228;
wire  _GEN1237 = io_x[18] ? _GEN1236 : _GEN1221;
wire  _GEN1238 = io_x[33] ? _GEN1237 : _GEN1215;
wire  _GEN1239 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1240 = io_x[27] ? _GEN1239 : _GEN343;
wire  _GEN1241 = io_x[19] ? _GEN1240 : _GEN345;
wire  _GEN1242 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1243 = io_x[27] ? _GEN1242 : _GEN343;
wire  _GEN1244 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1245 = io_x[27] ? _GEN1244 : _GEN343;
wire  _GEN1246 = io_x[19] ? _GEN1245 : _GEN1243;
wire  _GEN1247 = io_x[23] ? _GEN1246 : _GEN1241;
wire  _GEN1248 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1249 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1250 = io_x[27] ? _GEN1249 : _GEN1248;
wire  _GEN1251 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1252 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1253 = io_x[27] ? _GEN1252 : _GEN1251;
wire  _GEN1254 = io_x[19] ? _GEN1253 : _GEN1250;
wire  _GEN1255 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1256 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1257 = io_x[27] ? _GEN1256 : _GEN1255;
wire  _GEN1258 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1259 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1260 = io_x[27] ? _GEN1259 : _GEN1258;
wire  _GEN1261 = io_x[19] ? _GEN1260 : _GEN1257;
wire  _GEN1262 = io_x[23] ? _GEN1261 : _GEN1254;
wire  _GEN1263 = io_x[18] ? _GEN1262 : _GEN1247;
wire  _GEN1264 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1265 = io_x[27] ? _GEN1264 : _GEN343;
wire  _GEN1266 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1267 = io_x[19] ? _GEN1266 : _GEN1265;
wire  _GEN1268 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1269 = io_x[27] ? _GEN1268 : _GEN336;
wire  _GEN1270 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1271 = io_x[27] ? _GEN1270 : _GEN343;
wire  _GEN1272 = io_x[19] ? _GEN1271 : _GEN1269;
wire  _GEN1273 = io_x[23] ? _GEN1272 : _GEN1267;
wire  _GEN1274 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1275 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1276 = io_x[27] ? _GEN1275 : _GEN1274;
wire  _GEN1277 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1278 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1279 = io_x[27] ? _GEN1278 : _GEN1277;
wire  _GEN1280 = io_x[19] ? _GEN1279 : _GEN1276;
wire  _GEN1281 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1282 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1283 = io_x[27] ? _GEN1282 : _GEN1281;
wire  _GEN1284 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1285 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1286 = io_x[27] ? _GEN1285 : _GEN1284;
wire  _GEN1287 = io_x[19] ? _GEN1286 : _GEN1283;
wire  _GEN1288 = io_x[23] ? _GEN1287 : _GEN1280;
wire  _GEN1289 = io_x[18] ? _GEN1288 : _GEN1273;
wire  _GEN1290 = io_x[33] ? _GEN1289 : _GEN1263;
wire  _GEN1291 = io_x[31] ? _GEN1290 : _GEN1238;
wire  _GEN1292 = io_x[28] ? _GEN1291 : _GEN1190;
wire  _GEN1293 = io_x[26] ? _GEN1292 : _GEN1118;
wire  _GEN1294 = io_x[20] ? _GEN1293 : _GEN980;
wire  _GEN1295 = io_x[24] ? _GEN1294 : _GEN760;
wire  _GEN1296 = io_x[18] ? _GEN362 : _GEN331;
wire  _GEN1297 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1298 = io_x[27] ? _GEN1297 : _GEN343;
wire  _GEN1299 = io_x[19] ? _GEN1298 : _GEN345;
wire  _GEN1300 = io_x[23] ? _GEN1299 : _GEN370;
wire  _GEN1301 = io_x[18] ? _GEN362 : _GEN1300;
wire  _GEN1302 = io_x[33] ? _GEN1301 : _GEN1296;
wire  _GEN1303 = io_x[23] ? _GEN332 : _GEN370;
wire  _GEN1304 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1305 = io_x[27] ? _GEN1304 : _GEN343;
wire  _GEN1306 = io_x[19] ? _GEN1305 : _GEN338;
wire  _GEN1307 = io_x[23] ? _GEN1306 : _GEN332;
wire  _GEN1308 = io_x[18] ? _GEN1307 : _GEN1303;
wire  _GEN1309 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1310 = io_x[19] ? _GEN1309 : _GEN345;
wire  _GEN1311 = io_x[23] ? _GEN332 : _GEN1310;
wire  _GEN1312 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1313 = io_x[27] ? _GEN1312 : _GEN343;
wire  _GEN1314 = io_x[19] ? _GEN1313 : _GEN345;
wire  _GEN1315 = io_x[23] ? _GEN1314 : _GEN332;
wire  _GEN1316 = io_x[18] ? _GEN1315 : _GEN1311;
wire  _GEN1317 = io_x[33] ? _GEN1316 : _GEN1308;
wire  _GEN1318 = io_x[31] ? _GEN1317 : _GEN1302;
wire  _GEN1319 = io_x[23] ? _GEN332 : _GEN370;
wire  _GEN1320 = io_x[18] ? _GEN1319 : _GEN331;
wire  _GEN1321 = io_x[23] ? _GEN332 : _GEN370;
wire  _GEN1322 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1323 = io_x[19] ? _GEN1322 : _GEN345;
wire  _GEN1324 = io_x[23] ? _GEN1323 : _GEN332;
wire  _GEN1325 = io_x[18] ? _GEN1324 : _GEN1321;
wire  _GEN1326 = io_x[33] ? _GEN1325 : _GEN1320;
wire  _GEN1327 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1328 = io_x[19] ? _GEN1327 : _GEN345;
wire  _GEN1329 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1330 = io_x[19] ? _GEN1329 : _GEN345;
wire  _GEN1331 = io_x[23] ? _GEN1330 : _GEN1328;
wire  _GEN1332 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1333 = io_x[23] ? _GEN370 : _GEN1332;
wire  _GEN1334 = io_x[18] ? _GEN1333 : _GEN1331;
wire  _GEN1335 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1336 = io_x[19] ? _GEN1335 : _GEN345;
wire  _GEN1337 = io_x[23] ? _GEN332 : _GEN1336;
wire  _GEN1338 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1339 = io_x[23] ? _GEN370 : _GEN1338;
wire  _GEN1340 = io_x[18] ? _GEN1339 : _GEN1337;
wire  _GEN1341 = io_x[33] ? _GEN1340 : _GEN1334;
wire  _GEN1342 = io_x[31] ? _GEN1341 : _GEN1326;
wire  _GEN1343 = io_x[28] ? _GEN1342 : _GEN1318;
wire  _GEN1344 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1345 = io_x[19] ? _GEN1344 : _GEN345;
wire  _GEN1346 = io_x[23] ? _GEN1345 : _GEN370;
wire  _GEN1347 = io_x[18] ? _GEN1346 : _GEN362;
wire  _GEN1348 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1349 = io_x[19] ? _GEN1348 : _GEN345;
wire  _GEN1350 = io_x[23] ? _GEN1349 : _GEN332;
wire  _GEN1351 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1352 = io_x[27] ? _GEN1351 : _GEN336;
wire  _GEN1353 = io_x[19] ? _GEN1352 : _GEN345;
wire  _GEN1354 = io_x[23] ? _GEN1353 : _GEN370;
wire  _GEN1355 = io_x[18] ? _GEN1354 : _GEN1350;
wire  _GEN1356 = io_x[33] ? _GEN1355 : _GEN1347;
wire  _GEN1357 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1358 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1359 = io_x[27] ? _GEN1358 : _GEN1357;
wire  _GEN1360 = io_x[19] ? _GEN1359 : _GEN345;
wire  _GEN1361 = io_x[23] ? _GEN1360 : _GEN332;
wire  _GEN1362 = io_x[18] ? _GEN1361 : _GEN331;
wire  _GEN1363 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN1364 = io_x[23] ? _GEN1363 : _GEN332;
wire  _GEN1365 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1366 = io_x[19] ? _GEN345 : _GEN1365;
wire  _GEN1367 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1368 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1369 = io_x[27] ? _GEN1368 : _GEN343;
wire  _GEN1370 = io_x[19] ? _GEN1369 : _GEN1367;
wire  _GEN1371 = io_x[23] ? _GEN1370 : _GEN1366;
wire  _GEN1372 = io_x[18] ? _GEN1371 : _GEN1364;
wire  _GEN1373 = io_x[33] ? _GEN1372 : _GEN1362;
wire  _GEN1374 = io_x[31] ? _GEN1373 : _GEN1356;
wire  _GEN1375 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1376 = io_x[19] ? _GEN1375 : _GEN345;
wire  _GEN1377 = io_x[23] ? _GEN332 : _GEN1376;
wire  _GEN1378 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1379 = io_x[27] ? _GEN343 : _GEN1378;
wire  _GEN1380 = io_x[19] ? _GEN1379 : _GEN345;
wire  _GEN1381 = io_x[23] ? _GEN1380 : _GEN332;
wire  _GEN1382 = io_x[18] ? _GEN1381 : _GEN1377;
wire  _GEN1383 = io_x[18] ? _GEN331 : _GEN362;
wire  _GEN1384 = io_x[33] ? _GEN1383 : _GEN1382;
wire  _GEN1385 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1386 = io_x[23] ? _GEN1385 : _GEN332;
wire  _GEN1387 = io_x[18] ? _GEN1386 : _GEN362;
wire  _GEN1388 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1389 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1390 = io_x[27] ? _GEN343 : _GEN1389;
wire  _GEN1391 = io_x[19] ? _GEN1390 : _GEN345;
wire  _GEN1392 = io_x[23] ? _GEN1391 : _GEN1388;
wire  _GEN1393 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1394 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1395 = io_x[27] ? _GEN1394 : _GEN1393;
wire  _GEN1396 = io_x[19] ? _GEN1395 : _GEN345;
wire  _GEN1397 = io_x[23] ? _GEN1396 : _GEN332;
wire  _GEN1398 = io_x[18] ? _GEN1397 : _GEN1392;
wire  _GEN1399 = io_x[33] ? _GEN1398 : _GEN1387;
wire  _GEN1400 = io_x[31] ? _GEN1399 : _GEN1384;
wire  _GEN1401 = io_x[28] ? _GEN1400 : _GEN1374;
wire  _GEN1402 = io_x[26] ? _GEN1401 : _GEN1343;
wire  _GEN1403 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1404 = io_x[19] ? _GEN1403 : _GEN345;
wire  _GEN1405 = io_x[23] ? _GEN1404 : _GEN332;
wire  _GEN1406 = io_x[18] ? _GEN331 : _GEN1405;
wire  _GEN1407 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1408 = io_x[23] ? _GEN1407 : _GEN332;
wire  _GEN1409 = io_x[18] ? _GEN1408 : _GEN362;
wire  _GEN1410 = io_x[33] ? _GEN1409 : _GEN1406;
wire  _GEN1411 = 1'b0;
wire  _GEN1412 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1413 = io_x[27] ? _GEN1412 : _GEN343;
wire  _GEN1414 = io_x[19] ? _GEN1413 : _GEN338;
wire  _GEN1415 = io_x[23] ? _GEN1414 : _GEN370;
wire  _GEN1416 = io_x[18] ? _GEN1415 : _GEN362;
wire  _GEN1417 = io_x[33] ? _GEN1416 : _GEN1411;
wire  _GEN1418 = io_x[31] ? _GEN1417 : _GEN1410;
wire  _GEN1419 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1420 = io_x[19] ? _GEN345 : _GEN1419;
wire  _GEN1421 = io_x[23] ? _GEN1420 : _GEN332;
wire  _GEN1422 = io_x[18] ? _GEN362 : _GEN1421;
wire  _GEN1423 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1424 = io_x[19] ? _GEN338 : _GEN1423;
wire  _GEN1425 = io_x[23] ? _GEN1424 : _GEN332;
wire  _GEN1426 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN1427 = io_x[18] ? _GEN1426 : _GEN1425;
wire  _GEN1428 = io_x[33] ? _GEN1427 : _GEN1422;
wire  _GEN1429 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1430 = io_x[27] ? _GEN1429 : _GEN336;
wire  _GEN1431 = io_x[19] ? _GEN345 : _GEN1430;
wire  _GEN1432 = io_x[23] ? _GEN1431 : _GEN332;
wire  _GEN1433 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1434 = io_x[19] ? _GEN1433 : _GEN345;
wire  _GEN1435 = io_x[23] ? _GEN1434 : _GEN370;
wire  _GEN1436 = io_x[18] ? _GEN1435 : _GEN1432;
wire  _GEN1437 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1438 = io_x[19] ? _GEN345 : _GEN1437;
wire  _GEN1439 = io_x[23] ? _GEN1438 : _GEN332;
wire  _GEN1440 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1441 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1442 = io_x[27] ? _GEN1441 : _GEN1440;
wire  _GEN1443 = io_x[19] ? _GEN1442 : _GEN345;
wire  _GEN1444 = io_x[23] ? _GEN1443 : _GEN370;
wire  _GEN1445 = io_x[18] ? _GEN1444 : _GEN1439;
wire  _GEN1446 = io_x[33] ? _GEN1445 : _GEN1436;
wire  _GEN1447 = io_x[31] ? _GEN1446 : _GEN1428;
wire  _GEN1448 = io_x[28] ? _GEN1447 : _GEN1418;
wire  _GEN1449 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1450 = io_x[27] ? _GEN336 : _GEN1449;
wire  _GEN1451 = io_x[19] ? _GEN345 : _GEN1450;
wire  _GEN1452 = io_x[23] ? _GEN1451 : _GEN332;
wire  _GEN1453 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1454 = io_x[27] ? _GEN1453 : _GEN336;
wire  _GEN1455 = io_x[19] ? _GEN1454 : _GEN345;
wire  _GEN1456 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1457 = io_x[27] ? _GEN1456 : _GEN343;
wire  _GEN1458 = io_x[19] ? _GEN1457 : _GEN345;
wire  _GEN1459 = io_x[23] ? _GEN1458 : _GEN1455;
wire  _GEN1460 = io_x[18] ? _GEN1459 : _GEN1452;
wire  _GEN1461 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1462 = io_x[27] ? _GEN343 : _GEN1461;
wire  _GEN1463 = io_x[19] ? _GEN1462 : _GEN345;
wire  _GEN1464 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1465 = io_x[27] ? _GEN336 : _GEN1464;
wire  _GEN1466 = io_x[19] ? _GEN345 : _GEN1465;
wire  _GEN1467 = io_x[23] ? _GEN1466 : _GEN1463;
wire  _GEN1468 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1469 = io_x[27] ? _GEN1468 : _GEN343;
wire  _GEN1470 = io_x[19] ? _GEN1469 : _GEN345;
wire  _GEN1471 = io_x[23] ? _GEN332 : _GEN1470;
wire  _GEN1472 = io_x[18] ? _GEN1471 : _GEN1467;
wire  _GEN1473 = io_x[33] ? _GEN1472 : _GEN1460;
wire  _GEN1474 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN1475 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1476 = io_x[27] ? _GEN1475 : _GEN343;
wire  _GEN1477 = io_x[19] ? _GEN1476 : _GEN345;
wire  _GEN1478 = io_x[23] ? _GEN1477 : _GEN332;
wire  _GEN1479 = io_x[18] ? _GEN1478 : _GEN1474;
wire  _GEN1480 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1481 = io_x[19] ? _GEN338 : _GEN1480;
wire  _GEN1482 = io_x[23] ? _GEN1481 : _GEN332;
wire  _GEN1483 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1484 = io_x[27] ? _GEN1483 : _GEN343;
wire  _GEN1485 = io_x[19] ? _GEN1484 : _GEN345;
wire  _GEN1486 = io_x[23] ? _GEN1485 : _GEN332;
wire  _GEN1487 = io_x[18] ? _GEN1486 : _GEN1482;
wire  _GEN1488 = io_x[33] ? _GEN1487 : _GEN1479;
wire  _GEN1489 = io_x[31] ? _GEN1488 : _GEN1473;
wire  _GEN1490 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1491 = io_x[23] ? _GEN1490 : _GEN332;
wire  _GEN1492 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN1493 = io_x[18] ? _GEN1492 : _GEN1491;
wire  _GEN1494 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1495 = io_x[23] ? _GEN1494 : _GEN332;
wire  _GEN1496 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1497 = io_x[27] ? _GEN336 : _GEN1496;
wire  _GEN1498 = io_x[19] ? _GEN1497 : _GEN345;
wire  _GEN1499 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1500 = io_x[19] ? _GEN1499 : _GEN345;
wire  _GEN1501 = io_x[23] ? _GEN1500 : _GEN1498;
wire  _GEN1502 = io_x[18] ? _GEN1501 : _GEN1495;
wire  _GEN1503 = io_x[33] ? _GEN1502 : _GEN1493;
wire  _GEN1504 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN1505 = io_x[23] ? _GEN1504 : _GEN332;
wire  _GEN1506 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1507 = io_x[27] ? _GEN1506 : _GEN336;
wire  _GEN1508 = io_x[19] ? _GEN338 : _GEN1507;
wire  _GEN1509 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1510 = io_x[27] ? _GEN1509 : _GEN343;
wire  _GEN1511 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1512 = io_x[27] ? _GEN1511 : _GEN343;
wire  _GEN1513 = io_x[19] ? _GEN1512 : _GEN1510;
wire  _GEN1514 = io_x[23] ? _GEN1513 : _GEN1508;
wire  _GEN1515 = io_x[18] ? _GEN1514 : _GEN1505;
wire  _GEN1516 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN1517 = io_x[23] ? _GEN1516 : _GEN332;
wire  _GEN1518 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1519 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1520 = io_x[27] ? _GEN1519 : _GEN1518;
wire  _GEN1521 = io_x[19] ? _GEN1520 : _GEN345;
wire  _GEN1522 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1523 = io_x[27] ? _GEN1522 : _GEN343;
wire  _GEN1524 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1525 = io_x[27] ? _GEN1524 : _GEN343;
wire  _GEN1526 = io_x[19] ? _GEN1525 : _GEN1523;
wire  _GEN1527 = io_x[23] ? _GEN1526 : _GEN1521;
wire  _GEN1528 = io_x[18] ? _GEN1527 : _GEN1517;
wire  _GEN1529 = io_x[33] ? _GEN1528 : _GEN1515;
wire  _GEN1530 = io_x[31] ? _GEN1529 : _GEN1503;
wire  _GEN1531 = io_x[28] ? _GEN1530 : _GEN1489;
wire  _GEN1532 = io_x[26] ? _GEN1531 : _GEN1448;
wire  _GEN1533 = io_x[20] ? _GEN1532 : _GEN1402;
wire  _GEN1534 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1535 = io_x[27] ? _GEN1534 : _GEN343;
wire  _GEN1536 = io_x[19] ? _GEN1535 : _GEN338;
wire  _GEN1537 = io_x[23] ? _GEN332 : _GEN1536;
wire  _GEN1538 = io_x[18] ? _GEN1537 : _GEN362;
wire  _GEN1539 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1540 = io_x[19] ? _GEN338 : _GEN1539;
wire  _GEN1541 = io_x[23] ? _GEN332 : _GEN1540;
wire  _GEN1542 = io_x[18] ? _GEN1541 : _GEN331;
wire  _GEN1543 = io_x[33] ? _GEN1542 : _GEN1538;
wire  _GEN1544 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN1545 = io_x[18] ? _GEN1544 : _GEN331;
wire  _GEN1546 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1547 = io_x[27] ? _GEN1546 : _GEN343;
wire  _GEN1548 = io_x[19] ? _GEN1547 : _GEN345;
wire  _GEN1549 = io_x[23] ? _GEN1548 : _GEN370;
wire  _GEN1550 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1551 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1552 = io_x[27] ? _GEN1551 : _GEN343;
wire  _GEN1553 = io_x[19] ? _GEN1552 : _GEN1550;
wire  _GEN1554 = io_x[23] ? _GEN370 : _GEN1553;
wire  _GEN1555 = io_x[18] ? _GEN1554 : _GEN1549;
wire  _GEN1556 = io_x[33] ? _GEN1555 : _GEN1545;
wire  _GEN1557 = io_x[31] ? _GEN1556 : _GEN1543;
wire  _GEN1558 = io_x[18] ? _GEN331 : _GEN362;
wire  _GEN1559 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1560 = io_x[27] ? _GEN1559 : _GEN343;
wire  _GEN1561 = io_x[19] ? _GEN1560 : _GEN338;
wire  _GEN1562 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1563 = io_x[19] ? _GEN1562 : _GEN345;
wire  _GEN1564 = io_x[23] ? _GEN1563 : _GEN1561;
wire  _GEN1565 = io_x[18] ? _GEN1564 : _GEN362;
wire  _GEN1566 = io_x[33] ? _GEN1565 : _GEN1558;
wire  _GEN1567 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1568 = io_x[23] ? _GEN332 : _GEN1567;
wire  _GEN1569 = io_x[18] ? _GEN1568 : _GEN331;
wire  _GEN1570 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1571 = io_x[27] ? _GEN1570 : _GEN343;
wire  _GEN1572 = io_x[19] ? _GEN1571 : _GEN345;
wire  _GEN1573 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1574 = io_x[19] ? _GEN1573 : _GEN345;
wire  _GEN1575 = io_x[23] ? _GEN1574 : _GEN1572;
wire  _GEN1576 = io_x[18] ? _GEN1575 : _GEN362;
wire  _GEN1577 = io_x[33] ? _GEN1576 : _GEN1569;
wire  _GEN1578 = io_x[31] ? _GEN1577 : _GEN1566;
wire  _GEN1579 = io_x[28] ? _GEN1578 : _GEN1557;
wire  _GEN1580 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN1581 = io_x[23] ? _GEN370 : _GEN1580;
wire  _GEN1582 = io_x[18] ? _GEN1581 : _GEN331;
wire  _GEN1583 = io_x[33] ? _GEN1411 : _GEN1582;
wire  _GEN1584 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1585 = io_x[19] ? _GEN1584 : _GEN345;
wire  _GEN1586 = io_x[23] ? _GEN1585 : _GEN332;
wire  _GEN1587 = io_x[18] ? _GEN1586 : _GEN362;
wire  _GEN1588 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1589 = io_x[19] ? _GEN1588 : _GEN345;
wire  _GEN1590 = io_x[23] ? _GEN1589 : _GEN332;
wire  _GEN1591 = io_x[18] ? _GEN1590 : _GEN331;
wire  _GEN1592 = io_x[33] ? _GEN1591 : _GEN1587;
wire  _GEN1593 = io_x[31] ? _GEN1592 : _GEN1583;
wire  _GEN1594 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1595 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1596 = io_x[27] ? _GEN1595 : _GEN343;
wire  _GEN1597 = io_x[19] ? _GEN1596 : _GEN345;
wire  _GEN1598 = io_x[23] ? _GEN1597 : _GEN1594;
wire  _GEN1599 = io_x[18] ? _GEN1598 : _GEN362;
wire  _GEN1600 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1601 = io_x[19] ? _GEN345 : _GEN1600;
wire  _GEN1602 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1603 = io_x[27] ? _GEN1602 : _GEN343;
wire  _GEN1604 = io_x[19] ? _GEN1603 : _GEN345;
wire  _GEN1605 = io_x[23] ? _GEN1604 : _GEN1601;
wire  _GEN1606 = io_x[18] ? _GEN1605 : _GEN362;
wire  _GEN1607 = io_x[33] ? _GEN1606 : _GEN1599;
wire  _GEN1608 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1609 = io_x[27] ? _GEN1608 : _GEN343;
wire  _GEN1610 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1611 = io_x[27] ? _GEN1610 : _GEN343;
wire  _GEN1612 = io_x[19] ? _GEN1611 : _GEN1609;
wire  _GEN1613 = io_x[23] ? _GEN1612 : _GEN370;
wire  _GEN1614 = io_x[18] ? _GEN331 : _GEN1613;
wire  _GEN1615 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1616 = io_x[27] ? _GEN1615 : _GEN343;
wire  _GEN1617 = io_x[19] ? _GEN345 : _GEN1616;
wire  _GEN1618 = io_x[23] ? _GEN1617 : _GEN370;
wire  _GEN1619 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1620 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1621 = io_x[27] ? _GEN1620 : _GEN1619;
wire  _GEN1622 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1623 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1624 = io_x[27] ? _GEN1623 : _GEN1622;
wire  _GEN1625 = io_x[19] ? _GEN1624 : _GEN1621;
wire  _GEN1626 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1627 = io_x[27] ? _GEN1626 : _GEN343;
wire  _GEN1628 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1629 = io_x[27] ? _GEN1628 : _GEN343;
wire  _GEN1630 = io_x[19] ? _GEN1629 : _GEN1627;
wire  _GEN1631 = io_x[23] ? _GEN1630 : _GEN1625;
wire  _GEN1632 = io_x[18] ? _GEN1631 : _GEN1618;
wire  _GEN1633 = io_x[33] ? _GEN1632 : _GEN1614;
wire  _GEN1634 = io_x[31] ? _GEN1633 : _GEN1607;
wire  _GEN1635 = io_x[28] ? _GEN1634 : _GEN1593;
wire  _GEN1636 = io_x[26] ? _GEN1635 : _GEN1579;
wire  _GEN1637 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1638 = io_x[19] ? _GEN345 : _GEN1637;
wire  _GEN1639 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1640 = io_x[23] ? _GEN1639 : _GEN1638;
wire  _GEN1641 = io_x[18] ? _GEN362 : _GEN1640;
wire  _GEN1642 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1643 = io_x[19] ? _GEN345 : _GEN1642;
wire  _GEN1644 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1645 = io_x[23] ? _GEN1644 : _GEN1643;
wire  _GEN1646 = io_x[18] ? _GEN331 : _GEN1645;
wire  _GEN1647 = io_x[33] ? _GEN1646 : _GEN1641;
wire  _GEN1648 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1649 = io_x[23] ? _GEN332 : _GEN1648;
wire  _GEN1650 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1651 = io_x[27] ? _GEN1650 : _GEN343;
wire  _GEN1652 = io_x[19] ? _GEN1651 : _GEN345;
wire  _GEN1653 = io_x[23] ? _GEN1652 : _GEN332;
wire  _GEN1654 = io_x[18] ? _GEN1653 : _GEN1649;
wire  _GEN1655 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1656 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1657 = io_x[27] ? _GEN1656 : _GEN343;
wire  _GEN1658 = io_x[19] ? _GEN1657 : _GEN345;
wire  _GEN1659 = io_x[23] ? _GEN1658 : _GEN1655;
wire  _GEN1660 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1661 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1662 = io_x[27] ? _GEN1661 : _GEN1660;
wire  _GEN1663 = io_x[19] ? _GEN1662 : _GEN338;
wire  _GEN1664 = io_x[23] ? _GEN1663 : _GEN332;
wire  _GEN1665 = io_x[18] ? _GEN1664 : _GEN1659;
wire  _GEN1666 = io_x[33] ? _GEN1665 : _GEN1654;
wire  _GEN1667 = io_x[31] ? _GEN1666 : _GEN1647;
wire  _GEN1668 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1669 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1670 = io_x[27] ? _GEN336 : _GEN1669;
wire  _GEN1671 = io_x[19] ? _GEN1670 : _GEN1668;
wire  _GEN1672 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1673 = io_x[23] ? _GEN1672 : _GEN1671;
wire  _GEN1674 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1675 = io_x[19] ? _GEN1674 : _GEN338;
wire  _GEN1676 = io_x[23] ? _GEN1675 : _GEN370;
wire  _GEN1677 = io_x[18] ? _GEN1676 : _GEN1673;
wire  _GEN1678 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1679 = io_x[27] ? _GEN343 : _GEN1678;
wire  _GEN1680 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1681 = io_x[19] ? _GEN1680 : _GEN1679;
wire  _GEN1682 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1683 = io_x[27] ? _GEN1682 : _GEN336;
wire  _GEN1684 = io_x[19] ? _GEN1683 : _GEN338;
wire  _GEN1685 = io_x[23] ? _GEN1684 : _GEN1681;
wire  _GEN1686 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1687 = io_x[27] ? _GEN1686 : _GEN343;
wire  _GEN1688 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1689 = io_x[27] ? _GEN1688 : _GEN343;
wire  _GEN1690 = io_x[19] ? _GEN1689 : _GEN1687;
wire  _GEN1691 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1692 = io_x[23] ? _GEN1691 : _GEN1690;
wire  _GEN1693 = io_x[18] ? _GEN1692 : _GEN1685;
wire  _GEN1694 = io_x[33] ? _GEN1693 : _GEN1677;
wire  _GEN1695 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1696 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1697 = io_x[27] ? _GEN1696 : _GEN343;
wire  _GEN1698 = io_x[19] ? _GEN1697 : _GEN345;
wire  _GEN1699 = io_x[23] ? _GEN1698 : _GEN1695;
wire  _GEN1700 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1701 = io_x[27] ? _GEN343 : _GEN1700;
wire  _GEN1702 = io_x[19] ? _GEN1701 : _GEN338;
wire  _GEN1703 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1704 = io_x[27] ? _GEN1703 : _GEN343;
wire  _GEN1705 = io_x[19] ? _GEN1704 : _GEN345;
wire  _GEN1706 = io_x[23] ? _GEN1705 : _GEN1702;
wire  _GEN1707 = io_x[18] ? _GEN1706 : _GEN1699;
wire  _GEN1708 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1709 = io_x[19] ? _GEN1708 : _GEN338;
wire  _GEN1710 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1711 = io_x[27] ? _GEN1710 : _GEN343;
wire  _GEN1712 = io_x[19] ? _GEN1711 : _GEN345;
wire  _GEN1713 = io_x[23] ? _GEN1712 : _GEN1709;
wire  _GEN1714 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1715 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1716 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1717 = io_x[27] ? _GEN1716 : _GEN1715;
wire  _GEN1718 = io_x[19] ? _GEN1717 : _GEN345;
wire  _GEN1719 = io_x[23] ? _GEN1718 : _GEN1714;
wire  _GEN1720 = io_x[18] ? _GEN1719 : _GEN1713;
wire  _GEN1721 = io_x[33] ? _GEN1720 : _GEN1707;
wire  _GEN1722 = io_x[31] ? _GEN1721 : _GEN1694;
wire  _GEN1723 = io_x[28] ? _GEN1722 : _GEN1667;
wire  _GEN1724 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1725 = io_x[27] ? _GEN1724 : _GEN343;
wire  _GEN1726 = io_x[19] ? _GEN1725 : _GEN345;
wire  _GEN1727 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1728 = io_x[19] ? _GEN1727 : _GEN345;
wire  _GEN1729 = io_x[23] ? _GEN1728 : _GEN1726;
wire  _GEN1730 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1731 = io_x[27] ? _GEN343 : _GEN1730;
wire  _GEN1732 = io_x[19] ? _GEN1731 : _GEN345;
wire  _GEN1733 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1734 = io_x[27] ? _GEN1733 : _GEN343;
wire  _GEN1735 = io_x[19] ? _GEN1734 : _GEN345;
wire  _GEN1736 = io_x[23] ? _GEN1735 : _GEN1732;
wire  _GEN1737 = io_x[18] ? _GEN1736 : _GEN1729;
wire  _GEN1738 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1739 = io_x[19] ? _GEN338 : _GEN1738;
wire  _GEN1740 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1741 = io_x[27] ? _GEN1740 : _GEN343;
wire  _GEN1742 = io_x[19] ? _GEN1741 : _GEN345;
wire  _GEN1743 = io_x[23] ? _GEN1742 : _GEN1739;
wire  _GEN1744 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1745 = io_x[27] ? _GEN336 : _GEN1744;
wire  _GEN1746 = io_x[19] ? _GEN1745 : _GEN345;
wire  _GEN1747 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1748 = io_x[27] ? _GEN1747 : _GEN343;
wire  _GEN1749 = io_x[19] ? _GEN1748 : _GEN345;
wire  _GEN1750 = io_x[23] ? _GEN1749 : _GEN1746;
wire  _GEN1751 = io_x[18] ? _GEN1750 : _GEN1743;
wire  _GEN1752 = io_x[33] ? _GEN1751 : _GEN1737;
wire  _GEN1753 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1754 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1755 = io_x[27] ? _GEN1754 : _GEN343;
wire  _GEN1756 = io_x[19] ? _GEN1755 : _GEN1753;
wire  _GEN1757 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1758 = io_x[27] ? _GEN1757 : _GEN343;
wire  _GEN1759 = io_x[19] ? _GEN1758 : _GEN345;
wire  _GEN1760 = io_x[23] ? _GEN1759 : _GEN1756;
wire  _GEN1761 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1762 = io_x[27] ? _GEN1761 : _GEN343;
wire  _GEN1763 = io_x[19] ? _GEN338 : _GEN1762;
wire  _GEN1764 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1765 = io_x[27] ? _GEN1764 : _GEN343;
wire  _GEN1766 = io_x[19] ? _GEN1765 : _GEN338;
wire  _GEN1767 = io_x[23] ? _GEN1766 : _GEN1763;
wire  _GEN1768 = io_x[18] ? _GEN1767 : _GEN1760;
wire  _GEN1769 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1770 = io_x[27] ? _GEN1769 : _GEN343;
wire  _GEN1771 = io_x[19] ? _GEN1770 : _GEN338;
wire  _GEN1772 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1773 = io_x[27] ? _GEN1772 : _GEN343;
wire  _GEN1774 = io_x[19] ? _GEN1773 : _GEN345;
wire  _GEN1775 = io_x[23] ? _GEN1774 : _GEN1771;
wire  _GEN1776 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN1777 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1778 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1779 = io_x[27] ? _GEN1778 : _GEN1777;
wire  _GEN1780 = io_x[19] ? _GEN1779 : _GEN345;
wire  _GEN1781 = io_x[23] ? _GEN1780 : _GEN1776;
wire  _GEN1782 = io_x[18] ? _GEN1781 : _GEN1775;
wire  _GEN1783 = io_x[33] ? _GEN1782 : _GEN1768;
wire  _GEN1784 = io_x[31] ? _GEN1783 : _GEN1752;
wire  _GEN1785 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1786 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1787 = io_x[27] ? _GEN336 : _GEN1786;
wire  _GEN1788 = io_x[19] ? _GEN1787 : _GEN1785;
wire  _GEN1789 = io_x[23] ? _GEN1788 : _GEN370;
wire  _GEN1790 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1791 = io_x[27] ? _GEN343 : _GEN1790;
wire  _GEN1792 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1793 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1794 = io_x[27] ? _GEN1793 : _GEN1792;
wire  _GEN1795 = io_x[19] ? _GEN1794 : _GEN1791;
wire  _GEN1796 = io_x[23] ? _GEN1795 : _GEN332;
wire  _GEN1797 = io_x[18] ? _GEN1796 : _GEN1789;
wire  _GEN1798 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1799 = io_x[19] ? _GEN338 : _GEN1798;
wire  _GEN1800 = io_x[23] ? _GEN370 : _GEN1799;
wire  _GEN1801 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1802 = io_x[27] ? _GEN343 : _GEN1801;
wire  _GEN1803 = io_x[19] ? _GEN1802 : _GEN345;
wire  _GEN1804 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1805 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1806 = io_x[27] ? _GEN1805 : _GEN1804;
wire  _GEN1807 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1808 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1809 = io_x[27] ? _GEN1808 : _GEN1807;
wire  _GEN1810 = io_x[19] ? _GEN1809 : _GEN1806;
wire  _GEN1811 = io_x[23] ? _GEN1810 : _GEN1803;
wire  _GEN1812 = io_x[18] ? _GEN1811 : _GEN1800;
wire  _GEN1813 = io_x[33] ? _GEN1812 : _GEN1797;
wire  _GEN1814 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1815 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1816 = io_x[19] ? _GEN1815 : _GEN1814;
wire  _GEN1817 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1818 = io_x[27] ? _GEN1817 : _GEN336;
wire  _GEN1819 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1820 = io_x[27] ? _GEN1819 : _GEN343;
wire  _GEN1821 = io_x[19] ? _GEN1820 : _GEN1818;
wire  _GEN1822 = io_x[23] ? _GEN1821 : _GEN1816;
wire  _GEN1823 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1824 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1825 = io_x[27] ? _GEN1824 : _GEN1823;
wire  _GEN1826 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1827 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1828 = io_x[27] ? _GEN1827 : _GEN1826;
wire  _GEN1829 = io_x[19] ? _GEN1828 : _GEN1825;
wire  _GEN1830 = io_x[23] ? _GEN1829 : _GEN370;
wire  _GEN1831 = io_x[18] ? _GEN1830 : _GEN1822;
wire  _GEN1832 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1833 = io_x[27] ? _GEN1832 : _GEN343;
wire  _GEN1834 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1835 = io_x[19] ? _GEN1834 : _GEN1833;
wire  _GEN1836 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1837 = io_x[27] ? _GEN1836 : _GEN336;
wire  _GEN1838 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1839 = io_x[27] ? _GEN1838 : _GEN343;
wire  _GEN1840 = io_x[19] ? _GEN1839 : _GEN1837;
wire  _GEN1841 = io_x[23] ? _GEN1840 : _GEN1835;
wire  _GEN1842 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1843 = io_x[27] ? _GEN1842 : _GEN336;
wire  _GEN1844 = io_x[19] ? _GEN1843 : _GEN338;
wire  _GEN1845 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1846 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1847 = io_x[27] ? _GEN1846 : _GEN1845;
wire  _GEN1848 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1849 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1850 = io_x[27] ? _GEN1849 : _GEN1848;
wire  _GEN1851 = io_x[19] ? _GEN1850 : _GEN1847;
wire  _GEN1852 = io_x[23] ? _GEN1851 : _GEN1844;
wire  _GEN1853 = io_x[18] ? _GEN1852 : _GEN1841;
wire  _GEN1854 = io_x[33] ? _GEN1853 : _GEN1831;
wire  _GEN1855 = io_x[31] ? _GEN1854 : _GEN1813;
wire  _GEN1856 = io_x[28] ? _GEN1855 : _GEN1784;
wire  _GEN1857 = io_x[26] ? _GEN1856 : _GEN1723;
wire  _GEN1858 = io_x[20] ? _GEN1857 : _GEN1636;
wire  _GEN1859 = io_x[24] ? _GEN1858 : _GEN1533;
wire  _GEN1860 = io_x[78] ? _GEN1859 : _GEN1295;
wire  _GEN1861 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1862 = io_x[23] ? _GEN1861 : _GEN370;
wire  _GEN1863 = io_x[18] ? _GEN362 : _GEN1862;
wire  _GEN1864 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1865 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1866 = io_x[27] ? _GEN1865 : _GEN1864;
wire  _GEN1867 = io_x[19] ? _GEN1866 : _GEN338;
wire  _GEN1868 = io_x[23] ? _GEN1867 : _GEN332;
wire  _GEN1869 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1870 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1871 = io_x[27] ? _GEN1870 : _GEN1869;
wire  _GEN1872 = io_x[19] ? _GEN1871 : _GEN338;
wire  _GEN1873 = io_x[23] ? _GEN1872 : _GEN332;
wire  _GEN1874 = io_x[18] ? _GEN1873 : _GEN1868;
wire  _GEN1875 = io_x[33] ? _GEN1874 : _GEN1863;
wire  _GEN1876 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1877 = io_x[27] ? _GEN1876 : _GEN343;
wire  _GEN1878 = io_x[19] ? _GEN1877 : _GEN345;
wire  _GEN1879 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1880 = io_x[19] ? _GEN1879 : _GEN345;
wire  _GEN1881 = io_x[23] ? _GEN1880 : _GEN1878;
wire  _GEN1882 = io_x[18] ? _GEN362 : _GEN1881;
wire  _GEN1883 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN1884 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1885 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1886 = io_x[27] ? _GEN1885 : _GEN1884;
wire  _GEN1887 = io_x[19] ? _GEN1886 : _GEN345;
wire  _GEN1888 = io_x[23] ? _GEN1887 : _GEN1883;
wire  _GEN1889 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1890 = io_x[27] ? _GEN1889 : _GEN343;
wire  _GEN1891 = io_x[19] ? _GEN1890 : _GEN345;
wire  _GEN1892 = io_x[23] ? _GEN1891 : _GEN370;
wire  _GEN1893 = io_x[18] ? _GEN1892 : _GEN1888;
wire  _GEN1894 = io_x[33] ? _GEN1893 : _GEN1882;
wire  _GEN1895 = io_x[31] ? _GEN1894 : _GEN1875;
wire  _GEN1896 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN1897 = io_x[18] ? _GEN362 : _GEN1896;
wire  _GEN1898 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1899 = io_x[19] ? _GEN1898 : _GEN345;
wire  _GEN1900 = io_x[23] ? _GEN370 : _GEN1899;
wire  _GEN1901 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1902 = io_x[27] ? _GEN1901 : _GEN343;
wire  _GEN1903 = io_x[19] ? _GEN1902 : _GEN338;
wire  _GEN1904 = io_x[23] ? _GEN370 : _GEN1903;
wire  _GEN1905 = io_x[18] ? _GEN1904 : _GEN1900;
wire  _GEN1906 = io_x[33] ? _GEN1905 : _GEN1897;
wire  _GEN1907 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1908 = io_x[19] ? _GEN1907 : _GEN345;
wire  _GEN1909 = io_x[23] ? _GEN332 : _GEN1908;
wire  _GEN1910 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1911 = io_x[19] ? _GEN1910 : _GEN345;
wire  _GEN1912 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1913 = io_x[27] ? _GEN1912 : _GEN343;
wire  _GEN1914 = io_x[19] ? _GEN1913 : _GEN338;
wire  _GEN1915 = io_x[23] ? _GEN1914 : _GEN1911;
wire  _GEN1916 = io_x[18] ? _GEN1915 : _GEN1909;
wire  _GEN1917 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1918 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1919 = io_x[27] ? _GEN1918 : _GEN1917;
wire  _GEN1920 = io_x[19] ? _GEN1919 : _GEN338;
wire  _GEN1921 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1922 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1923 = io_x[27] ? _GEN1922 : _GEN1921;
wire  _GEN1924 = io_x[19] ? _GEN1923 : _GEN345;
wire  _GEN1925 = io_x[23] ? _GEN1924 : _GEN1920;
wire  _GEN1926 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1927 = io_x[27] ? _GEN1926 : _GEN336;
wire  _GEN1928 = io_x[19] ? _GEN1927 : _GEN345;
wire  _GEN1929 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1930 = io_x[27] ? _GEN1929 : _GEN343;
wire  _GEN1931 = io_x[19] ? _GEN1930 : _GEN345;
wire  _GEN1932 = io_x[23] ? _GEN1931 : _GEN1928;
wire  _GEN1933 = io_x[18] ? _GEN1932 : _GEN1925;
wire  _GEN1934 = io_x[33] ? _GEN1933 : _GEN1916;
wire  _GEN1935 = io_x[31] ? _GEN1934 : _GEN1906;
wire  _GEN1936 = io_x[28] ? _GEN1935 : _GEN1895;
wire  _GEN1937 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1938 = io_x[27] ? _GEN1937 : _GEN343;
wire  _GEN1939 = io_x[19] ? _GEN1938 : _GEN345;
wire  _GEN1940 = io_x[23] ? _GEN1939 : _GEN332;
wire  _GEN1941 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN1942 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN1943 = io_x[23] ? _GEN1942 : _GEN1941;
wire  _GEN1944 = io_x[18] ? _GEN1943 : _GEN1940;
wire  _GEN1945 = io_x[33] ? _GEN1944 : _GEN1411;
wire  _GEN1946 = io_x[18] ? _GEN331 : _GEN362;
wire  _GEN1947 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1948 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1949 = io_x[27] ? _GEN1948 : _GEN336;
wire  _GEN1950 = io_x[19] ? _GEN1949 : _GEN1947;
wire  _GEN1951 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1952 = io_x[27] ? _GEN1951 : _GEN343;
wire  _GEN1953 = io_x[19] ? _GEN1952 : _GEN345;
wire  _GEN1954 = io_x[23] ? _GEN1953 : _GEN1950;
wire  _GEN1955 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1956 = io_x[27] ? _GEN1955 : _GEN336;
wire  _GEN1957 = io_x[19] ? _GEN1956 : _GEN345;
wire  _GEN1958 = io_x[23] ? _GEN1957 : _GEN370;
wire  _GEN1959 = io_x[18] ? _GEN1958 : _GEN1954;
wire  _GEN1960 = io_x[33] ? _GEN1959 : _GEN1946;
wire  _GEN1961 = io_x[31] ? _GEN1960 : _GEN1945;
wire  _GEN1962 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1963 = io_x[27] ? _GEN343 : _GEN1962;
wire  _GEN1964 = io_x[19] ? _GEN1963 : _GEN338;
wire  _GEN1965 = io_x[23] ? _GEN332 : _GEN1964;
wire  _GEN1966 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN1967 = io_x[19] ? _GEN1966 : _GEN345;
wire  _GEN1968 = io_x[23] ? _GEN1967 : _GEN370;
wire  _GEN1969 = io_x[18] ? _GEN1968 : _GEN1965;
wire  _GEN1970 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN1971 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1972 = io_x[27] ? _GEN343 : _GEN1971;
wire  _GEN1973 = io_x[19] ? _GEN1972 : _GEN345;
wire  _GEN1974 = io_x[23] ? _GEN1973 : _GEN1970;
wire  _GEN1975 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1976 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1977 = io_x[27] ? _GEN1976 : _GEN1975;
wire  _GEN1978 = io_x[19] ? _GEN1977 : _GEN338;
wire  _GEN1979 = io_x[23] ? _GEN1978 : _GEN332;
wire  _GEN1980 = io_x[18] ? _GEN1979 : _GEN1974;
wire  _GEN1981 = io_x[33] ? _GEN1980 : _GEN1969;
wire  _GEN1982 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN1983 = io_x[18] ? _GEN331 : _GEN1982;
wire  _GEN1984 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN1985 = io_x[27] ? _GEN336 : _GEN1984;
wire  _GEN1986 = io_x[19] ? _GEN1985 : _GEN345;
wire  _GEN1987 = io_x[23] ? _GEN1986 : _GEN332;
wire  _GEN1988 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN1989 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN1990 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN1991 = io_x[27] ? _GEN1990 : _GEN336;
wire  _GEN1992 = io_x[19] ? _GEN1991 : _GEN1989;
wire  _GEN1993 = io_x[23] ? _GEN1992 : _GEN1988;
wire  _GEN1994 = io_x[18] ? _GEN1993 : _GEN1987;
wire  _GEN1995 = io_x[33] ? _GEN1994 : _GEN1983;
wire  _GEN1996 = io_x[31] ? _GEN1995 : _GEN1981;
wire  _GEN1997 = io_x[28] ? _GEN1996 : _GEN1961;
wire  _GEN1998 = io_x[26] ? _GEN1997 : _GEN1936;
wire  _GEN1999 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2000 = io_x[27] ? _GEN1999 : _GEN343;
wire  _GEN2001 = io_x[19] ? _GEN2000 : _GEN338;
wire  _GEN2002 = io_x[23] ? _GEN2001 : _GEN370;
wire  _GEN2003 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2004 = io_x[23] ? _GEN2003 : _GEN332;
wire  _GEN2005 = io_x[18] ? _GEN2004 : _GEN2002;
wire  _GEN2006 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2007 = io_x[27] ? _GEN2006 : _GEN343;
wire  _GEN2008 = io_x[19] ? _GEN2007 : _GEN345;
wire  _GEN2009 = io_x[23] ? _GEN2008 : _GEN370;
wire  _GEN2010 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2011 = io_x[27] ? _GEN2010 : _GEN336;
wire  _GEN2012 = io_x[19] ? _GEN2011 : _GEN338;
wire  _GEN2013 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2014 = io_x[27] ? _GEN343 : _GEN2013;
wire  _GEN2015 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2016 = io_x[27] ? _GEN2015 : _GEN343;
wire  _GEN2017 = io_x[19] ? _GEN2016 : _GEN2014;
wire  _GEN2018 = io_x[23] ? _GEN2017 : _GEN2012;
wire  _GEN2019 = io_x[18] ? _GEN2018 : _GEN2009;
wire  _GEN2020 = io_x[33] ? _GEN2019 : _GEN2005;
wire  _GEN2021 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2022 = io_x[27] ? _GEN2021 : _GEN343;
wire  _GEN2023 = io_x[19] ? _GEN2022 : _GEN338;
wire  _GEN2024 = io_x[23] ? _GEN2023 : _GEN332;
wire  _GEN2025 = io_x[18] ? _GEN331 : _GEN2024;
wire  _GEN2026 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2027 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2028 = io_x[27] ? _GEN2027 : _GEN343;
wire  _GEN2029 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2030 = io_x[27] ? _GEN2029 : _GEN343;
wire  _GEN2031 = io_x[19] ? _GEN2030 : _GEN2028;
wire  _GEN2032 = io_x[23] ? _GEN2031 : _GEN2026;
wire  _GEN2033 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2034 = io_x[27] ? _GEN343 : _GEN2033;
wire  _GEN2035 = io_x[19] ? _GEN2034 : _GEN338;
wire  _GEN2036 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2037 = io_x[27] ? _GEN2036 : _GEN343;
wire  _GEN2038 = io_x[19] ? _GEN2037 : _GEN338;
wire  _GEN2039 = io_x[23] ? _GEN2038 : _GEN2035;
wire  _GEN2040 = io_x[18] ? _GEN2039 : _GEN2032;
wire  _GEN2041 = io_x[33] ? _GEN2040 : _GEN2025;
wire  _GEN2042 = io_x[31] ? _GEN2041 : _GEN2020;
wire  _GEN2043 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN2044 = io_x[18] ? _GEN2043 : _GEN331;
wire  _GEN2045 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2046 = io_x[19] ? _GEN2045 : _GEN345;
wire  _GEN2047 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2048 = io_x[23] ? _GEN2047 : _GEN2046;
wire  _GEN2049 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2050 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2051 = io_x[27] ? _GEN2050 : _GEN2049;
wire  _GEN2052 = io_x[19] ? _GEN2051 : _GEN345;
wire  _GEN2053 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2054 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2055 = io_x[27] ? _GEN2054 : _GEN2053;
wire  _GEN2056 = io_x[19] ? _GEN2055 : _GEN345;
wire  _GEN2057 = io_x[23] ? _GEN2056 : _GEN2052;
wire  _GEN2058 = io_x[18] ? _GEN2057 : _GEN2048;
wire  _GEN2059 = io_x[33] ? _GEN2058 : _GEN2044;
wire  _GEN2060 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2061 = io_x[19] ? _GEN338 : _GEN2060;
wire  _GEN2062 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2063 = io_x[27] ? _GEN2062 : _GEN343;
wire  _GEN2064 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2065 = io_x[19] ? _GEN2064 : _GEN2063;
wire  _GEN2066 = io_x[23] ? _GEN2065 : _GEN2061;
wire  _GEN2067 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2068 = io_x[27] ? _GEN2067 : _GEN343;
wire  _GEN2069 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2070 = io_x[27] ? _GEN343 : _GEN2069;
wire  _GEN2071 = io_x[19] ? _GEN2070 : _GEN2068;
wire  _GEN2072 = io_x[23] ? _GEN2071 : _GEN370;
wire  _GEN2073 = io_x[18] ? _GEN2072 : _GEN2066;
wire  _GEN2074 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2075 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2076 = io_x[27] ? _GEN343 : _GEN2075;
wire  _GEN2077 = io_x[19] ? _GEN2076 : _GEN2074;
wire  _GEN2078 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2079 = io_x[27] ? _GEN2078 : _GEN343;
wire  _GEN2080 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2081 = io_x[27] ? _GEN2080 : _GEN343;
wire  _GEN2082 = io_x[19] ? _GEN2081 : _GEN2079;
wire  _GEN2083 = io_x[23] ? _GEN2082 : _GEN2077;
wire  _GEN2084 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2085 = io_x[19] ? _GEN2084 : _GEN338;
wire  _GEN2086 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2087 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2088 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2089 = io_x[27] ? _GEN2088 : _GEN2087;
wire  _GEN2090 = io_x[19] ? _GEN2089 : _GEN2086;
wire  _GEN2091 = io_x[23] ? _GEN2090 : _GEN2085;
wire  _GEN2092 = io_x[18] ? _GEN2091 : _GEN2083;
wire  _GEN2093 = io_x[33] ? _GEN2092 : _GEN2073;
wire  _GEN2094 = io_x[31] ? _GEN2093 : _GEN2059;
wire  _GEN2095 = io_x[28] ? _GEN2094 : _GEN2042;
wire  _GEN2096 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2097 = io_x[27] ? _GEN2096 : _GEN336;
wire  _GEN2098 = io_x[19] ? _GEN345 : _GEN2097;
wire  _GEN2099 = io_x[23] ? _GEN2098 : _GEN370;
wire  _GEN2100 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2101 = io_x[27] ? _GEN336 : _GEN2100;
wire  _GEN2102 = io_x[19] ? _GEN2101 : _GEN338;
wire  _GEN2103 = io_x[23] ? _GEN2102 : _GEN332;
wire  _GEN2104 = io_x[18] ? _GEN2103 : _GEN2099;
wire  _GEN2105 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2106 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2107 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2108 = io_x[27] ? _GEN2107 : _GEN2106;
wire  _GEN2109 = io_x[19] ? _GEN2108 : _GEN2105;
wire  _GEN2110 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2111 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2112 = io_x[27] ? _GEN2111 : _GEN2110;
wire  _GEN2113 = io_x[19] ? _GEN345 : _GEN2112;
wire  _GEN2114 = io_x[23] ? _GEN2113 : _GEN2109;
wire  _GEN2115 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2116 = io_x[19] ? _GEN2115 : _GEN345;
wire  _GEN2117 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2118 = io_x[19] ? _GEN2117 : _GEN338;
wire  _GEN2119 = io_x[23] ? _GEN2118 : _GEN2116;
wire  _GEN2120 = io_x[18] ? _GEN2119 : _GEN2114;
wire  _GEN2121 = io_x[33] ? _GEN2120 : _GEN2104;
wire  _GEN2122 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2123 = io_x[19] ? _GEN345 : _GEN2122;
wire  _GEN2124 = io_x[23] ? _GEN332 : _GEN2123;
wire  _GEN2125 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2126 = io_x[27] ? _GEN2125 : _GEN343;
wire  _GEN2127 = io_x[19] ? _GEN345 : _GEN2126;
wire  _GEN2128 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2129 = io_x[27] ? _GEN2128 : _GEN343;
wire  _GEN2130 = io_x[19] ? _GEN2129 : _GEN345;
wire  _GEN2131 = io_x[23] ? _GEN2130 : _GEN2127;
wire  _GEN2132 = io_x[18] ? _GEN2131 : _GEN2124;
wire  _GEN2133 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2134 = io_x[19] ? _GEN345 : _GEN2133;
wire  _GEN2135 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2136 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2137 = io_x[27] ? _GEN2136 : _GEN2135;
wire  _GEN2138 = io_x[19] ? _GEN2137 : _GEN345;
wire  _GEN2139 = io_x[23] ? _GEN2138 : _GEN2134;
wire  _GEN2140 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2141 = io_x[27] ? _GEN2140 : _GEN343;
wire  _GEN2142 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2143 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2144 = io_x[27] ? _GEN2143 : _GEN2142;
wire  _GEN2145 = io_x[19] ? _GEN2144 : _GEN2141;
wire  _GEN2146 = io_x[23] ? _GEN2145 : _GEN332;
wire  _GEN2147 = io_x[18] ? _GEN2146 : _GEN2139;
wire  _GEN2148 = io_x[33] ? _GEN2147 : _GEN2132;
wire  _GEN2149 = io_x[31] ? _GEN2148 : _GEN2121;
wire  _GEN2150 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2151 = io_x[27] ? _GEN343 : _GEN2150;
wire  _GEN2152 = io_x[19] ? _GEN2151 : _GEN338;
wire  _GEN2153 = io_x[23] ? _GEN2152 : _GEN332;
wire  _GEN2154 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2155 = io_x[27] ? _GEN343 : _GEN2154;
wire  _GEN2156 = io_x[19] ? _GEN345 : _GEN2155;
wire  _GEN2157 = io_x[23] ? _GEN370 : _GEN2156;
wire  _GEN2158 = io_x[18] ? _GEN2157 : _GEN2153;
wire  _GEN2159 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2160 = io_x[19] ? _GEN2159 : _GEN345;
wire  _GEN2161 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2162 = io_x[27] ? _GEN2161 : _GEN336;
wire  _GEN2163 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2164 = io_x[27] ? _GEN343 : _GEN2163;
wire  _GEN2165 = io_x[19] ? _GEN2164 : _GEN2162;
wire  _GEN2166 = io_x[23] ? _GEN2165 : _GEN2160;
wire  _GEN2167 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2168 = io_x[27] ? _GEN343 : _GEN2167;
wire  _GEN2169 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2170 = io_x[27] ? _GEN343 : _GEN2169;
wire  _GEN2171 = io_x[19] ? _GEN2170 : _GEN2168;
wire  _GEN2172 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2173 = io_x[27] ? _GEN2172 : _GEN336;
wire  _GEN2174 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2175 = io_x[27] ? _GEN343 : _GEN2174;
wire  _GEN2176 = io_x[19] ? _GEN2175 : _GEN2173;
wire  _GEN2177 = io_x[23] ? _GEN2176 : _GEN2171;
wire  _GEN2178 = io_x[18] ? _GEN2177 : _GEN2166;
wire  _GEN2179 = io_x[33] ? _GEN2178 : _GEN2158;
wire  _GEN2180 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2181 = io_x[27] ? _GEN2180 : _GEN343;
wire  _GEN2182 = io_x[19] ? _GEN2181 : _GEN338;
wire  _GEN2183 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2184 = io_x[23] ? _GEN2183 : _GEN2182;
wire  _GEN2185 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2186 = io_x[27] ? _GEN2185 : _GEN343;
wire  _GEN2187 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2188 = io_x[27] ? _GEN2187 : _GEN343;
wire  _GEN2189 = io_x[19] ? _GEN2188 : _GEN2186;
wire  _GEN2190 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2191 = io_x[27] ? _GEN2190 : _GEN343;
wire  _GEN2192 = io_x[19] ? _GEN2191 : _GEN345;
wire  _GEN2193 = io_x[23] ? _GEN2192 : _GEN2189;
wire  _GEN2194 = io_x[18] ? _GEN2193 : _GEN2184;
wire  _GEN2195 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2196 = io_x[27] ? _GEN2195 : _GEN343;
wire  _GEN2197 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2198 = io_x[27] ? _GEN336 : _GEN2197;
wire  _GEN2199 = io_x[19] ? _GEN2198 : _GEN2196;
wire  _GEN2200 = io_x[23] ? _GEN2199 : _GEN370;
wire  _GEN2201 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2202 = io_x[27] ? _GEN2201 : _GEN343;
wire  _GEN2203 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2204 = io_x[27] ? _GEN2203 : _GEN336;
wire  _GEN2205 = io_x[19] ? _GEN2204 : _GEN2202;
wire  _GEN2206 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2207 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2208 = io_x[27] ? _GEN2207 : _GEN2206;
wire  _GEN2209 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2210 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2211 = io_x[27] ? _GEN2210 : _GEN2209;
wire  _GEN2212 = io_x[19] ? _GEN2211 : _GEN2208;
wire  _GEN2213 = io_x[23] ? _GEN2212 : _GEN2205;
wire  _GEN2214 = io_x[18] ? _GEN2213 : _GEN2200;
wire  _GEN2215 = io_x[33] ? _GEN2214 : _GEN2194;
wire  _GEN2216 = io_x[31] ? _GEN2215 : _GEN2179;
wire  _GEN2217 = io_x[28] ? _GEN2216 : _GEN2149;
wire  _GEN2218 = io_x[26] ? _GEN2217 : _GEN2095;
wire  _GEN2219 = io_x[20] ? _GEN2218 : _GEN1998;
wire  _GEN2220 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN2221 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2222 = io_x[27] ? _GEN2221 : _GEN343;
wire  _GEN2223 = io_x[19] ? _GEN2222 : _GEN345;
wire  _GEN2224 = io_x[23] ? _GEN2223 : _GEN370;
wire  _GEN2225 = io_x[18] ? _GEN2224 : _GEN2220;
wire  _GEN2226 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2227 = io_x[27] ? _GEN2226 : _GEN343;
wire  _GEN2228 = io_x[19] ? _GEN2227 : _GEN345;
wire  _GEN2229 = io_x[23] ? _GEN2228 : _GEN332;
wire  _GEN2230 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2231 = io_x[19] ? _GEN2230 : _GEN338;
wire  _GEN2232 = io_x[23] ? _GEN332 : _GEN2231;
wire  _GEN2233 = io_x[18] ? _GEN2232 : _GEN2229;
wire  _GEN2234 = io_x[33] ? _GEN2233 : _GEN2225;
wire  _GEN2235 = io_x[23] ? _GEN332 : _GEN370;
wire  _GEN2236 = io_x[23] ? _GEN332 : _GEN370;
wire  _GEN2237 = io_x[18] ? _GEN2236 : _GEN2235;
wire  _GEN2238 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2239 = io_x[27] ? _GEN2238 : _GEN343;
wire  _GEN2240 = io_x[19] ? _GEN2239 : _GEN338;
wire  _GEN2241 = io_x[23] ? _GEN2240 : _GEN370;
wire  _GEN2242 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2243 = io_x[27] ? _GEN2242 : _GEN343;
wire  _GEN2244 = io_x[19] ? _GEN345 : _GEN2243;
wire  _GEN2245 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2246 = io_x[27] ? _GEN2245 : _GEN343;
wire  _GEN2247 = io_x[19] ? _GEN2246 : _GEN338;
wire  _GEN2248 = io_x[23] ? _GEN2247 : _GEN2244;
wire  _GEN2249 = io_x[18] ? _GEN2248 : _GEN2241;
wire  _GEN2250 = io_x[33] ? _GEN2249 : _GEN2237;
wire  _GEN2251 = io_x[31] ? _GEN2250 : _GEN2234;
wire  _GEN2252 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2253 = io_x[19] ? _GEN345 : _GEN2252;
wire  _GEN2254 = io_x[23] ? _GEN370 : _GEN2253;
wire  _GEN2255 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2256 = io_x[19] ? _GEN2255 : _GEN345;
wire  _GEN2257 = io_x[23] ? _GEN2256 : _GEN332;
wire  _GEN2258 = io_x[18] ? _GEN2257 : _GEN2254;
wire  _GEN2259 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2260 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2261 = io_x[27] ? _GEN2260 : _GEN343;
wire  _GEN2262 = io_x[19] ? _GEN2261 : _GEN2259;
wire  _GEN2263 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2264 = io_x[27] ? _GEN2263 : _GEN343;
wire  _GEN2265 = io_x[19] ? _GEN2264 : _GEN345;
wire  _GEN2266 = io_x[23] ? _GEN2265 : _GEN2262;
wire  _GEN2267 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2268 = io_x[27] ? _GEN2267 : _GEN343;
wire  _GEN2269 = io_x[19] ? _GEN2268 : _GEN338;
wire  _GEN2270 = io_x[23] ? _GEN2269 : _GEN332;
wire  _GEN2271 = io_x[18] ? _GEN2270 : _GEN2266;
wire  _GEN2272 = io_x[33] ? _GEN2271 : _GEN2258;
wire  _GEN2273 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN2274 = io_x[18] ? _GEN2273 : _GEN331;
wire  _GEN2275 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2276 = io_x[27] ? _GEN343 : _GEN2275;
wire  _GEN2277 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2278 = io_x[27] ? _GEN2277 : _GEN343;
wire  _GEN2279 = io_x[19] ? _GEN2278 : _GEN2276;
wire  _GEN2280 = io_x[23] ? _GEN2279 : _GEN332;
wire  _GEN2281 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2282 = io_x[27] ? _GEN336 : _GEN2281;
wire  _GEN2283 = io_x[19] ? _GEN345 : _GEN2282;
wire  _GEN2284 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2285 = io_x[27] ? _GEN336 : _GEN2284;
wire  _GEN2286 = io_x[19] ? _GEN2285 : _GEN338;
wire  _GEN2287 = io_x[23] ? _GEN2286 : _GEN2283;
wire  _GEN2288 = io_x[18] ? _GEN2287 : _GEN2280;
wire  _GEN2289 = io_x[33] ? _GEN2288 : _GEN2274;
wire  _GEN2290 = io_x[31] ? _GEN2289 : _GEN2272;
wire  _GEN2291 = io_x[28] ? _GEN2290 : _GEN2251;
wire  _GEN2292 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2293 = io_x[19] ? _GEN345 : _GEN2292;
wire  _GEN2294 = io_x[23] ? _GEN332 : _GEN2293;
wire  _GEN2295 = io_x[18] ? _GEN2294 : _GEN362;
wire  _GEN2296 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2297 = io_x[27] ? _GEN2296 : _GEN343;
wire  _GEN2298 = io_x[19] ? _GEN2297 : _GEN345;
wire  _GEN2299 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2300 = io_x[27] ? _GEN343 : _GEN2299;
wire  _GEN2301 = io_x[19] ? _GEN2300 : _GEN345;
wire  _GEN2302 = io_x[23] ? _GEN2301 : _GEN2298;
wire  _GEN2303 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2304 = io_x[27] ? _GEN343 : _GEN2303;
wire  _GEN2305 = io_x[19] ? _GEN2304 : _GEN338;
wire  _GEN2306 = io_x[23] ? _GEN332 : _GEN2305;
wire  _GEN2307 = io_x[18] ? _GEN2306 : _GEN2302;
wire  _GEN2308 = io_x[33] ? _GEN2307 : _GEN2295;
wire  _GEN2309 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2310 = io_x[27] ? _GEN2309 : _GEN343;
wire  _GEN2311 = io_x[19] ? _GEN2310 : _GEN338;
wire  _GEN2312 = io_x[23] ? _GEN370 : _GEN2311;
wire  _GEN2313 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2314 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2315 = io_x[27] ? _GEN2314 : _GEN2313;
wire  _GEN2316 = io_x[19] ? _GEN2315 : _GEN345;
wire  _GEN2317 = io_x[23] ? _GEN2316 : _GEN332;
wire  _GEN2318 = io_x[18] ? _GEN2317 : _GEN2312;
wire  _GEN2319 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2320 = io_x[27] ? _GEN2319 : _GEN343;
wire  _GEN2321 = io_x[19] ? _GEN2320 : _GEN345;
wire  _GEN2322 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2323 = io_x[27] ? _GEN336 : _GEN2322;
wire  _GEN2324 = io_x[19] ? _GEN2323 : _GEN338;
wire  _GEN2325 = io_x[23] ? _GEN2324 : _GEN2321;
wire  _GEN2326 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2327 = io_x[27] ? _GEN336 : _GEN2326;
wire  _GEN2328 = io_x[19] ? _GEN338 : _GEN2327;
wire  _GEN2329 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2330 = io_x[27] ? _GEN2329 : _GEN336;
wire  _GEN2331 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2332 = io_x[27] ? _GEN2331 : _GEN343;
wire  _GEN2333 = io_x[19] ? _GEN2332 : _GEN2330;
wire  _GEN2334 = io_x[23] ? _GEN2333 : _GEN2328;
wire  _GEN2335 = io_x[18] ? _GEN2334 : _GEN2325;
wire  _GEN2336 = io_x[33] ? _GEN2335 : _GEN2318;
wire  _GEN2337 = io_x[31] ? _GEN2336 : _GEN2308;
wire  _GEN2338 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2339 = io_x[27] ? _GEN2338 : _GEN343;
wire  _GEN2340 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2341 = io_x[27] ? _GEN343 : _GEN2340;
wire  _GEN2342 = io_x[19] ? _GEN2341 : _GEN2339;
wire  _GEN2343 = io_x[23] ? _GEN2342 : _GEN370;
wire  _GEN2344 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2345 = io_x[19] ? _GEN2344 : _GEN345;
wire  _GEN2346 = io_x[23] ? _GEN332 : _GEN2345;
wire  _GEN2347 = io_x[18] ? _GEN2346 : _GEN2343;
wire  _GEN2348 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2349 = io_x[27] ? _GEN343 : _GEN2348;
wire  _GEN2350 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2351 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2352 = io_x[27] ? _GEN2351 : _GEN2350;
wire  _GEN2353 = io_x[19] ? _GEN2352 : _GEN2349;
wire  _GEN2354 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2355 = io_x[27] ? _GEN2354 : _GEN343;
wire  _GEN2356 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2357 = io_x[27] ? _GEN343 : _GEN2356;
wire  _GEN2358 = io_x[19] ? _GEN2357 : _GEN2355;
wire  _GEN2359 = io_x[23] ? _GEN2358 : _GEN2353;
wire  _GEN2360 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2361 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2362 = io_x[19] ? _GEN2361 : _GEN2360;
wire  _GEN2363 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2364 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2365 = io_x[27] ? _GEN2364 : _GEN336;
wire  _GEN2366 = io_x[19] ? _GEN2365 : _GEN2363;
wire  _GEN2367 = io_x[23] ? _GEN2366 : _GEN2362;
wire  _GEN2368 = io_x[18] ? _GEN2367 : _GEN2359;
wire  _GEN2369 = io_x[33] ? _GEN2368 : _GEN2347;
wire  _GEN2370 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2371 = io_x[23] ? _GEN2370 : _GEN332;
wire  _GEN2372 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2373 = io_x[27] ? _GEN2372 : _GEN336;
wire  _GEN2374 = io_x[19] ? _GEN2373 : _GEN345;
wire  _GEN2375 = io_x[23] ? _GEN2374 : _GEN332;
wire  _GEN2376 = io_x[18] ? _GEN2375 : _GEN2371;
wire  _GEN2377 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2378 = io_x[27] ? _GEN343 : _GEN2377;
wire  _GEN2379 = io_x[19] ? _GEN2378 : _GEN338;
wire  _GEN2380 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2381 = io_x[27] ? _GEN2380 : _GEN343;
wire  _GEN2382 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2383 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2384 = io_x[27] ? _GEN2383 : _GEN2382;
wire  _GEN2385 = io_x[19] ? _GEN2384 : _GEN2381;
wire  _GEN2386 = io_x[23] ? _GEN2385 : _GEN2379;
wire  _GEN2387 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2388 = io_x[27] ? _GEN336 : _GEN2387;
wire  _GEN2389 = io_x[19] ? _GEN345 : _GEN2388;
wire  _GEN2390 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2391 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2392 = io_x[27] ? _GEN2391 : _GEN2390;
wire  _GEN2393 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2394 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2395 = io_x[27] ? _GEN2394 : _GEN2393;
wire  _GEN2396 = io_x[19] ? _GEN2395 : _GEN2392;
wire  _GEN2397 = io_x[23] ? _GEN2396 : _GEN2389;
wire  _GEN2398 = io_x[18] ? _GEN2397 : _GEN2386;
wire  _GEN2399 = io_x[33] ? _GEN2398 : _GEN2376;
wire  _GEN2400 = io_x[31] ? _GEN2399 : _GEN2369;
wire  _GEN2401 = io_x[28] ? _GEN2400 : _GEN2337;
wire  _GEN2402 = io_x[26] ? _GEN2401 : _GEN2291;
wire  _GEN2403 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2404 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2405 = io_x[27] ? _GEN2404 : _GEN343;
wire  _GEN2406 = io_x[19] ? _GEN2405 : _GEN2403;
wire  _GEN2407 = io_x[23] ? _GEN332 : _GEN2406;
wire  _GEN2408 = io_x[18] ? _GEN2407 : _GEN331;
wire  _GEN2409 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2410 = io_x[27] ? _GEN2409 : _GEN336;
wire  _GEN2411 = io_x[19] ? _GEN2410 : _GEN338;
wire  _GEN2412 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2413 = io_x[27] ? _GEN2412 : _GEN336;
wire  _GEN2414 = io_x[19] ? _GEN2413 : _GEN338;
wire  _GEN2415 = io_x[23] ? _GEN2414 : _GEN2411;
wire  _GEN2416 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2417 = io_x[27] ? _GEN2416 : _GEN343;
wire  _GEN2418 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2419 = io_x[27] ? _GEN2418 : _GEN336;
wire  _GEN2420 = io_x[19] ? _GEN2419 : _GEN2417;
wire  _GEN2421 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2422 = io_x[27] ? _GEN2421 : _GEN343;
wire  _GEN2423 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2424 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2425 = io_x[27] ? _GEN2424 : _GEN2423;
wire  _GEN2426 = io_x[19] ? _GEN2425 : _GEN2422;
wire  _GEN2427 = io_x[23] ? _GEN2426 : _GEN2420;
wire  _GEN2428 = io_x[18] ? _GEN2427 : _GEN2415;
wire  _GEN2429 = io_x[33] ? _GEN2428 : _GEN2408;
wire  _GEN2430 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2431 = io_x[19] ? _GEN345 : _GEN2430;
wire  _GEN2432 = io_x[23] ? _GEN2431 : _GEN332;
wire  _GEN2433 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2434 = io_x[19] ? _GEN338 : _GEN2433;
wire  _GEN2435 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2436 = io_x[27] ? _GEN2435 : _GEN343;
wire  _GEN2437 = io_x[19] ? _GEN2436 : _GEN338;
wire  _GEN2438 = io_x[23] ? _GEN2437 : _GEN2434;
wire  _GEN2439 = io_x[18] ? _GEN2438 : _GEN2432;
wire  _GEN2440 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2441 = io_x[27] ? _GEN2440 : _GEN343;
wire  _GEN2442 = io_x[19] ? _GEN2441 : _GEN345;
wire  _GEN2443 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2444 = io_x[27] ? _GEN2443 : _GEN336;
wire  _GEN2445 = io_x[19] ? _GEN2444 : _GEN345;
wire  _GEN2446 = io_x[23] ? _GEN2445 : _GEN2442;
wire  _GEN2447 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2448 = io_x[27] ? _GEN2447 : _GEN343;
wire  _GEN2449 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2450 = io_x[27] ? _GEN2449 : _GEN343;
wire  _GEN2451 = io_x[19] ? _GEN2450 : _GEN2448;
wire  _GEN2452 = io_x[23] ? _GEN370 : _GEN2451;
wire  _GEN2453 = io_x[18] ? _GEN2452 : _GEN2446;
wire  _GEN2454 = io_x[33] ? _GEN2453 : _GEN2439;
wire  _GEN2455 = io_x[31] ? _GEN2454 : _GEN2429;
wire  _GEN2456 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2457 = io_x[19] ? _GEN2456 : _GEN338;
wire  _GEN2458 = io_x[23] ? _GEN2457 : _GEN332;
wire  _GEN2459 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2460 = io_x[27] ? _GEN2459 : _GEN343;
wire  _GEN2461 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2462 = io_x[27] ? _GEN2461 : _GEN336;
wire  _GEN2463 = io_x[19] ? _GEN2462 : _GEN2460;
wire  _GEN2464 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2465 = io_x[27] ? _GEN2464 : _GEN343;
wire  _GEN2466 = io_x[19] ? _GEN2465 : _GEN345;
wire  _GEN2467 = io_x[23] ? _GEN2466 : _GEN2463;
wire  _GEN2468 = io_x[18] ? _GEN2467 : _GEN2458;
wire  _GEN2469 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2470 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2471 = io_x[27] ? _GEN2470 : _GEN2469;
wire  _GEN2472 = io_x[19] ? _GEN2471 : _GEN338;
wire  _GEN2473 = io_x[23] ? _GEN2472 : _GEN332;
wire  _GEN2474 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2475 = io_x[27] ? _GEN2474 : _GEN343;
wire  _GEN2476 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2477 = io_x[27] ? _GEN2476 : _GEN343;
wire  _GEN2478 = io_x[19] ? _GEN2477 : _GEN2475;
wire  _GEN2479 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2480 = io_x[27] ? _GEN343 : _GEN2479;
wire  _GEN2481 = io_x[19] ? _GEN2480 : _GEN338;
wire  _GEN2482 = io_x[23] ? _GEN2481 : _GEN2478;
wire  _GEN2483 = io_x[18] ? _GEN2482 : _GEN2473;
wire  _GEN2484 = io_x[33] ? _GEN2483 : _GEN2468;
wire  _GEN2485 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2486 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2487 = io_x[19] ? _GEN2486 : _GEN2485;
wire  _GEN2488 = io_x[23] ? _GEN2487 : _GEN332;
wire  _GEN2489 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2490 = io_x[27] ? _GEN336 : _GEN2489;
wire  _GEN2491 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2492 = io_x[27] ? _GEN2491 : _GEN343;
wire  _GEN2493 = io_x[19] ? _GEN2492 : _GEN2490;
wire  _GEN2494 = io_x[23] ? _GEN2493 : _GEN370;
wire  _GEN2495 = io_x[18] ? _GEN2494 : _GEN2488;
wire  _GEN2496 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2497 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2498 = io_x[27] ? _GEN2497 : _GEN2496;
wire  _GEN2499 = io_x[19] ? _GEN2498 : _GEN338;
wire  _GEN2500 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2501 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2502 = io_x[27] ? _GEN2501 : _GEN2500;
wire  _GEN2503 = io_x[19] ? _GEN2502 : _GEN345;
wire  _GEN2504 = io_x[23] ? _GEN2503 : _GEN2499;
wire  _GEN2505 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2506 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2507 = io_x[27] ? _GEN2506 : _GEN2505;
wire  _GEN2508 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2509 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2510 = io_x[27] ? _GEN2509 : _GEN2508;
wire  _GEN2511 = io_x[19] ? _GEN2510 : _GEN2507;
wire  _GEN2512 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2513 = io_x[27] ? _GEN2512 : _GEN343;
wire  _GEN2514 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2515 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2516 = io_x[27] ? _GEN2515 : _GEN2514;
wire  _GEN2517 = io_x[19] ? _GEN2516 : _GEN2513;
wire  _GEN2518 = io_x[23] ? _GEN2517 : _GEN2511;
wire  _GEN2519 = io_x[18] ? _GEN2518 : _GEN2504;
wire  _GEN2520 = io_x[33] ? _GEN2519 : _GEN2495;
wire  _GEN2521 = io_x[31] ? _GEN2520 : _GEN2484;
wire  _GEN2522 = io_x[28] ? _GEN2521 : _GEN2455;
wire  _GEN2523 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2524 = io_x[19] ? _GEN2523 : _GEN345;
wire  _GEN2525 = io_x[23] ? _GEN2524 : _GEN370;
wire  _GEN2526 = io_x[18] ? _GEN2525 : _GEN362;
wire  _GEN2527 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2528 = io_x[19] ? _GEN2527 : _GEN345;
wire  _GEN2529 = io_x[23] ? _GEN2528 : _GEN332;
wire  _GEN2530 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2531 = io_x[27] ? _GEN2530 : _GEN336;
wire  _GEN2532 = io_x[19] ? _GEN2531 : _GEN345;
wire  _GEN2533 = io_x[23] ? _GEN2532 : _GEN370;
wire  _GEN2534 = io_x[18] ? _GEN2533 : _GEN2529;
wire  _GEN2535 = io_x[33] ? _GEN2534 : _GEN2526;
wire  _GEN2536 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2537 = io_x[27] ? _GEN2536 : _GEN343;
wire  _GEN2538 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2539 = io_x[19] ? _GEN2538 : _GEN2537;
wire  _GEN2540 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2541 = io_x[27] ? _GEN2540 : _GEN343;
wire  _GEN2542 = io_x[19] ? _GEN2541 : _GEN345;
wire  _GEN2543 = io_x[23] ? _GEN2542 : _GEN2539;
wire  _GEN2544 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2545 = io_x[27] ? _GEN2544 : _GEN343;
wire  _GEN2546 = io_x[19] ? _GEN2545 : _GEN345;
wire  _GEN2547 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2548 = io_x[27] ? _GEN2547 : _GEN343;
wire  _GEN2549 = io_x[19] ? _GEN2548 : _GEN338;
wire  _GEN2550 = io_x[23] ? _GEN2549 : _GEN2546;
wire  _GEN2551 = io_x[18] ? _GEN2550 : _GEN2543;
wire  _GEN2552 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2553 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2554 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2555 = io_x[27] ? _GEN2554 : _GEN2553;
wire  _GEN2556 = io_x[19] ? _GEN2555 : _GEN2552;
wire  _GEN2557 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2558 = io_x[27] ? _GEN343 : _GEN2557;
wire  _GEN2559 = io_x[19] ? _GEN338 : _GEN2558;
wire  _GEN2560 = io_x[23] ? _GEN2559 : _GEN2556;
wire  _GEN2561 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2562 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2563 = io_x[27] ? _GEN2562 : _GEN2561;
wire  _GEN2564 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2565 = io_x[27] ? _GEN2564 : _GEN343;
wire  _GEN2566 = io_x[19] ? _GEN2565 : _GEN2563;
wire  _GEN2567 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2568 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2569 = io_x[27] ? _GEN2568 : _GEN2567;
wire  _GEN2570 = io_x[19] ? _GEN2569 : _GEN345;
wire  _GEN2571 = io_x[23] ? _GEN2570 : _GEN2566;
wire  _GEN2572 = io_x[18] ? _GEN2571 : _GEN2560;
wire  _GEN2573 = io_x[33] ? _GEN2572 : _GEN2551;
wire  _GEN2574 = io_x[31] ? _GEN2573 : _GEN2535;
wire  _GEN2575 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2576 = io_x[19] ? _GEN2575 : _GEN338;
wire  _GEN2577 = io_x[23] ? _GEN332 : _GEN2576;
wire  _GEN2578 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2579 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2580 = io_x[27] ? _GEN2579 : _GEN2578;
wire  _GEN2581 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2582 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2583 = io_x[27] ? _GEN2582 : _GEN2581;
wire  _GEN2584 = io_x[19] ? _GEN2583 : _GEN2580;
wire  _GEN2585 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2586 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2587 = io_x[27] ? _GEN2586 : _GEN343;
wire  _GEN2588 = io_x[19] ? _GEN2587 : _GEN2585;
wire  _GEN2589 = io_x[23] ? _GEN2588 : _GEN2584;
wire  _GEN2590 = io_x[18] ? _GEN2589 : _GEN2577;
wire  _GEN2591 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2592 = io_x[27] ? _GEN343 : _GEN2591;
wire  _GEN2593 = io_x[19] ? _GEN2592 : _GEN338;
wire  _GEN2594 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2595 = io_x[27] ? _GEN336 : _GEN2594;
wire  _GEN2596 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2597 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2598 = io_x[27] ? _GEN2597 : _GEN2596;
wire  _GEN2599 = io_x[19] ? _GEN2598 : _GEN2595;
wire  _GEN2600 = io_x[23] ? _GEN2599 : _GEN2593;
wire  _GEN2601 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2602 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2603 = io_x[27] ? _GEN2602 : _GEN2601;
wire  _GEN2604 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2605 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2606 = io_x[27] ? _GEN2605 : _GEN2604;
wire  _GEN2607 = io_x[19] ? _GEN2606 : _GEN2603;
wire  _GEN2608 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2609 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2610 = io_x[27] ? _GEN2609 : _GEN2608;
wire  _GEN2611 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2612 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2613 = io_x[27] ? _GEN2612 : _GEN2611;
wire  _GEN2614 = io_x[19] ? _GEN2613 : _GEN2610;
wire  _GEN2615 = io_x[23] ? _GEN2614 : _GEN2607;
wire  _GEN2616 = io_x[18] ? _GEN2615 : _GEN2600;
wire  _GEN2617 = io_x[33] ? _GEN2616 : _GEN2590;
wire  _GEN2618 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2619 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2620 = io_x[27] ? _GEN2619 : _GEN343;
wire  _GEN2621 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2622 = io_x[27] ? _GEN2621 : _GEN336;
wire  _GEN2623 = io_x[19] ? _GEN2622 : _GEN2620;
wire  _GEN2624 = io_x[23] ? _GEN2623 : _GEN2618;
wire  _GEN2625 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2626 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2627 = io_x[27] ? _GEN2626 : _GEN343;
wire  _GEN2628 = io_x[19] ? _GEN2627 : _GEN2625;
wire  _GEN2629 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2630 = io_x[27] ? _GEN2629 : _GEN343;
wire  _GEN2631 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2632 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2633 = io_x[27] ? _GEN2632 : _GEN2631;
wire  _GEN2634 = io_x[19] ? _GEN2633 : _GEN2630;
wire  _GEN2635 = io_x[23] ? _GEN2634 : _GEN2628;
wire  _GEN2636 = io_x[18] ? _GEN2635 : _GEN2624;
wire  _GEN2637 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2638 = io_x[27] ? _GEN2637 : _GEN343;
wire  _GEN2639 = io_x[19] ? _GEN2638 : _GEN345;
wire  _GEN2640 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2641 = io_x[27] ? _GEN2640 : _GEN336;
wire  _GEN2642 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2643 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2644 = io_x[27] ? _GEN2643 : _GEN2642;
wire  _GEN2645 = io_x[19] ? _GEN2644 : _GEN2641;
wire  _GEN2646 = io_x[23] ? _GEN2645 : _GEN2639;
wire  _GEN2647 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2648 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2649 = io_x[27] ? _GEN2648 : _GEN2647;
wire  _GEN2650 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2651 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2652 = io_x[27] ? _GEN2651 : _GEN2650;
wire  _GEN2653 = io_x[19] ? _GEN2652 : _GEN2649;
wire  _GEN2654 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2655 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2656 = io_x[27] ? _GEN2655 : _GEN2654;
wire  _GEN2657 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2658 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2659 = io_x[27] ? _GEN2658 : _GEN2657;
wire  _GEN2660 = io_x[19] ? _GEN2659 : _GEN2656;
wire  _GEN2661 = io_x[23] ? _GEN2660 : _GEN2653;
wire  _GEN2662 = io_x[18] ? _GEN2661 : _GEN2646;
wire  _GEN2663 = io_x[33] ? _GEN2662 : _GEN2636;
wire  _GEN2664 = io_x[31] ? _GEN2663 : _GEN2617;
wire  _GEN2665 = io_x[28] ? _GEN2664 : _GEN2574;
wire  _GEN2666 = io_x[26] ? _GEN2665 : _GEN2522;
wire  _GEN2667 = io_x[20] ? _GEN2666 : _GEN2402;
wire  _GEN2668 = io_x[24] ? _GEN2667 : _GEN2219;
wire  _GEN2669 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN2670 = io_x[18] ? _GEN362 : _GEN2669;
wire  _GEN2671 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2672 = io_x[27] ? _GEN2671 : _GEN343;
wire  _GEN2673 = io_x[19] ? _GEN2672 : _GEN338;
wire  _GEN2674 = io_x[23] ? _GEN2673 : _GEN332;
wire  _GEN2675 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2676 = io_x[19] ? _GEN338 : _GEN2675;
wire  _GEN2677 = io_x[23] ? _GEN2676 : _GEN332;
wire  _GEN2678 = io_x[18] ? _GEN2677 : _GEN2674;
wire  _GEN2679 = io_x[33] ? _GEN2678 : _GEN2670;
wire  _GEN2680 = io_x[23] ? _GEN332 : _GEN370;
wire  _GEN2681 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2682 = io_x[27] ? _GEN2681 : _GEN343;
wire  _GEN2683 = io_x[19] ? _GEN2682 : _GEN345;
wire  _GEN2684 = io_x[23] ? _GEN2683 : _GEN332;
wire  _GEN2685 = io_x[18] ? _GEN2684 : _GEN2680;
wire  _GEN2686 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2687 = io_x[27] ? _GEN2686 : _GEN343;
wire  _GEN2688 = io_x[19] ? _GEN2687 : _GEN345;
wire  _GEN2689 = io_x[23] ? _GEN2688 : _GEN332;
wire  _GEN2690 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2691 = io_x[27] ? _GEN2690 : _GEN343;
wire  _GEN2692 = io_x[19] ? _GEN2691 : _GEN345;
wire  _GEN2693 = io_x[23] ? _GEN2692 : _GEN332;
wire  _GEN2694 = io_x[18] ? _GEN2693 : _GEN2689;
wire  _GEN2695 = io_x[33] ? _GEN2694 : _GEN2685;
wire  _GEN2696 = io_x[31] ? _GEN2695 : _GEN2679;
wire  _GEN2697 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2698 = io_x[27] ? _GEN343 : _GEN2697;
wire  _GEN2699 = io_x[19] ? _GEN2698 : _GEN345;
wire  _GEN2700 = io_x[23] ? _GEN332 : _GEN2699;
wire  _GEN2701 = io_x[18] ? _GEN362 : _GEN2700;
wire  _GEN2702 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN2703 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2704 = io_x[27] ? _GEN2703 : _GEN343;
wire  _GEN2705 = io_x[19] ? _GEN2704 : _GEN338;
wire  _GEN2706 = io_x[23] ? _GEN2705 : _GEN2702;
wire  _GEN2707 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2708 = io_x[27] ? _GEN2707 : _GEN343;
wire  _GEN2709 = io_x[19] ? _GEN2708 : _GEN338;
wire  _GEN2710 = io_x[23] ? _GEN2709 : _GEN332;
wire  _GEN2711 = io_x[18] ? _GEN2710 : _GEN2706;
wire  _GEN2712 = io_x[33] ? _GEN2711 : _GEN2701;
wire  _GEN2713 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN2714 = io_x[18] ? _GEN2713 : _GEN331;
wire  _GEN2715 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2716 = io_x[19] ? _GEN338 : _GEN2715;
wire  _GEN2717 = io_x[23] ? _GEN2716 : _GEN370;
wire  _GEN2718 = io_x[18] ? _GEN2717 : _GEN331;
wire  _GEN2719 = io_x[33] ? _GEN2718 : _GEN2714;
wire  _GEN2720 = io_x[31] ? _GEN2719 : _GEN2712;
wire  _GEN2721 = io_x[28] ? _GEN2720 : _GEN2696;
wire  _GEN2722 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2723 = io_x[27] ? _GEN2722 : _GEN343;
wire  _GEN2724 = io_x[19] ? _GEN2723 : _GEN345;
wire  _GEN2725 = io_x[23] ? _GEN332 : _GEN2724;
wire  _GEN2726 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2727 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN2728 = io_x[23] ? _GEN2727 : _GEN2726;
wire  _GEN2729 = io_x[18] ? _GEN2728 : _GEN2725;
wire  _GEN2730 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2731 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2732 = io_x[19] ? _GEN2731 : _GEN345;
wire  _GEN2733 = io_x[23] ? _GEN2732 : _GEN2730;
wire  _GEN2734 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2735 = io_x[19] ? _GEN338 : _GEN2734;
wire  _GEN2736 = io_x[23] ? _GEN370 : _GEN2735;
wire  _GEN2737 = io_x[18] ? _GEN2736 : _GEN2733;
wire  _GEN2738 = io_x[33] ? _GEN2737 : _GEN2729;
wire  _GEN2739 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN2740 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2741 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2742 = io_x[27] ? _GEN2741 : _GEN336;
wire  _GEN2743 = io_x[19] ? _GEN2742 : _GEN2740;
wire  _GEN2744 = io_x[23] ? _GEN2743 : _GEN2739;
wire  _GEN2745 = io_x[18] ? _GEN2744 : _GEN362;
wire  _GEN2746 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2747 = io_x[19] ? _GEN345 : _GEN2746;
wire  _GEN2748 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2749 = io_x[19] ? _GEN2748 : _GEN338;
wire  _GEN2750 = io_x[23] ? _GEN2749 : _GEN2747;
wire  _GEN2751 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2752 = io_x[19] ? _GEN2751 : _GEN345;
wire  _GEN2753 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2754 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2755 = io_x[19] ? _GEN2754 : _GEN2753;
wire  _GEN2756 = io_x[23] ? _GEN2755 : _GEN2752;
wire  _GEN2757 = io_x[18] ? _GEN2756 : _GEN2750;
wire  _GEN2758 = io_x[33] ? _GEN2757 : _GEN2745;
wire  _GEN2759 = io_x[31] ? _GEN2758 : _GEN2738;
wire  _GEN2760 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2761 = io_x[27] ? _GEN343 : _GEN2760;
wire  _GEN2762 = io_x[19] ? _GEN2761 : _GEN345;
wire  _GEN2763 = io_x[23] ? _GEN2762 : _GEN370;
wire  _GEN2764 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2765 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2766 = io_x[27] ? _GEN343 : _GEN2765;
wire  _GEN2767 = io_x[19] ? _GEN2766 : _GEN2764;
wire  _GEN2768 = io_x[23] ? _GEN2767 : _GEN370;
wire  _GEN2769 = io_x[18] ? _GEN2768 : _GEN2763;
wire  _GEN2770 = io_x[33] ? _GEN2769 : _GEN1411;
wire  _GEN2771 = io_x[23] ? _GEN332 : _GEN370;
wire  _GEN2772 = io_x[18] ? _GEN2771 : _GEN362;
wire  _GEN2773 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN2774 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2775 = io_x[19] ? _GEN2774 : _GEN345;
wire  _GEN2776 = io_x[23] ? _GEN2775 : _GEN2773;
wire  _GEN2777 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2778 = io_x[19] ? _GEN345 : _GEN2777;
wire  _GEN2779 = io_x[23] ? _GEN2778 : _GEN370;
wire  _GEN2780 = io_x[18] ? _GEN2779 : _GEN2776;
wire  _GEN2781 = io_x[33] ? _GEN2780 : _GEN2772;
wire  _GEN2782 = io_x[31] ? _GEN2781 : _GEN2770;
wire  _GEN2783 = io_x[28] ? _GEN2782 : _GEN2759;
wire  _GEN2784 = io_x[26] ? _GEN2783 : _GEN2721;
wire  _GEN2785 = 1'b1;
wire  _GEN2786 = io_x[23] ? _GEN332 : _GEN370;
wire  _GEN2787 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2788 = io_x[27] ? _GEN2787 : _GEN343;
wire  _GEN2789 = io_x[19] ? _GEN2788 : _GEN345;
wire  _GEN2790 = io_x[23] ? _GEN2789 : _GEN332;
wire  _GEN2791 = io_x[18] ? _GEN2790 : _GEN2786;
wire  _GEN2792 = io_x[33] ? _GEN2791 : _GEN2785;
wire  _GEN2793 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN2794 = io_x[23] ? _GEN2793 : _GEN370;
wire  _GEN2795 = io_x[18] ? _GEN2794 : _GEN331;
wire  _GEN2796 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2797 = io_x[27] ? _GEN2796 : _GEN343;
wire  _GEN2798 = io_x[19] ? _GEN2797 : _GEN345;
wire  _GEN2799 = io_x[23] ? _GEN2798 : _GEN332;
wire  _GEN2800 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2801 = io_x[27] ? _GEN2800 : _GEN343;
wire  _GEN2802 = io_x[19] ? _GEN2801 : _GEN338;
wire  _GEN2803 = io_x[23] ? _GEN2802 : _GEN332;
wire  _GEN2804 = io_x[18] ? _GEN2803 : _GEN2799;
wire  _GEN2805 = io_x[33] ? _GEN2804 : _GEN2795;
wire  _GEN2806 = io_x[31] ? _GEN2805 : _GEN2792;
wire  _GEN2807 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2808 = io_x[23] ? _GEN2807 : _GEN370;
wire  _GEN2809 = io_x[18] ? _GEN2808 : _GEN362;
wire  _GEN2810 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN2811 = io_x[23] ? _GEN332 : _GEN2810;
wire  _GEN2812 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2813 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2814 = io_x[19] ? _GEN2813 : _GEN2812;
wire  _GEN2815 = io_x[23] ? _GEN2814 : _GEN370;
wire  _GEN2816 = io_x[18] ? _GEN2815 : _GEN2811;
wire  _GEN2817 = io_x[33] ? _GEN2816 : _GEN2809;
wire  _GEN2818 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2819 = io_x[23] ? _GEN2818 : _GEN332;
wire  _GEN2820 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2821 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2822 = io_x[27] ? _GEN2821 : _GEN2820;
wire  _GEN2823 = io_x[19] ? _GEN2822 : _GEN338;
wire  _GEN2824 = io_x[23] ? _GEN2823 : _GEN332;
wire  _GEN2825 = io_x[18] ? _GEN2824 : _GEN2819;
wire  _GEN2826 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2827 = io_x[27] ? _GEN2826 : _GEN336;
wire  _GEN2828 = io_x[19] ? _GEN2827 : _GEN338;
wire  _GEN2829 = io_x[23] ? _GEN2828 : _GEN370;
wire  _GEN2830 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2831 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2832 = io_x[27] ? _GEN2831 : _GEN2830;
wire  _GEN2833 = io_x[19] ? _GEN2832 : _GEN338;
wire  _GEN2834 = io_x[23] ? _GEN2833 : _GEN332;
wire  _GEN2835 = io_x[18] ? _GEN2834 : _GEN2829;
wire  _GEN2836 = io_x[33] ? _GEN2835 : _GEN2825;
wire  _GEN2837 = io_x[31] ? _GEN2836 : _GEN2817;
wire  _GEN2838 = io_x[28] ? _GEN2837 : _GEN2806;
wire  _GEN2839 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2840 = io_x[19] ? _GEN345 : _GEN2839;
wire  _GEN2841 = io_x[23] ? _GEN2840 : _GEN332;
wire  _GEN2842 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2843 = io_x[19] ? _GEN338 : _GEN2842;
wire  _GEN2844 = io_x[23] ? _GEN2843 : _GEN332;
wire  _GEN2845 = io_x[18] ? _GEN2844 : _GEN2841;
wire  _GEN2846 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2847 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2848 = io_x[27] ? _GEN343 : _GEN2847;
wire  _GEN2849 = io_x[19] ? _GEN345 : _GEN2848;
wire  _GEN2850 = io_x[23] ? _GEN2849 : _GEN2846;
wire  _GEN2851 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2852 = io_x[19] ? _GEN2851 : _GEN345;
wire  _GEN2853 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2854 = io_x[27] ? _GEN336 : _GEN2853;
wire  _GEN2855 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2856 = io_x[19] ? _GEN2855 : _GEN2854;
wire  _GEN2857 = io_x[23] ? _GEN2856 : _GEN2852;
wire  _GEN2858 = io_x[18] ? _GEN2857 : _GEN2850;
wire  _GEN2859 = io_x[33] ? _GEN2858 : _GEN2845;
wire  _GEN2860 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2861 = io_x[23] ? _GEN2860 : _GEN332;
wire  _GEN2862 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2863 = io_x[19] ? _GEN345 : _GEN2862;
wire  _GEN2864 = io_x[23] ? _GEN2863 : _GEN370;
wire  _GEN2865 = io_x[18] ? _GEN2864 : _GEN2861;
wire  _GEN2866 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2867 = io_x[27] ? _GEN343 : _GEN2866;
wire  _GEN2868 = io_x[19] ? _GEN338 : _GEN2867;
wire  _GEN2869 = io_x[23] ? _GEN2868 : _GEN332;
wire  _GEN2870 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2871 = io_x[19] ? _GEN2870 : _GEN338;
wire  _GEN2872 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2873 = io_x[27] ? _GEN2872 : _GEN336;
wire  _GEN2874 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2875 = io_x[27] ? _GEN2874 : _GEN343;
wire  _GEN2876 = io_x[19] ? _GEN2875 : _GEN2873;
wire  _GEN2877 = io_x[23] ? _GEN2876 : _GEN2871;
wire  _GEN2878 = io_x[18] ? _GEN2877 : _GEN2869;
wire  _GEN2879 = io_x[33] ? _GEN2878 : _GEN2865;
wire  _GEN2880 = io_x[31] ? _GEN2879 : _GEN2859;
wire  _GEN2881 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2882 = io_x[27] ? _GEN343 : _GEN2881;
wire  _GEN2883 = io_x[19] ? _GEN345 : _GEN2882;
wire  _GEN2884 = io_x[23] ? _GEN370 : _GEN2883;
wire  _GEN2885 = io_x[18] ? _GEN2884 : _GEN331;
wire  _GEN2886 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2887 = io_x[19] ? _GEN2886 : _GEN345;
wire  _GEN2888 = io_x[23] ? _GEN370 : _GEN2887;
wire  _GEN2889 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2890 = io_x[19] ? _GEN2889 : _GEN345;
wire  _GEN2891 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2892 = io_x[27] ? _GEN2891 : _GEN336;
wire  _GEN2893 = io_x[19] ? _GEN2892 : _GEN338;
wire  _GEN2894 = io_x[23] ? _GEN2893 : _GEN2890;
wire  _GEN2895 = io_x[18] ? _GEN2894 : _GEN2888;
wire  _GEN2896 = io_x[33] ? _GEN2895 : _GEN2885;
wire  _GEN2897 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN2898 = io_x[23] ? _GEN2897 : _GEN332;
wire  _GEN2899 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2900 = io_x[19] ? _GEN2899 : _GEN345;
wire  _GEN2901 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2902 = io_x[23] ? _GEN2901 : _GEN2900;
wire  _GEN2903 = io_x[18] ? _GEN2902 : _GEN2898;
wire  _GEN2904 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2905 = io_x[27] ? _GEN2904 : _GEN343;
wire  _GEN2906 = io_x[19] ? _GEN345 : _GEN2905;
wire  _GEN2907 = io_x[23] ? _GEN2906 : _GEN332;
wire  _GEN2908 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2909 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2910 = io_x[27] ? _GEN2909 : _GEN2908;
wire  _GEN2911 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2912 = io_x[27] ? _GEN2911 : _GEN336;
wire  _GEN2913 = io_x[19] ? _GEN2912 : _GEN2910;
wire  _GEN2914 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2915 = io_x[27] ? _GEN2914 : _GEN343;
wire  _GEN2916 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2917 = io_x[27] ? _GEN2916 : _GEN336;
wire  _GEN2918 = io_x[19] ? _GEN2917 : _GEN2915;
wire  _GEN2919 = io_x[23] ? _GEN2918 : _GEN2913;
wire  _GEN2920 = io_x[18] ? _GEN2919 : _GEN2907;
wire  _GEN2921 = io_x[33] ? _GEN2920 : _GEN2903;
wire  _GEN2922 = io_x[31] ? _GEN2921 : _GEN2896;
wire  _GEN2923 = io_x[28] ? _GEN2922 : _GEN2880;
wire  _GEN2924 = io_x[26] ? _GEN2923 : _GEN2838;
wire  _GEN2925 = io_x[20] ? _GEN2924 : _GEN2784;
wire  _GEN2926 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2927 = io_x[27] ? _GEN2926 : _GEN343;
wire  _GEN2928 = io_x[19] ? _GEN338 : _GEN2927;
wire  _GEN2929 = io_x[23] ? _GEN370 : _GEN2928;
wire  _GEN2930 = io_x[18] ? _GEN2929 : _GEN362;
wire  _GEN2931 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2932 = io_x[19] ? _GEN2931 : _GEN338;
wire  _GEN2933 = io_x[23] ? _GEN2932 : _GEN370;
wire  _GEN2934 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2935 = io_x[27] ? _GEN2934 : _GEN343;
wire  _GEN2936 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2937 = io_x[27] ? _GEN2936 : _GEN343;
wire  _GEN2938 = io_x[19] ? _GEN2937 : _GEN2935;
wire  _GEN2939 = io_x[23] ? _GEN332 : _GEN2938;
wire  _GEN2940 = io_x[18] ? _GEN2939 : _GEN2933;
wire  _GEN2941 = io_x[33] ? _GEN2940 : _GEN2930;
wire  _GEN2942 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN2943 = io_x[23] ? _GEN332 : _GEN2942;
wire  _GEN2944 = io_x[18] ? _GEN2943 : _GEN331;
wire  _GEN2945 = io_x[23] ? _GEN370 : _GEN332;
wire  _GEN2946 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN2947 = io_x[27] ? _GEN2946 : _GEN336;
wire  _GEN2948 = io_x[19] ? _GEN2947 : _GEN338;
wire  _GEN2949 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2950 = io_x[27] ? _GEN2949 : _GEN343;
wire  _GEN2951 = io_x[19] ? _GEN2950 : _GEN345;
wire  _GEN2952 = io_x[23] ? _GEN2951 : _GEN2948;
wire  _GEN2953 = io_x[18] ? _GEN2952 : _GEN2945;
wire  _GEN2954 = io_x[33] ? _GEN2953 : _GEN2944;
wire  _GEN2955 = io_x[31] ? _GEN2954 : _GEN2941;
wire  _GEN2956 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2957 = io_x[23] ? _GEN332 : _GEN2956;
wire  _GEN2958 = io_x[18] ? _GEN2957 : _GEN362;
wire  _GEN2959 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2960 = io_x[19] ? _GEN2959 : _GEN345;
wire  _GEN2961 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2962 = io_x[19] ? _GEN2961 : _GEN345;
wire  _GEN2963 = io_x[23] ? _GEN2962 : _GEN2960;
wire  _GEN2964 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2965 = io_x[19] ? _GEN2964 : _GEN338;
wire  _GEN2966 = io_x[23] ? _GEN2965 : _GEN332;
wire  _GEN2967 = io_x[18] ? _GEN2966 : _GEN2963;
wire  _GEN2968 = io_x[33] ? _GEN2967 : _GEN2958;
wire  _GEN2969 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN2970 = io_x[23] ? _GEN332 : _GEN2969;
wire  _GEN2971 = io_x[18] ? _GEN2970 : _GEN331;
wire  _GEN2972 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN2973 = io_x[23] ? _GEN2972 : _GEN332;
wire  _GEN2974 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2975 = io_x[19] ? _GEN345 : _GEN2974;
wire  _GEN2976 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2977 = io_x[19] ? _GEN2976 : _GEN345;
wire  _GEN2978 = io_x[23] ? _GEN2977 : _GEN2975;
wire  _GEN2979 = io_x[18] ? _GEN2978 : _GEN2973;
wire  _GEN2980 = io_x[33] ? _GEN2979 : _GEN2971;
wire  _GEN2981 = io_x[31] ? _GEN2980 : _GEN2968;
wire  _GEN2982 = io_x[28] ? _GEN2981 : _GEN2955;
wire  _GEN2983 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2984 = io_x[19] ? _GEN338 : _GEN2983;
wire  _GEN2985 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2986 = io_x[23] ? _GEN2985 : _GEN2984;
wire  _GEN2987 = io_x[18] ? _GEN2986 : _GEN362;
wire  _GEN2988 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN2989 = io_x[19] ? _GEN2988 : _GEN345;
wire  _GEN2990 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN2991 = io_x[19] ? _GEN2990 : _GEN345;
wire  _GEN2992 = io_x[23] ? _GEN2991 : _GEN2989;
wire  _GEN2993 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN2994 = io_x[27] ? _GEN343 : _GEN2993;
wire  _GEN2995 = io_x[19] ? _GEN338 : _GEN2994;
wire  _GEN2996 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN2997 = io_x[23] ? _GEN2996 : _GEN2995;
wire  _GEN2998 = io_x[18] ? _GEN2997 : _GEN2992;
wire  _GEN2999 = io_x[33] ? _GEN2998 : _GEN2987;
wire  _GEN3000 = io_x[18] ? _GEN362 : _GEN331;
wire  _GEN3001 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3002 = io_x[19] ? _GEN3001 : _GEN345;
wire  _GEN3003 = io_x[23] ? _GEN3002 : _GEN332;
wire  _GEN3004 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3005 = io_x[27] ? _GEN343 : _GEN3004;
wire  _GEN3006 = io_x[19] ? _GEN3005 : _GEN338;
wire  _GEN3007 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3008 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3009 = io_x[19] ? _GEN3008 : _GEN3007;
wire  _GEN3010 = io_x[23] ? _GEN3009 : _GEN3006;
wire  _GEN3011 = io_x[18] ? _GEN3010 : _GEN3003;
wire  _GEN3012 = io_x[33] ? _GEN3011 : _GEN3000;
wire  _GEN3013 = io_x[31] ? _GEN3012 : _GEN2999;
wire  _GEN3014 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3015 = io_x[27] ? _GEN343 : _GEN3014;
wire  _GEN3016 = io_x[19] ? _GEN3015 : _GEN345;
wire  _GEN3017 = io_x[23] ? _GEN3016 : _GEN332;
wire  _GEN3018 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3019 = io_x[27] ? _GEN3018 : _GEN343;
wire  _GEN3020 = io_x[19] ? _GEN3019 : _GEN338;
wire  _GEN3021 = io_x[23] ? _GEN3020 : _GEN332;
wire  _GEN3022 = io_x[18] ? _GEN3021 : _GEN3017;
wire  _GEN3023 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3024 = io_x[27] ? _GEN343 : _GEN3023;
wire  _GEN3025 = io_x[19] ? _GEN3024 : _GEN345;
wire  _GEN3026 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3027 = io_x[19] ? _GEN3026 : _GEN345;
wire  _GEN3028 = io_x[23] ? _GEN3027 : _GEN3025;
wire  _GEN3029 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3030 = io_x[27] ? _GEN343 : _GEN3029;
wire  _GEN3031 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3032 = io_x[27] ? _GEN343 : _GEN3031;
wire  _GEN3033 = io_x[19] ? _GEN3032 : _GEN3030;
wire  _GEN3034 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3035 = io_x[19] ? _GEN345 : _GEN3034;
wire  _GEN3036 = io_x[23] ? _GEN3035 : _GEN3033;
wire  _GEN3037 = io_x[18] ? _GEN3036 : _GEN3028;
wire  _GEN3038 = io_x[33] ? _GEN3037 : _GEN3022;
wire  _GEN3039 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3040 = io_x[27] ? _GEN3039 : _GEN343;
wire  _GEN3041 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3042 = io_x[19] ? _GEN3041 : _GEN3040;
wire  _GEN3043 = io_x[23] ? _GEN3042 : _GEN332;
wire  _GEN3044 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3045 = io_x[19] ? _GEN3044 : _GEN345;
wire  _GEN3046 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3047 = io_x[27] ? _GEN3046 : _GEN343;
wire  _GEN3048 = io_x[19] ? _GEN3047 : _GEN345;
wire  _GEN3049 = io_x[23] ? _GEN3048 : _GEN3045;
wire  _GEN3050 = io_x[18] ? _GEN3049 : _GEN3043;
wire  _GEN3051 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3052 = io_x[27] ? _GEN3051 : _GEN343;
wire  _GEN3053 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3054 = io_x[27] ? _GEN3053 : _GEN343;
wire  _GEN3055 = io_x[19] ? _GEN3054 : _GEN3052;
wire  _GEN3056 = io_x[23] ? _GEN3055 : _GEN370;
wire  _GEN3057 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3058 = io_x[27] ? _GEN336 : _GEN3057;
wire  _GEN3059 = io_x[19] ? _GEN338 : _GEN3058;
wire  _GEN3060 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3061 = io_x[27] ? _GEN3060 : _GEN343;
wire  _GEN3062 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3063 = io_x[27] ? _GEN3062 : _GEN343;
wire  _GEN3064 = io_x[19] ? _GEN3063 : _GEN3061;
wire  _GEN3065 = io_x[23] ? _GEN3064 : _GEN3059;
wire  _GEN3066 = io_x[18] ? _GEN3065 : _GEN3056;
wire  _GEN3067 = io_x[33] ? _GEN3066 : _GEN3050;
wire  _GEN3068 = io_x[31] ? _GEN3067 : _GEN3038;
wire  _GEN3069 = io_x[28] ? _GEN3068 : _GEN3013;
wire  _GEN3070 = io_x[26] ? _GEN3069 : _GEN2982;
wire  _GEN3071 = io_x[23] ? _GEN332 : _GEN370;
wire  _GEN3072 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3073 = io_x[27] ? _GEN3072 : _GEN343;
wire  _GEN3074 = io_x[19] ? _GEN345 : _GEN3073;
wire  _GEN3075 = io_x[23] ? _GEN370 : _GEN3074;
wire  _GEN3076 = io_x[18] ? _GEN3075 : _GEN3071;
wire  _GEN3077 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3078 = io_x[19] ? _GEN338 : _GEN3077;
wire  _GEN3079 = io_x[23] ? _GEN332 : _GEN3078;
wire  _GEN3080 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3081 = io_x[27] ? _GEN3080 : _GEN343;
wire  _GEN3082 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3083 = io_x[19] ? _GEN3082 : _GEN3081;
wire  _GEN3084 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3085 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3086 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3087 = io_x[27] ? _GEN3086 : _GEN3085;
wire  _GEN3088 = io_x[19] ? _GEN3087 : _GEN3084;
wire  _GEN3089 = io_x[23] ? _GEN3088 : _GEN3083;
wire  _GEN3090 = io_x[18] ? _GEN3089 : _GEN3079;
wire  _GEN3091 = io_x[33] ? _GEN3090 : _GEN3076;
wire  _GEN3092 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3093 = io_x[27] ? _GEN3092 : _GEN343;
wire  _GEN3094 = io_x[19] ? _GEN345 : _GEN3093;
wire  _GEN3095 = io_x[23] ? _GEN332 : _GEN3094;
wire  _GEN3096 = io_x[18] ? _GEN3095 : _GEN362;
wire  _GEN3097 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3098 = io_x[27] ? _GEN3097 : _GEN343;
wire  _GEN3099 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3100 = io_x[19] ? _GEN3099 : _GEN3098;
wire  _GEN3101 = io_x[23] ? _GEN3100 : _GEN332;
wire  _GEN3102 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3103 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3104 = io_x[19] ? _GEN3103 : _GEN3102;
wire  _GEN3105 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3106 = io_x[19] ? _GEN3105 : _GEN345;
wire  _GEN3107 = io_x[23] ? _GEN3106 : _GEN3104;
wire  _GEN3108 = io_x[18] ? _GEN3107 : _GEN3101;
wire  _GEN3109 = io_x[33] ? _GEN3108 : _GEN3096;
wire  _GEN3110 = io_x[31] ? _GEN3109 : _GEN3091;
wire  _GEN3111 = io_x[19] ? _GEN338 : _GEN345;
wire  _GEN3112 = io_x[23] ? _GEN332 : _GEN3111;
wire  _GEN3113 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3114 = io_x[27] ? _GEN3113 : _GEN343;
wire  _GEN3115 = io_x[19] ? _GEN338 : _GEN3114;
wire  _GEN3116 = io_x[23] ? _GEN370 : _GEN3115;
wire  _GEN3117 = io_x[18] ? _GEN3116 : _GEN3112;
wire  _GEN3118 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3119 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3120 = io_x[19] ? _GEN3119 : _GEN3118;
wire  _GEN3121 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3122 = io_x[19] ? _GEN3121 : _GEN338;
wire  _GEN3123 = io_x[23] ? _GEN3122 : _GEN3120;
wire  _GEN3124 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3125 = io_x[19] ? _GEN3124 : _GEN345;
wire  _GEN3126 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3127 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3128 = io_x[27] ? _GEN343 : _GEN3127;
wire  _GEN3129 = io_x[19] ? _GEN3128 : _GEN3126;
wire  _GEN3130 = io_x[23] ? _GEN3129 : _GEN3125;
wire  _GEN3131 = io_x[18] ? _GEN3130 : _GEN3123;
wire  _GEN3132 = io_x[33] ? _GEN3131 : _GEN3117;
wire  _GEN3133 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN3134 = io_x[23] ? _GEN3133 : _GEN332;
wire  _GEN3135 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3136 = io_x[27] ? _GEN3135 : _GEN336;
wire  _GEN3137 = io_x[19] ? _GEN345 : _GEN3136;
wire  _GEN3138 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3139 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3140 = io_x[27] ? _GEN3139 : _GEN343;
wire  _GEN3141 = io_x[19] ? _GEN3140 : _GEN3138;
wire  _GEN3142 = io_x[23] ? _GEN3141 : _GEN3137;
wire  _GEN3143 = io_x[18] ? _GEN3142 : _GEN3134;
wire  _GEN3144 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3145 = io_x[19] ? _GEN3144 : _GEN345;
wire  _GEN3146 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3147 = io_x[27] ? _GEN3146 : _GEN343;
wire  _GEN3148 = io_x[19] ? _GEN338 : _GEN3147;
wire  _GEN3149 = io_x[23] ? _GEN3148 : _GEN3145;
wire  _GEN3150 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3151 = io_x[27] ? _GEN343 : _GEN3150;
wire  _GEN3152 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3153 = io_x[27] ? _GEN343 : _GEN3152;
wire  _GEN3154 = io_x[19] ? _GEN3153 : _GEN3151;
wire  _GEN3155 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3156 = io_x[27] ? _GEN3155 : _GEN336;
wire  _GEN3157 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3158 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3159 = io_x[27] ? _GEN3158 : _GEN3157;
wire  _GEN3160 = io_x[19] ? _GEN3159 : _GEN3156;
wire  _GEN3161 = io_x[23] ? _GEN3160 : _GEN3154;
wire  _GEN3162 = io_x[18] ? _GEN3161 : _GEN3149;
wire  _GEN3163 = io_x[33] ? _GEN3162 : _GEN3143;
wire  _GEN3164 = io_x[31] ? _GEN3163 : _GEN3132;
wire  _GEN3165 = io_x[28] ? _GEN3164 : _GEN3110;
wire  _GEN3166 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3167 = io_x[19] ? _GEN345 : _GEN3166;
wire  _GEN3168 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3169 = io_x[19] ? _GEN345 : _GEN3168;
wire  _GEN3170 = io_x[23] ? _GEN3169 : _GEN3167;
wire  _GEN3171 = io_x[18] ? _GEN3170 : _GEN331;
wire  _GEN3172 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3173 = io_x[19] ? _GEN3172 : _GEN338;
wire  _GEN3174 = io_x[23] ? _GEN3173 : _GEN370;
wire  _GEN3175 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3176 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3177 = io_x[19] ? _GEN3176 : _GEN3175;
wire  _GEN3178 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3179 = io_x[27] ? _GEN3178 : _GEN343;
wire  _GEN3180 = io_x[19] ? _GEN3179 : _GEN345;
wire  _GEN3181 = io_x[23] ? _GEN3180 : _GEN3177;
wire  _GEN3182 = io_x[18] ? _GEN3181 : _GEN3174;
wire  _GEN3183 = io_x[33] ? _GEN3182 : _GEN3171;
wire  _GEN3184 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN3185 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3186 = io_x[19] ? _GEN3185 : _GEN338;
wire  _GEN3187 = io_x[23] ? _GEN3186 : _GEN3184;
wire  _GEN3188 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3189 = io_x[27] ? _GEN3188 : _GEN343;
wire  _GEN3190 = io_x[19] ? _GEN345 : _GEN3189;
wire  _GEN3191 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3192 = io_x[27] ? _GEN3191 : _GEN343;
wire  _GEN3193 = io_x[19] ? _GEN3192 : _GEN345;
wire  _GEN3194 = io_x[23] ? _GEN3193 : _GEN3190;
wire  _GEN3195 = io_x[18] ? _GEN3194 : _GEN3187;
wire  _GEN3196 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3197 = io_x[27] ? _GEN3196 : _GEN343;
wire  _GEN3198 = io_x[19] ? _GEN3197 : _GEN338;
wire  _GEN3199 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3200 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3201 = io_x[27] ? _GEN3200 : _GEN343;
wire  _GEN3202 = io_x[19] ? _GEN3201 : _GEN3199;
wire  _GEN3203 = io_x[23] ? _GEN3202 : _GEN3198;
wire  _GEN3204 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3205 = io_x[27] ? _GEN3204 : _GEN343;
wire  _GEN3206 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3207 = io_x[27] ? _GEN3206 : _GEN336;
wire  _GEN3208 = io_x[19] ? _GEN3207 : _GEN3205;
wire  _GEN3209 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3210 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3211 = io_x[27] ? _GEN3210 : _GEN3209;
wire  _GEN3212 = io_x[19] ? _GEN3211 : _GEN338;
wire  _GEN3213 = io_x[23] ? _GEN3212 : _GEN3208;
wire  _GEN3214 = io_x[18] ? _GEN3213 : _GEN3203;
wire  _GEN3215 = io_x[33] ? _GEN3214 : _GEN3195;
wire  _GEN3216 = io_x[31] ? _GEN3215 : _GEN3183;
wire  _GEN3217 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN3218 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3219 = io_x[27] ? _GEN3218 : _GEN343;
wire  _GEN3220 = io_x[19] ? _GEN3219 : _GEN345;
wire  _GEN3221 = io_x[23] ? _GEN3220 : _GEN3217;
wire  _GEN3222 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3223 = io_x[27] ? _GEN343 : _GEN3222;
wire  _GEN3224 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3225 = io_x[27] ? _GEN336 : _GEN3224;
wire  _GEN3226 = io_x[19] ? _GEN3225 : _GEN3223;
wire  _GEN3227 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3228 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3229 = io_x[27] ? _GEN3228 : _GEN343;
wire  _GEN3230 = io_x[19] ? _GEN3229 : _GEN3227;
wire  _GEN3231 = io_x[23] ? _GEN3230 : _GEN3226;
wire  _GEN3232 = io_x[18] ? _GEN3231 : _GEN3221;
wire  _GEN3233 = io_x[27] ? _GEN343 : _GEN336;
wire  _GEN3234 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3235 = io_x[27] ? _GEN343 : _GEN3234;
wire  _GEN3236 = io_x[19] ? _GEN3235 : _GEN3233;
wire  _GEN3237 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3238 = io_x[27] ? _GEN336 : _GEN3237;
wire  _GEN3239 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3240 = io_x[27] ? _GEN3239 : _GEN336;
wire  _GEN3241 = io_x[19] ? _GEN3240 : _GEN3238;
wire  _GEN3242 = io_x[23] ? _GEN3241 : _GEN3236;
wire  _GEN3243 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3244 = io_x[27] ? _GEN343 : _GEN3243;
wire  _GEN3245 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3246 = io_x[27] ? _GEN336 : _GEN3245;
wire  _GEN3247 = io_x[19] ? _GEN3246 : _GEN3244;
wire  _GEN3248 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3249 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3250 = io_x[27] ? _GEN3249 : _GEN3248;
wire  _GEN3251 = io_x[19] ? _GEN3250 : _GEN345;
wire  _GEN3252 = io_x[23] ? _GEN3251 : _GEN3247;
wire  _GEN3253 = io_x[18] ? _GEN3252 : _GEN3242;
wire  _GEN3254 = io_x[33] ? _GEN3253 : _GEN3232;
wire  _GEN3255 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3256 = io_x[27] ? _GEN3255 : _GEN336;
wire  _GEN3257 = io_x[19] ? _GEN3256 : _GEN338;
wire  _GEN3258 = io_x[23] ? _GEN3257 : _GEN370;
wire  _GEN3259 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3260 = io_x[27] ? _GEN336 : _GEN3259;
wire  _GEN3261 = io_x[19] ? _GEN345 : _GEN3260;
wire  _GEN3262 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3263 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3264 = io_x[27] ? _GEN3263 : _GEN3262;
wire  _GEN3265 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3266 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3267 = io_x[27] ? _GEN3266 : _GEN3265;
wire  _GEN3268 = io_x[19] ? _GEN3267 : _GEN3264;
wire  _GEN3269 = io_x[23] ? _GEN3268 : _GEN3261;
wire  _GEN3270 = io_x[18] ? _GEN3269 : _GEN3258;
wire  _GEN3271 = io_x[27] ? _GEN336 : _GEN343;
wire  _GEN3272 = io_x[19] ? _GEN338 : _GEN3271;
wire  _GEN3273 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3274 = io_x[27] ? _GEN3273 : _GEN336;
wire  _GEN3275 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3276 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3277 = io_x[27] ? _GEN3276 : _GEN3275;
wire  _GEN3278 = io_x[19] ? _GEN3277 : _GEN3274;
wire  _GEN3279 = io_x[23] ? _GEN3278 : _GEN3272;
wire  _GEN3280 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3281 = io_x[27] ? _GEN336 : _GEN3280;
wire  _GEN3282 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3283 = io_x[27] ? _GEN3282 : _GEN336;
wire  _GEN3284 = io_x[19] ? _GEN3283 : _GEN3281;
wire  _GEN3285 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3286 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3287 = io_x[27] ? _GEN3286 : _GEN3285;
wire  _GEN3288 = io_x[77] ? _GEN334 : _GEN333;
wire  _GEN3289 = io_x[77] ? _GEN333 : _GEN334;
wire  _GEN3290 = io_x[27] ? _GEN3289 : _GEN3288;
wire  _GEN3291 = io_x[19] ? _GEN3290 : _GEN3287;
wire  _GEN3292 = io_x[23] ? _GEN3291 : _GEN3284;
wire  _GEN3293 = io_x[18] ? _GEN3292 : _GEN3279;
wire  _GEN3294 = io_x[33] ? _GEN3293 : _GEN3270;
wire  _GEN3295 = io_x[31] ? _GEN3294 : _GEN3254;
wire  _GEN3296 = io_x[28] ? _GEN3295 : _GEN3216;
wire  _GEN3297 = io_x[26] ? _GEN3296 : _GEN3165;
wire  _GEN3298 = io_x[20] ? _GEN3297 : _GEN3070;
wire  _GEN3299 = io_x[24] ? _GEN3298 : _GEN2925;
wire  _GEN3300 = io_x[78] ? _GEN3299 : _GEN2668;
wire  _GEN3301 = io_x[72] ? _GEN3300 : _GEN1860;
assign io_y[18] = _GEN3301;
wire  _GEN3302 = 1'b1;
wire  _GEN3303 = 1'b0;
wire  _GEN3304 = 1'b1;
wire  _GEN3305 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3306 = 1'b1;
wire  _GEN3307 = io_x[26] ? _GEN3306 : _GEN3305;
wire  _GEN3308 = 1'b1;
wire  _GEN3309 = io_x[73] ? _GEN3308 : _GEN3307;
wire  _GEN3310 = io_x[33] ? _GEN3309 : _GEN3302;
wire  _GEN3311 = 1'b0;
wire  _GEN3312 = 1'b0;
wire  _GEN3313 = 1'b1;
wire  _GEN3314 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3315 = io_x[30] ? _GEN3314 : _GEN3304;
wire  _GEN3316 = io_x[26] ? _GEN3315 : _GEN3311;
wire  _GEN3317 = io_x[73] ? _GEN3308 : _GEN3316;
wire  _GEN3318 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3319 = io_x[30] ? _GEN3318 : _GEN3304;
wire  _GEN3320 = io_x[26] ? _GEN3319 : _GEN3311;
wire  _GEN3321 = io_x[73] ? _GEN3308 : _GEN3320;
wire  _GEN3322 = io_x[33] ? _GEN3321 : _GEN3317;
wire  _GEN3323 = io_x[28] ? _GEN3322 : _GEN3310;
wire  _GEN3324 = 1'b0;
wire  _GEN3325 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3326 = io_x[73] ? _GEN3325 : _GEN3324;
wire  _GEN3327 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3328 = io_x[30] ? _GEN3327 : _GEN3304;
wire  _GEN3329 = io_x[26] ? _GEN3328 : _GEN3311;
wire  _GEN3330 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3331 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3332 = io_x[30] ? _GEN3331 : _GEN3330;
wire  _GEN3333 = io_x[26] ? _GEN3311 : _GEN3332;
wire  _GEN3334 = io_x[73] ? _GEN3333 : _GEN3329;
wire  _GEN3335 = io_x[33] ? _GEN3334 : _GEN3326;
wire  _GEN3336 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3337 = io_x[26] ? _GEN3336 : _GEN3306;
wire  _GEN3338 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3339 = io_x[73] ? _GEN3338 : _GEN3337;
wire  _GEN3340 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3341 = io_x[30] ? _GEN3340 : _GEN3304;
wire  _GEN3342 = io_x[26] ? _GEN3341 : _GEN3306;
wire  _GEN3343 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3344 = io_x[30] ? _GEN3343 : _GEN3304;
wire  _GEN3345 = io_x[26] ? _GEN3311 : _GEN3344;
wire  _GEN3346 = io_x[73] ? _GEN3345 : _GEN3342;
wire  _GEN3347 = io_x[33] ? _GEN3346 : _GEN3339;
wire  _GEN3348 = io_x[28] ? _GEN3347 : _GEN3335;
wire  _GEN3349 = io_x[18] ? _GEN3348 : _GEN3323;
wire  _GEN3350 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3351 = io_x[26] ? _GEN3350 : _GEN3306;
wire  _GEN3352 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3353 = io_x[26] ? _GEN3352 : _GEN3306;
wire  _GEN3354 = io_x[73] ? _GEN3353 : _GEN3351;
wire  _GEN3355 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3356 = io_x[30] ? _GEN3355 : _GEN3303;
wire  _GEN3357 = io_x[26] ? _GEN3356 : _GEN3306;
wire  _GEN3358 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3359 = io_x[26] ? _GEN3358 : _GEN3306;
wire  _GEN3360 = io_x[73] ? _GEN3359 : _GEN3357;
wire  _GEN3361 = io_x[33] ? _GEN3360 : _GEN3354;
wire  _GEN3362 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3363 = io_x[30] ? _GEN3362 : _GEN3304;
wire  _GEN3364 = io_x[26] ? _GEN3363 : _GEN3311;
wire  _GEN3365 = io_x[73] ? _GEN3308 : _GEN3364;
wire  _GEN3366 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3367 = io_x[26] ? _GEN3366 : _GEN3311;
wire  _GEN3368 = io_x[73] ? _GEN3324 : _GEN3367;
wire  _GEN3369 = io_x[33] ? _GEN3368 : _GEN3365;
wire  _GEN3370 = io_x[28] ? _GEN3369 : _GEN3361;
wire  _GEN3371 = 1'b0;
wire  _GEN3372 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3373 = io_x[30] ? _GEN3372 : _GEN3304;
wire  _GEN3374 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3375 = io_x[30] ? _GEN3374 : _GEN3304;
wire  _GEN3376 = io_x[26] ? _GEN3375 : _GEN3373;
wire  _GEN3377 = io_x[73] ? _GEN3324 : _GEN3376;
wire  _GEN3378 = io_x[33] ? _GEN3377 : _GEN3371;
wire  _GEN3379 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3380 = io_x[30] ? _GEN3379 : _GEN3304;
wire  _GEN3381 = io_x[26] ? _GEN3380 : _GEN3306;
wire  _GEN3382 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3383 = io_x[73] ? _GEN3382 : _GEN3381;
wire  _GEN3384 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3385 = io_x[30] ? _GEN3384 : _GEN3303;
wire  _GEN3386 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3387 = io_x[26] ? _GEN3386 : _GEN3385;
wire  _GEN3388 = io_x[73] ? _GEN3387 : _GEN3324;
wire  _GEN3389 = io_x[33] ? _GEN3388 : _GEN3383;
wire  _GEN3390 = io_x[28] ? _GEN3389 : _GEN3378;
wire  _GEN3391 = io_x[18] ? _GEN3390 : _GEN3370;
wire  _GEN3392 = io_x[25] ? _GEN3391 : _GEN3349;
wire  _GEN3393 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3394 = io_x[73] ? _GEN3324 : _GEN3393;
wire  _GEN3395 = io_x[33] ? _GEN3394 : _GEN3371;
wire  _GEN3396 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3397 = io_x[30] ? _GEN3304 : _GEN3396;
wire  _GEN3398 = io_x[26] ? _GEN3311 : _GEN3397;
wire  _GEN3399 = io_x[73] ? _GEN3308 : _GEN3398;
wire  _GEN3400 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3401 = io_x[30] ? _GEN3304 : _GEN3400;
wire  _GEN3402 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3403 = io_x[26] ? _GEN3402 : _GEN3401;
wire  _GEN3404 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3405 = io_x[30] ? _GEN3404 : _GEN3304;
wire  _GEN3406 = io_x[26] ? _GEN3405 : _GEN3306;
wire  _GEN3407 = io_x[73] ? _GEN3406 : _GEN3403;
wire  _GEN3408 = io_x[33] ? _GEN3407 : _GEN3399;
wire  _GEN3409 = io_x[28] ? _GEN3408 : _GEN3395;
wire  _GEN3410 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3411 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN3412 = io_x[73] ? _GEN3411 : _GEN3410;
wire  _GEN3413 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3414 = io_x[26] ? _GEN3413 : _GEN3311;
wire  _GEN3415 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3416 = io_x[26] ? _GEN3415 : _GEN3306;
wire  _GEN3417 = io_x[73] ? _GEN3416 : _GEN3414;
wire  _GEN3418 = io_x[33] ? _GEN3417 : _GEN3412;
wire  _GEN3419 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3420 = io_x[26] ? _GEN3419 : _GEN3311;
wire  _GEN3421 = io_x[73] ? _GEN3420 : _GEN3324;
wire  _GEN3422 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3423 = io_x[30] ? _GEN3422 : _GEN3303;
wire  _GEN3424 = io_x[26] ? _GEN3423 : _GEN3306;
wire  _GEN3425 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3426 = io_x[26] ? _GEN3425 : _GEN3306;
wire  _GEN3427 = io_x[73] ? _GEN3426 : _GEN3424;
wire  _GEN3428 = io_x[33] ? _GEN3427 : _GEN3421;
wire  _GEN3429 = io_x[28] ? _GEN3428 : _GEN3418;
wire  _GEN3430 = io_x[18] ? _GEN3429 : _GEN3409;
wire  _GEN3431 = io_x[73] ? _GEN3324 : _GEN3308;
wire  _GEN3432 = io_x[33] ? _GEN3431 : _GEN3302;
wire  _GEN3433 = io_x[73] ? _GEN3308 : _GEN3324;
wire  _GEN3434 = io_x[33] ? _GEN3433 : _GEN3302;
wire  _GEN3435 = io_x[28] ? _GEN3434 : _GEN3432;
wire  _GEN3436 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3437 = io_x[26] ? _GEN3436 : _GEN3306;
wire  _GEN3438 = io_x[73] ? _GEN3324 : _GEN3437;
wire  _GEN3439 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3440 = io_x[30] ? _GEN3439 : _GEN3304;
wire  _GEN3441 = io_x[26] ? _GEN3311 : _GEN3440;
wire  _GEN3442 = io_x[73] ? _GEN3308 : _GEN3441;
wire  _GEN3443 = io_x[33] ? _GEN3442 : _GEN3438;
wire  _GEN3444 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3445 = io_x[30] ? _GEN3444 : _GEN3304;
wire  _GEN3446 = io_x[26] ? _GEN3445 : _GEN3306;
wire  _GEN3447 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3448 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3449 = io_x[26] ? _GEN3448 : _GEN3447;
wire  _GEN3450 = io_x[73] ? _GEN3449 : _GEN3446;
wire  _GEN3451 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3452 = io_x[30] ? _GEN3451 : _GEN3304;
wire  _GEN3453 = io_x[26] ? _GEN3452 : _GEN3306;
wire  _GEN3454 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3455 = io_x[30] ? _GEN3303 : _GEN3454;
wire  _GEN3456 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3457 = io_x[26] ? _GEN3456 : _GEN3455;
wire  _GEN3458 = io_x[73] ? _GEN3457 : _GEN3453;
wire  _GEN3459 = io_x[33] ? _GEN3458 : _GEN3450;
wire  _GEN3460 = io_x[28] ? _GEN3459 : _GEN3443;
wire  _GEN3461 = io_x[18] ? _GEN3460 : _GEN3435;
wire  _GEN3462 = io_x[25] ? _GEN3461 : _GEN3430;
wire  _GEN3463 = io_x[29] ? _GEN3462 : _GEN3392;
wire  _GEN3464 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3465 = io_x[73] ? _GEN3308 : _GEN3464;
wire  _GEN3466 = io_x[33] ? _GEN3465 : _GEN3302;
wire  _GEN3467 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3468 = io_x[73] ? _GEN3308 : _GEN3467;
wire  _GEN3469 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3470 = io_x[30] ? _GEN3469 : _GEN3304;
wire  _GEN3471 = io_x[26] ? _GEN3311 : _GEN3470;
wire  _GEN3472 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3473 = io_x[73] ? _GEN3472 : _GEN3471;
wire  _GEN3474 = io_x[33] ? _GEN3473 : _GEN3468;
wire  _GEN3475 = io_x[28] ? _GEN3474 : _GEN3466;
wire  _GEN3476 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3477 = io_x[30] ? _GEN3476 : _GEN3304;
wire  _GEN3478 = io_x[26] ? _GEN3477 : _GEN3311;
wire  _GEN3479 = io_x[73] ? _GEN3308 : _GEN3478;
wire  _GEN3480 = io_x[33] ? _GEN3371 : _GEN3479;
wire  _GEN3481 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3482 = io_x[26] ? _GEN3481 : _GEN3306;
wire  _GEN3483 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3484 = io_x[30] ? _GEN3303 : _GEN3483;
wire  _GEN3485 = io_x[26] ? _GEN3484 : _GEN3306;
wire  _GEN3486 = io_x[73] ? _GEN3485 : _GEN3482;
wire  _GEN3487 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3488 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3489 = io_x[30] ? _GEN3488 : _GEN3487;
wire  _GEN3490 = io_x[26] ? _GEN3489 : _GEN3306;
wire  _GEN3491 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3492 = io_x[30] ? _GEN3303 : _GEN3491;
wire  _GEN3493 = io_x[26] ? _GEN3492 : _GEN3311;
wire  _GEN3494 = io_x[73] ? _GEN3493 : _GEN3490;
wire  _GEN3495 = io_x[33] ? _GEN3494 : _GEN3486;
wire  _GEN3496 = io_x[28] ? _GEN3495 : _GEN3480;
wire  _GEN3497 = io_x[18] ? _GEN3496 : _GEN3475;
wire  _GEN3498 = 1'b1;
wire  _GEN3499 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN3500 = io_x[73] ? _GEN3499 : _GEN3308;
wire  _GEN3501 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3502 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3503 = io_x[30] ? _GEN3502 : _GEN3501;
wire  _GEN3504 = io_x[26] ? _GEN3503 : _GEN3306;
wire  _GEN3505 = io_x[73] ? _GEN3308 : _GEN3504;
wire  _GEN3506 = io_x[33] ? _GEN3505 : _GEN3500;
wire  _GEN3507 = io_x[28] ? _GEN3506 : _GEN3498;
wire  _GEN3508 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3509 = io_x[73] ? _GEN3308 : _GEN3508;
wire  _GEN3510 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3511 = io_x[73] ? _GEN3510 : _GEN3324;
wire  _GEN3512 = io_x[33] ? _GEN3511 : _GEN3509;
wire  _GEN3513 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3514 = io_x[30] ? _GEN3513 : _GEN3304;
wire  _GEN3515 = io_x[26] ? _GEN3311 : _GEN3514;
wire  _GEN3516 = io_x[73] ? _GEN3324 : _GEN3515;
wire  _GEN3517 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3518 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3519 = io_x[30] ? _GEN3303 : _GEN3518;
wire  _GEN3520 = io_x[26] ? _GEN3519 : _GEN3517;
wire  _GEN3521 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3522 = io_x[26] ? _GEN3311 : _GEN3521;
wire  _GEN3523 = io_x[73] ? _GEN3522 : _GEN3520;
wire  _GEN3524 = io_x[33] ? _GEN3523 : _GEN3516;
wire  _GEN3525 = io_x[28] ? _GEN3524 : _GEN3512;
wire  _GEN3526 = io_x[18] ? _GEN3525 : _GEN3507;
wire  _GEN3527 = io_x[25] ? _GEN3526 : _GEN3497;
wire  _GEN3528 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3529 = io_x[30] ? _GEN3303 : _GEN3528;
wire  _GEN3530 = io_x[26] ? _GEN3529 : _GEN3306;
wire  _GEN3531 = io_x[73] ? _GEN3308 : _GEN3530;
wire  _GEN3532 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3533 = io_x[26] ? _GEN3532 : _GEN3306;
wire  _GEN3534 = io_x[73] ? _GEN3308 : _GEN3533;
wire  _GEN3535 = io_x[33] ? _GEN3534 : _GEN3531;
wire  _GEN3536 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3537 = io_x[30] ? _GEN3303 : _GEN3536;
wire  _GEN3538 = io_x[26] ? _GEN3537 : _GEN3306;
wire  _GEN3539 = io_x[73] ? _GEN3324 : _GEN3538;
wire  _GEN3540 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3541 = io_x[30] ? _GEN3304 : _GEN3540;
wire  _GEN3542 = io_x[26] ? _GEN3541 : _GEN3306;
wire  _GEN3543 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3544 = io_x[30] ? _GEN3543 : _GEN3303;
wire  _GEN3545 = io_x[26] ? _GEN3544 : _GEN3311;
wire  _GEN3546 = io_x[73] ? _GEN3545 : _GEN3542;
wire  _GEN3547 = io_x[33] ? _GEN3546 : _GEN3539;
wire  _GEN3548 = io_x[28] ? _GEN3547 : _GEN3535;
wire  _GEN3549 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3550 = io_x[26] ? _GEN3549 : _GEN3311;
wire  _GEN3551 = io_x[73] ? _GEN3550 : _GEN3324;
wire  _GEN3552 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3553 = io_x[30] ? _GEN3552 : _GEN3303;
wire  _GEN3554 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3555 = io_x[26] ? _GEN3554 : _GEN3553;
wire  _GEN3556 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN3557 = io_x[73] ? _GEN3556 : _GEN3555;
wire  _GEN3558 = io_x[33] ? _GEN3557 : _GEN3551;
wire  _GEN3559 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3560 = io_x[30] ? _GEN3559 : _GEN3304;
wire  _GEN3561 = io_x[26] ? _GEN3560 : _GEN3306;
wire  _GEN3562 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3563 = io_x[30] ? _GEN3562 : _GEN3304;
wire  _GEN3564 = io_x[26] ? _GEN3563 : _GEN3306;
wire  _GEN3565 = io_x[73] ? _GEN3564 : _GEN3561;
wire  _GEN3566 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3567 = io_x[30] ? _GEN3566 : _GEN3304;
wire  _GEN3568 = io_x[26] ? _GEN3567 : _GEN3306;
wire  _GEN3569 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3570 = io_x[26] ? _GEN3306 : _GEN3569;
wire  _GEN3571 = io_x[73] ? _GEN3570 : _GEN3568;
wire  _GEN3572 = io_x[33] ? _GEN3571 : _GEN3565;
wire  _GEN3573 = io_x[28] ? _GEN3572 : _GEN3558;
wire  _GEN3574 = io_x[18] ? _GEN3573 : _GEN3548;
wire  _GEN3575 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3576 = io_x[30] ? _GEN3303 : _GEN3575;
wire  _GEN3577 = io_x[26] ? _GEN3311 : _GEN3576;
wire  _GEN3578 = io_x[73] ? _GEN3308 : _GEN3577;
wire  _GEN3579 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3580 = io_x[30] ? _GEN3303 : _GEN3579;
wire  _GEN3581 = io_x[26] ? _GEN3306 : _GEN3580;
wire  _GEN3582 = io_x[73] ? _GEN3308 : _GEN3581;
wire  _GEN3583 = io_x[33] ? _GEN3582 : _GEN3578;
wire  _GEN3584 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3585 = io_x[26] ? _GEN3584 : _GEN3311;
wire  _GEN3586 = io_x[73] ? _GEN3308 : _GEN3585;
wire  _GEN3587 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3588 = io_x[30] ? _GEN3587 : _GEN3303;
wire  _GEN3589 = io_x[26] ? _GEN3588 : _GEN3306;
wire  _GEN3590 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3591 = io_x[26] ? _GEN3311 : _GEN3590;
wire  _GEN3592 = io_x[73] ? _GEN3591 : _GEN3589;
wire  _GEN3593 = io_x[33] ? _GEN3592 : _GEN3586;
wire  _GEN3594 = io_x[28] ? _GEN3593 : _GEN3583;
wire  _GEN3595 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3596 = io_x[30] ? _GEN3595 : _GEN3304;
wire  _GEN3597 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3598 = io_x[30] ? _GEN3303 : _GEN3597;
wire  _GEN3599 = io_x[26] ? _GEN3598 : _GEN3596;
wire  _GEN3600 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3601 = io_x[26] ? _GEN3311 : _GEN3600;
wire  _GEN3602 = io_x[73] ? _GEN3601 : _GEN3599;
wire  _GEN3603 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3604 = io_x[26] ? _GEN3311 : _GEN3603;
wire  _GEN3605 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3606 = io_x[30] ? _GEN3304 : _GEN3605;
wire  _GEN3607 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3608 = io_x[26] ? _GEN3607 : _GEN3606;
wire  _GEN3609 = io_x[73] ? _GEN3608 : _GEN3604;
wire  _GEN3610 = io_x[33] ? _GEN3609 : _GEN3602;
wire  _GEN3611 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3612 = io_x[26] ? _GEN3611 : _GEN3306;
wire  _GEN3613 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3614 = io_x[30] ? _GEN3613 : _GEN3304;
wire  _GEN3615 = io_x[26] ? _GEN3614 : _GEN3311;
wire  _GEN3616 = io_x[73] ? _GEN3615 : _GEN3612;
wire  _GEN3617 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3618 = io_x[30] ? _GEN3617 : _GEN3304;
wire  _GEN3619 = io_x[26] ? _GEN3618 : _GEN3306;
wire  _GEN3620 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3621 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3622 = io_x[26] ? _GEN3621 : _GEN3620;
wire  _GEN3623 = io_x[73] ? _GEN3622 : _GEN3619;
wire  _GEN3624 = io_x[33] ? _GEN3623 : _GEN3616;
wire  _GEN3625 = io_x[28] ? _GEN3624 : _GEN3610;
wire  _GEN3626 = io_x[18] ? _GEN3625 : _GEN3594;
wire  _GEN3627 = io_x[25] ? _GEN3626 : _GEN3574;
wire  _GEN3628 = io_x[29] ? _GEN3627 : _GEN3527;
wire  _GEN3629 = io_x[23] ? _GEN3628 : _GEN3463;
wire  _GEN3630 = io_x[73] ? _GEN3308 : _GEN3324;
wire  _GEN3631 = io_x[33] ? _GEN3371 : _GEN3630;
wire  _GEN3632 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3633 = io_x[26] ? _GEN3306 : _GEN3632;
wire  _GEN3634 = io_x[73] ? _GEN3308 : _GEN3633;
wire  _GEN3635 = io_x[33] ? _GEN3371 : _GEN3634;
wire  _GEN3636 = io_x[28] ? _GEN3635 : _GEN3631;
wire  _GEN3637 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3638 = io_x[26] ? _GEN3637 : _GEN3306;
wire  _GEN3639 = io_x[73] ? _GEN3324 : _GEN3638;
wire  _GEN3640 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3641 = io_x[26] ? _GEN3311 : _GEN3640;
wire  _GEN3642 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3643 = io_x[30] ? _GEN3642 : _GEN3304;
wire  _GEN3644 = io_x[26] ? _GEN3643 : _GEN3311;
wire  _GEN3645 = io_x[73] ? _GEN3644 : _GEN3641;
wire  _GEN3646 = io_x[33] ? _GEN3645 : _GEN3639;
wire  _GEN3647 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3648 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3649 = io_x[30] ? _GEN3648 : _GEN3304;
wire  _GEN3650 = io_x[26] ? _GEN3649 : _GEN3647;
wire  _GEN3651 = io_x[73] ? _GEN3324 : _GEN3650;
wire  _GEN3652 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3653 = io_x[30] ? _GEN3304 : _GEN3652;
wire  _GEN3654 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3655 = io_x[30] ? _GEN3654 : _GEN3304;
wire  _GEN3656 = io_x[26] ? _GEN3655 : _GEN3653;
wire  _GEN3657 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3658 = io_x[26] ? _GEN3657 : _GEN3306;
wire  _GEN3659 = io_x[73] ? _GEN3658 : _GEN3656;
wire  _GEN3660 = io_x[33] ? _GEN3659 : _GEN3651;
wire  _GEN3661 = io_x[28] ? _GEN3660 : _GEN3646;
wire  _GEN3662 = io_x[18] ? _GEN3661 : _GEN3636;
wire  _GEN3663 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3664 = io_x[30] ? _GEN3663 : _GEN3304;
wire  _GEN3665 = io_x[26] ? _GEN3664 : _GEN3306;
wire  _GEN3666 = io_x[73] ? _GEN3324 : _GEN3665;
wire  _GEN3667 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3668 = io_x[30] ? _GEN3304 : _GEN3667;
wire  _GEN3669 = io_x[26] ? _GEN3668 : _GEN3306;
wire  _GEN3670 = io_x[73] ? _GEN3308 : _GEN3669;
wire  _GEN3671 = io_x[33] ? _GEN3670 : _GEN3666;
wire  _GEN3672 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3673 = io_x[30] ? _GEN3304 : _GEN3672;
wire  _GEN3674 = io_x[26] ? _GEN3311 : _GEN3673;
wire  _GEN3675 = io_x[73] ? _GEN3308 : _GEN3674;
wire  _GEN3676 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3677 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3678 = io_x[26] ? _GEN3677 : _GEN3676;
wire  _GEN3679 = io_x[73] ? _GEN3308 : _GEN3678;
wire  _GEN3680 = io_x[33] ? _GEN3679 : _GEN3675;
wire  _GEN3681 = io_x[28] ? _GEN3680 : _GEN3671;
wire  _GEN3682 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3683 = io_x[30] ? _GEN3682 : _GEN3304;
wire  _GEN3684 = io_x[26] ? _GEN3683 : _GEN3306;
wire  _GEN3685 = io_x[73] ? _GEN3684 : _GEN3308;
wire  _GEN3686 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3687 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3688 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3689 = io_x[30] ? _GEN3688 : _GEN3687;
wire  _GEN3690 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3691 = io_x[26] ? _GEN3690 : _GEN3689;
wire  _GEN3692 = io_x[73] ? _GEN3691 : _GEN3686;
wire  _GEN3693 = io_x[33] ? _GEN3692 : _GEN3685;
wire  _GEN3694 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3695 = io_x[26] ? _GEN3694 : _GEN3306;
wire  _GEN3696 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3697 = io_x[30] ? _GEN3696 : _GEN3304;
wire  _GEN3698 = io_x[26] ? _GEN3697 : _GEN3311;
wire  _GEN3699 = io_x[73] ? _GEN3698 : _GEN3695;
wire  _GEN3700 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3701 = io_x[30] ? _GEN3700 : _GEN3304;
wire  _GEN3702 = io_x[26] ? _GEN3701 : _GEN3306;
wire  _GEN3703 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3704 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3705 = io_x[30] ? _GEN3704 : _GEN3304;
wire  _GEN3706 = io_x[26] ? _GEN3705 : _GEN3703;
wire  _GEN3707 = io_x[73] ? _GEN3706 : _GEN3702;
wire  _GEN3708 = io_x[33] ? _GEN3707 : _GEN3699;
wire  _GEN3709 = io_x[28] ? _GEN3708 : _GEN3693;
wire  _GEN3710 = io_x[18] ? _GEN3709 : _GEN3681;
wire  _GEN3711 = io_x[25] ? _GEN3710 : _GEN3662;
wire  _GEN3712 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3713 = io_x[26] ? _GEN3306 : _GEN3712;
wire  _GEN3714 = io_x[73] ? _GEN3713 : _GEN3324;
wire  _GEN3715 = io_x[33] ? _GEN3714 : _GEN3302;
wire  _GEN3716 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3717 = io_x[30] ? _GEN3716 : _GEN3304;
wire  _GEN3718 = io_x[26] ? _GEN3717 : _GEN3306;
wire  _GEN3719 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3720 = io_x[73] ? _GEN3719 : _GEN3718;
wire  _GEN3721 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3722 = io_x[26] ? _GEN3721 : _GEN3306;
wire  _GEN3723 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3724 = io_x[30] ? _GEN3723 : _GEN3303;
wire  _GEN3725 = io_x[26] ? _GEN3724 : _GEN3306;
wire  _GEN3726 = io_x[73] ? _GEN3725 : _GEN3722;
wire  _GEN3727 = io_x[33] ? _GEN3726 : _GEN3720;
wire  _GEN3728 = io_x[28] ? _GEN3727 : _GEN3715;
wire  _GEN3729 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3730 = io_x[26] ? _GEN3729 : _GEN3306;
wire  _GEN3731 = io_x[73] ? _GEN3308 : _GEN3730;
wire  _GEN3732 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3733 = io_x[30] ? _GEN3732 : _GEN3304;
wire  _GEN3734 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3735 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3736 = io_x[30] ? _GEN3735 : _GEN3734;
wire  _GEN3737 = io_x[26] ? _GEN3736 : _GEN3733;
wire  _GEN3738 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3739 = io_x[26] ? _GEN3738 : _GEN3311;
wire  _GEN3740 = io_x[73] ? _GEN3739 : _GEN3737;
wire  _GEN3741 = io_x[33] ? _GEN3740 : _GEN3731;
wire  _GEN3742 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3743 = io_x[30] ? _GEN3304 : _GEN3742;
wire  _GEN3744 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3745 = io_x[30] ? _GEN3744 : _GEN3304;
wire  _GEN3746 = io_x[26] ? _GEN3745 : _GEN3743;
wire  _GEN3747 = io_x[73] ? _GEN3324 : _GEN3746;
wire  _GEN3748 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3749 = io_x[30] ? _GEN3748 : _GEN3303;
wire  _GEN3750 = io_x[26] ? _GEN3311 : _GEN3749;
wire  _GEN3751 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3752 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3753 = io_x[30] ? _GEN3752 : _GEN3304;
wire  _GEN3754 = io_x[26] ? _GEN3753 : _GEN3751;
wire  _GEN3755 = io_x[73] ? _GEN3754 : _GEN3750;
wire  _GEN3756 = io_x[33] ? _GEN3755 : _GEN3747;
wire  _GEN3757 = io_x[28] ? _GEN3756 : _GEN3741;
wire  _GEN3758 = io_x[18] ? _GEN3757 : _GEN3728;
wire  _GEN3759 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3760 = io_x[30] ? _GEN3759 : _GEN3304;
wire  _GEN3761 = io_x[26] ? _GEN3760 : _GEN3306;
wire  _GEN3762 = io_x[73] ? _GEN3324 : _GEN3761;
wire  _GEN3763 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3764 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3765 = io_x[30] ? _GEN3764 : _GEN3763;
wire  _GEN3766 = io_x[26] ? _GEN3765 : _GEN3311;
wire  _GEN3767 = io_x[73] ? _GEN3324 : _GEN3766;
wire  _GEN3768 = io_x[33] ? _GEN3767 : _GEN3762;
wire  _GEN3769 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3770 = io_x[73] ? _GEN3308 : _GEN3769;
wire  _GEN3771 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3772 = io_x[30] ? _GEN3771 : _GEN3304;
wire  _GEN3773 = io_x[26] ? _GEN3772 : _GEN3306;
wire  _GEN3774 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3775 = io_x[30] ? _GEN3774 : _GEN3303;
wire  _GEN3776 = io_x[26] ? _GEN3775 : _GEN3306;
wire  _GEN3777 = io_x[73] ? _GEN3776 : _GEN3773;
wire  _GEN3778 = io_x[33] ? _GEN3777 : _GEN3770;
wire  _GEN3779 = io_x[28] ? _GEN3778 : _GEN3768;
wire  _GEN3780 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN3781 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3782 = io_x[30] ? _GEN3304 : _GEN3781;
wire  _GEN3783 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3784 = io_x[30] ? _GEN3304 : _GEN3783;
wire  _GEN3785 = io_x[26] ? _GEN3784 : _GEN3782;
wire  _GEN3786 = io_x[73] ? _GEN3785 : _GEN3780;
wire  _GEN3787 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3788 = io_x[30] ? _GEN3304 : _GEN3787;
wire  _GEN3789 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3790 = io_x[30] ? _GEN3789 : _GEN3304;
wire  _GEN3791 = io_x[26] ? _GEN3790 : _GEN3788;
wire  _GEN3792 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3793 = io_x[30] ? _GEN3792 : _GEN3303;
wire  _GEN3794 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3795 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3796 = io_x[30] ? _GEN3795 : _GEN3794;
wire  _GEN3797 = io_x[26] ? _GEN3796 : _GEN3793;
wire  _GEN3798 = io_x[73] ? _GEN3797 : _GEN3791;
wire  _GEN3799 = io_x[33] ? _GEN3798 : _GEN3786;
wire  _GEN3800 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3801 = io_x[30] ? _GEN3800 : _GEN3304;
wire  _GEN3802 = io_x[26] ? _GEN3801 : _GEN3306;
wire  _GEN3803 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3804 = io_x[26] ? _GEN3803 : _GEN3306;
wire  _GEN3805 = io_x[73] ? _GEN3804 : _GEN3802;
wire  _GEN3806 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3807 = io_x[30] ? _GEN3806 : _GEN3303;
wire  _GEN3808 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3809 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3810 = io_x[30] ? _GEN3809 : _GEN3808;
wire  _GEN3811 = io_x[26] ? _GEN3810 : _GEN3807;
wire  _GEN3812 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3813 = io_x[30] ? _GEN3812 : _GEN3304;
wire  _GEN3814 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3815 = io_x[30] ? _GEN3814 : _GEN3304;
wire  _GEN3816 = io_x[26] ? _GEN3815 : _GEN3813;
wire  _GEN3817 = io_x[73] ? _GEN3816 : _GEN3811;
wire  _GEN3818 = io_x[33] ? _GEN3817 : _GEN3805;
wire  _GEN3819 = io_x[28] ? _GEN3818 : _GEN3799;
wire  _GEN3820 = io_x[18] ? _GEN3819 : _GEN3779;
wire  _GEN3821 = io_x[25] ? _GEN3820 : _GEN3758;
wire  _GEN3822 = io_x[29] ? _GEN3821 : _GEN3711;
wire  _GEN3823 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3824 = io_x[30] ? _GEN3823 : _GEN3304;
wire  _GEN3825 = io_x[26] ? _GEN3824 : _GEN3306;
wire  _GEN3826 = io_x[73] ? _GEN3308 : _GEN3825;
wire  _GEN3827 = io_x[33] ? _GEN3826 : _GEN3302;
wire  _GEN3828 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3829 = io_x[73] ? _GEN3828 : _GEN3308;
wire  _GEN3830 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3831 = io_x[30] ? _GEN3830 : _GEN3303;
wire  _GEN3832 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3833 = io_x[30] ? _GEN3304 : _GEN3832;
wire  _GEN3834 = io_x[26] ? _GEN3833 : _GEN3831;
wire  _GEN3835 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3836 = io_x[73] ? _GEN3835 : _GEN3834;
wire  _GEN3837 = io_x[33] ? _GEN3836 : _GEN3829;
wire  _GEN3838 = io_x[28] ? _GEN3837 : _GEN3827;
wire  _GEN3839 = io_x[73] ? _GEN3324 : _GEN3308;
wire  _GEN3840 = io_x[33] ? _GEN3839 : _GEN3302;
wire  _GEN3841 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3842 = io_x[30] ? _GEN3841 : _GEN3303;
wire  _GEN3843 = io_x[26] ? _GEN3842 : _GEN3306;
wire  _GEN3844 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3845 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3846 = io_x[30] ? _GEN3845 : _GEN3844;
wire  _GEN3847 = io_x[26] ? _GEN3846 : _GEN3311;
wire  _GEN3848 = io_x[73] ? _GEN3847 : _GEN3843;
wire  _GEN3849 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3850 = io_x[30] ? _GEN3849 : _GEN3303;
wire  _GEN3851 = io_x[26] ? _GEN3850 : _GEN3306;
wire  _GEN3852 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3853 = io_x[30] ? _GEN3304 : _GEN3852;
wire  _GEN3854 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3855 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3856 = io_x[30] ? _GEN3855 : _GEN3854;
wire  _GEN3857 = io_x[26] ? _GEN3856 : _GEN3853;
wire  _GEN3858 = io_x[73] ? _GEN3857 : _GEN3851;
wire  _GEN3859 = io_x[33] ? _GEN3858 : _GEN3848;
wire  _GEN3860 = io_x[28] ? _GEN3859 : _GEN3840;
wire  _GEN3861 = io_x[18] ? _GEN3860 : _GEN3838;
wire  _GEN3862 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3863 = io_x[73] ? _GEN3308 : _GEN3862;
wire  _GEN3864 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3865 = io_x[26] ? _GEN3864 : _GEN3311;
wire  _GEN3866 = io_x[73] ? _GEN3308 : _GEN3865;
wire  _GEN3867 = io_x[33] ? _GEN3866 : _GEN3863;
wire  _GEN3868 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN3869 = io_x[73] ? _GEN3308 : _GEN3868;
wire  _GEN3870 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3871 = io_x[30] ? _GEN3870 : _GEN3304;
wire  _GEN3872 = io_x[26] ? _GEN3871 : _GEN3306;
wire  _GEN3873 = io_x[73] ? _GEN3308 : _GEN3872;
wire  _GEN3874 = io_x[33] ? _GEN3873 : _GEN3869;
wire  _GEN3875 = io_x[28] ? _GEN3874 : _GEN3867;
wire  _GEN3876 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3877 = io_x[30] ? _GEN3303 : _GEN3876;
wire  _GEN3878 = io_x[26] ? _GEN3311 : _GEN3877;
wire  _GEN3879 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3880 = io_x[30] ? _GEN3879 : _GEN3304;
wire  _GEN3881 = io_x[26] ? _GEN3880 : _GEN3311;
wire  _GEN3882 = io_x[73] ? _GEN3881 : _GEN3878;
wire  _GEN3883 = io_x[33] ? _GEN3882 : _GEN3371;
wire  _GEN3884 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3885 = io_x[30] ? _GEN3884 : _GEN3304;
wire  _GEN3886 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3887 = io_x[30] ? _GEN3886 : _GEN3304;
wire  _GEN3888 = io_x[26] ? _GEN3887 : _GEN3885;
wire  _GEN3889 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3890 = io_x[30] ? _GEN3889 : _GEN3304;
wire  _GEN3891 = io_x[26] ? _GEN3890 : _GEN3306;
wire  _GEN3892 = io_x[73] ? _GEN3891 : _GEN3888;
wire  _GEN3893 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3894 = io_x[30] ? _GEN3893 : _GEN3304;
wire  _GEN3895 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3896 = io_x[30] ? _GEN3895 : _GEN3304;
wire  _GEN3897 = io_x[26] ? _GEN3896 : _GEN3894;
wire  _GEN3898 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3899 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3900 = io_x[30] ? _GEN3899 : _GEN3898;
wire  _GEN3901 = io_x[26] ? _GEN3900 : _GEN3306;
wire  _GEN3902 = io_x[73] ? _GEN3901 : _GEN3897;
wire  _GEN3903 = io_x[33] ? _GEN3902 : _GEN3892;
wire  _GEN3904 = io_x[28] ? _GEN3903 : _GEN3883;
wire  _GEN3905 = io_x[18] ? _GEN3904 : _GEN3875;
wire  _GEN3906 = io_x[25] ? _GEN3905 : _GEN3861;
wire  _GEN3907 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3908 = io_x[30] ? _GEN3907 : _GEN3304;
wire  _GEN3909 = io_x[26] ? _GEN3311 : _GEN3908;
wire  _GEN3910 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3911 = io_x[26] ? _GEN3306 : _GEN3910;
wire  _GEN3912 = io_x[73] ? _GEN3911 : _GEN3909;
wire  _GEN3913 = io_x[33] ? _GEN3912 : _GEN3302;
wire  _GEN3914 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN3915 = io_x[73] ? _GEN3308 : _GEN3914;
wire  _GEN3916 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3917 = io_x[30] ? _GEN3916 : _GEN3304;
wire  _GEN3918 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3919 = io_x[30] ? _GEN3918 : _GEN3303;
wire  _GEN3920 = io_x[26] ? _GEN3919 : _GEN3917;
wire  _GEN3921 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN3922 = io_x[73] ? _GEN3921 : _GEN3920;
wire  _GEN3923 = io_x[33] ? _GEN3922 : _GEN3915;
wire  _GEN3924 = io_x[28] ? _GEN3923 : _GEN3913;
wire  _GEN3925 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3926 = io_x[30] ? _GEN3304 : _GEN3925;
wire  _GEN3927 = io_x[26] ? _GEN3926 : _GEN3306;
wire  _GEN3928 = io_x[73] ? _GEN3308 : _GEN3927;
wire  _GEN3929 = io_x[73] ? _GEN3308 : _GEN3324;
wire  _GEN3930 = io_x[33] ? _GEN3929 : _GEN3928;
wire  _GEN3931 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3932 = io_x[30] ? _GEN3303 : _GEN3931;
wire  _GEN3933 = io_x[26] ? _GEN3932 : _GEN3306;
wire  _GEN3934 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3935 = io_x[26] ? _GEN3934 : _GEN3306;
wire  _GEN3936 = io_x[73] ? _GEN3935 : _GEN3933;
wire  _GEN3937 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3938 = io_x[26] ? _GEN3937 : _GEN3306;
wire  _GEN3939 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3940 = io_x[26] ? _GEN3939 : _GEN3306;
wire  _GEN3941 = io_x[73] ? _GEN3940 : _GEN3938;
wire  _GEN3942 = io_x[33] ? _GEN3941 : _GEN3936;
wire  _GEN3943 = io_x[28] ? _GEN3942 : _GEN3930;
wire  _GEN3944 = io_x[18] ? _GEN3943 : _GEN3924;
wire  _GEN3945 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3946 = io_x[30] ? _GEN3304 : _GEN3945;
wire  _GEN3947 = io_x[26] ? _GEN3306 : _GEN3946;
wire  _GEN3948 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN3949 = io_x[73] ? _GEN3948 : _GEN3947;
wire  _GEN3950 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3951 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3952 = io_x[30] ? _GEN3951 : _GEN3950;
wire  _GEN3953 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3954 = io_x[30] ? _GEN3953 : _GEN3303;
wire  _GEN3955 = io_x[26] ? _GEN3954 : _GEN3952;
wire  _GEN3956 = io_x[73] ? _GEN3308 : _GEN3955;
wire  _GEN3957 = io_x[33] ? _GEN3956 : _GEN3949;
wire  _GEN3958 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3959 = io_x[30] ? _GEN3958 : _GEN3303;
wire  _GEN3960 = io_x[26] ? _GEN3959 : _GEN3306;
wire  _GEN3961 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN3962 = io_x[26] ? _GEN3961 : _GEN3311;
wire  _GEN3963 = io_x[73] ? _GEN3962 : _GEN3960;
wire  _GEN3964 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3965 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3966 = io_x[30] ? _GEN3965 : _GEN3964;
wire  _GEN3967 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3968 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3969 = io_x[30] ? _GEN3968 : _GEN3967;
wire  _GEN3970 = io_x[26] ? _GEN3969 : _GEN3966;
wire  _GEN3971 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3972 = io_x[30] ? _GEN3971 : _GEN3304;
wire  _GEN3973 = io_x[26] ? _GEN3972 : _GEN3311;
wire  _GEN3974 = io_x[73] ? _GEN3973 : _GEN3970;
wire  _GEN3975 = io_x[33] ? _GEN3974 : _GEN3963;
wire  _GEN3976 = io_x[28] ? _GEN3975 : _GEN3957;
wire  _GEN3977 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3978 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3979 = io_x[30] ? _GEN3978 : _GEN3977;
wire  _GEN3980 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN3981 = io_x[26] ? _GEN3980 : _GEN3979;
wire  _GEN3982 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3983 = io_x[30] ? _GEN3304 : _GEN3982;
wire  _GEN3984 = io_x[26] ? _GEN3306 : _GEN3983;
wire  _GEN3985 = io_x[73] ? _GEN3984 : _GEN3981;
wire  _GEN3986 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3987 = io_x[30] ? _GEN3986 : _GEN3304;
wire  _GEN3988 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3989 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3990 = io_x[30] ? _GEN3989 : _GEN3988;
wire  _GEN3991 = io_x[26] ? _GEN3990 : _GEN3987;
wire  _GEN3992 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN3993 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3994 = io_x[30] ? _GEN3993 : _GEN3992;
wire  _GEN3995 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN3996 = io_x[30] ? _GEN3303 : _GEN3995;
wire  _GEN3997 = io_x[26] ? _GEN3996 : _GEN3994;
wire  _GEN3998 = io_x[73] ? _GEN3997 : _GEN3991;
wire  _GEN3999 = io_x[33] ? _GEN3998 : _GEN3985;
wire  _GEN4000 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4001 = io_x[30] ? _GEN3304 : _GEN4000;
wire  _GEN4002 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4003 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4004 = io_x[30] ? _GEN4003 : _GEN4002;
wire  _GEN4005 = io_x[26] ? _GEN4004 : _GEN4001;
wire  _GEN4006 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4007 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4008 = io_x[30] ? _GEN4007 : _GEN4006;
wire  _GEN4009 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4010 = io_x[30] ? _GEN4009 : _GEN3304;
wire  _GEN4011 = io_x[26] ? _GEN4010 : _GEN4008;
wire  _GEN4012 = io_x[73] ? _GEN4011 : _GEN4005;
wire  _GEN4013 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4014 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4015 = io_x[30] ? _GEN4014 : _GEN4013;
wire  _GEN4016 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4017 = io_x[30] ? _GEN4016 : _GEN3304;
wire  _GEN4018 = io_x[26] ? _GEN4017 : _GEN4015;
wire  _GEN4019 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4020 = io_x[30] ? _GEN3304 : _GEN4019;
wire  _GEN4021 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4022 = io_x[30] ? _GEN4021 : _GEN3304;
wire  _GEN4023 = io_x[26] ? _GEN4022 : _GEN4020;
wire  _GEN4024 = io_x[73] ? _GEN4023 : _GEN4018;
wire  _GEN4025 = io_x[33] ? _GEN4024 : _GEN4012;
wire  _GEN4026 = io_x[28] ? _GEN4025 : _GEN3999;
wire  _GEN4027 = io_x[18] ? _GEN4026 : _GEN3976;
wire  _GEN4028 = io_x[25] ? _GEN4027 : _GEN3944;
wire  _GEN4029 = io_x[29] ? _GEN4028 : _GEN3906;
wire  _GEN4030 = io_x[23] ? _GEN4029 : _GEN3822;
wire  _GEN4031 = io_x[31] ? _GEN4030 : _GEN3629;
wire  _GEN4032 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4033 = io_x[30] ? _GEN4032 : _GEN3304;
wire  _GEN4034 = io_x[26] ? _GEN4033 : _GEN3306;
wire  _GEN4035 = io_x[73] ? _GEN3308 : _GEN4034;
wire  _GEN4036 = io_x[33] ? _GEN4035 : _GEN3302;
wire  _GEN4037 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN4038 = io_x[73] ? _GEN4037 : _GEN3308;
wire  _GEN4039 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4040 = io_x[26] ? _GEN4039 : _GEN3306;
wire  _GEN4041 = io_x[73] ? _GEN3324 : _GEN4040;
wire  _GEN4042 = io_x[33] ? _GEN4041 : _GEN4038;
wire  _GEN4043 = io_x[28] ? _GEN4042 : _GEN4036;
wire  _GEN4044 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4045 = io_x[30] ? _GEN4044 : _GEN3304;
wire  _GEN4046 = io_x[26] ? _GEN4045 : _GEN3306;
wire  _GEN4047 = io_x[73] ? _GEN4046 : _GEN3308;
wire  _GEN4048 = io_x[33] ? _GEN4047 : _GEN3371;
wire  _GEN4049 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4050 = io_x[30] ? _GEN4049 : _GEN3304;
wire  _GEN4051 = io_x[26] ? _GEN4050 : _GEN3306;
wire  _GEN4052 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN4053 = io_x[73] ? _GEN4052 : _GEN4051;
wire  _GEN4054 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4055 = io_x[30] ? _GEN4054 : _GEN3304;
wire  _GEN4056 = io_x[26] ? _GEN3311 : _GEN4055;
wire  _GEN4057 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4058 = io_x[30] ? _GEN4057 : _GEN3304;
wire  _GEN4059 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4060 = io_x[30] ? _GEN4059 : _GEN3303;
wire  _GEN4061 = io_x[26] ? _GEN4060 : _GEN4058;
wire  _GEN4062 = io_x[73] ? _GEN4061 : _GEN4056;
wire  _GEN4063 = io_x[33] ? _GEN4062 : _GEN4053;
wire  _GEN4064 = io_x[28] ? _GEN4063 : _GEN4048;
wire  _GEN4065 = io_x[18] ? _GEN4064 : _GEN4043;
wire  _GEN4066 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN4067 = io_x[73] ? _GEN4066 : _GEN3308;
wire  _GEN4068 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4069 = io_x[26] ? _GEN4068 : _GEN3306;
wire  _GEN4070 = io_x[73] ? _GEN3308 : _GEN4069;
wire  _GEN4071 = io_x[33] ? _GEN4070 : _GEN4067;
wire  _GEN4072 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4073 = io_x[26] ? _GEN4072 : _GEN3306;
wire  _GEN4074 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4075 = io_x[30] ? _GEN4074 : _GEN3304;
wire  _GEN4076 = io_x[26] ? _GEN3306 : _GEN4075;
wire  _GEN4077 = io_x[73] ? _GEN4076 : _GEN4073;
wire  _GEN4078 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4079 = io_x[30] ? _GEN4078 : _GEN3304;
wire  _GEN4080 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4081 = io_x[30] ? _GEN4080 : _GEN3303;
wire  _GEN4082 = io_x[26] ? _GEN4081 : _GEN4079;
wire  _GEN4083 = io_x[73] ? _GEN3308 : _GEN4082;
wire  _GEN4084 = io_x[33] ? _GEN4083 : _GEN4077;
wire  _GEN4085 = io_x[28] ? _GEN4084 : _GEN4071;
wire  _GEN4086 = 1'b0;
wire  _GEN4087 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4088 = io_x[30] ? _GEN4087 : _GEN3304;
wire  _GEN4089 = io_x[26] ? _GEN4088 : _GEN3311;
wire  _GEN4090 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4091 = io_x[26] ? _GEN4090 : _GEN3306;
wire  _GEN4092 = io_x[73] ? _GEN4091 : _GEN4089;
wire  _GEN4093 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4094 = io_x[30] ? _GEN4093 : _GEN3304;
wire  _GEN4095 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4096 = io_x[30] ? _GEN4095 : _GEN3304;
wire  _GEN4097 = io_x[26] ? _GEN4096 : _GEN4094;
wire  _GEN4098 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4099 = io_x[26] ? _GEN3306 : _GEN4098;
wire  _GEN4100 = io_x[73] ? _GEN4099 : _GEN4097;
wire  _GEN4101 = io_x[33] ? _GEN4100 : _GEN4092;
wire  _GEN4102 = io_x[28] ? _GEN4101 : _GEN4086;
wire  _GEN4103 = io_x[18] ? _GEN4102 : _GEN4085;
wire  _GEN4104 = io_x[25] ? _GEN4103 : _GEN4065;
wire  _GEN4105 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4106 = io_x[30] ? _GEN3304 : _GEN4105;
wire  _GEN4107 = io_x[26] ? _GEN4106 : _GEN3306;
wire  _GEN4108 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN4109 = io_x[73] ? _GEN4108 : _GEN4107;
wire  _GEN4110 = io_x[33] ? _GEN4109 : _GEN3302;
wire  _GEN4111 = io_x[73] ? _GEN3308 : _GEN3324;
wire  _GEN4112 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4113 = io_x[30] ? _GEN4112 : _GEN3304;
wire  _GEN4114 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4115 = io_x[26] ? _GEN4114 : _GEN4113;
wire  _GEN4116 = io_x[73] ? _GEN3324 : _GEN4115;
wire  _GEN4117 = io_x[33] ? _GEN4116 : _GEN4111;
wire  _GEN4118 = io_x[28] ? _GEN4117 : _GEN4110;
wire  _GEN4119 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4120 = io_x[26] ? _GEN4119 : _GEN3306;
wire  _GEN4121 = io_x[73] ? _GEN4120 : _GEN3324;
wire  _GEN4122 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4123 = io_x[30] ? _GEN4122 : _GEN3304;
wire  _GEN4124 = io_x[26] ? _GEN4123 : _GEN3311;
wire  _GEN4125 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4126 = io_x[30] ? _GEN3303 : _GEN4125;
wire  _GEN4127 = io_x[26] ? _GEN4126 : _GEN3306;
wire  _GEN4128 = io_x[73] ? _GEN4127 : _GEN4124;
wire  _GEN4129 = io_x[33] ? _GEN4128 : _GEN4121;
wire  _GEN4130 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4131 = io_x[26] ? _GEN4130 : _GEN3306;
wire  _GEN4132 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4133 = io_x[26] ? _GEN4132 : _GEN3306;
wire  _GEN4134 = io_x[73] ? _GEN4133 : _GEN4131;
wire  _GEN4135 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4136 = io_x[26] ? _GEN3311 : _GEN4135;
wire  _GEN4137 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4138 = io_x[26] ? _GEN4137 : _GEN3306;
wire  _GEN4139 = io_x[73] ? _GEN4138 : _GEN4136;
wire  _GEN4140 = io_x[33] ? _GEN4139 : _GEN4134;
wire  _GEN4141 = io_x[28] ? _GEN4140 : _GEN4129;
wire  _GEN4142 = io_x[18] ? _GEN4141 : _GEN4118;
wire  _GEN4143 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4144 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4145 = io_x[26] ? _GEN4144 : _GEN4143;
wire  _GEN4146 = io_x[73] ? _GEN4145 : _GEN3324;
wire  _GEN4147 = io_x[33] ? _GEN4146 : _GEN3371;
wire  _GEN4148 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4149 = io_x[26] ? _GEN4148 : _GEN3306;
wire  _GEN4150 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4151 = io_x[30] ? _GEN3303 : _GEN4150;
wire  _GEN4152 = io_x[26] ? _GEN4151 : _GEN3311;
wire  _GEN4153 = io_x[73] ? _GEN4152 : _GEN4149;
wire  _GEN4154 = io_x[33] ? _GEN4153 : _GEN3302;
wire  _GEN4155 = io_x[28] ? _GEN4154 : _GEN4147;
wire  _GEN4156 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4157 = io_x[26] ? _GEN3306 : _GEN4156;
wire  _GEN4158 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4159 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4160 = io_x[26] ? _GEN4159 : _GEN4158;
wire  _GEN4161 = io_x[73] ? _GEN4160 : _GEN4157;
wire  _GEN4162 = io_x[33] ? _GEN4161 : _GEN3302;
wire  _GEN4163 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4164 = io_x[30] ? _GEN4163 : _GEN3304;
wire  _GEN4165 = io_x[26] ? _GEN4164 : _GEN3306;
wire  _GEN4166 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4167 = io_x[30] ? _GEN3304 : _GEN4166;
wire  _GEN4168 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4169 = io_x[30] ? _GEN4168 : _GEN3304;
wire  _GEN4170 = io_x[26] ? _GEN4169 : _GEN4167;
wire  _GEN4171 = io_x[73] ? _GEN4170 : _GEN4165;
wire  _GEN4172 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4173 = io_x[30] ? _GEN4172 : _GEN3304;
wire  _GEN4174 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4175 = io_x[30] ? _GEN4174 : _GEN3303;
wire  _GEN4176 = io_x[26] ? _GEN4175 : _GEN4173;
wire  _GEN4177 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4178 = io_x[30] ? _GEN4177 : _GEN3304;
wire  _GEN4179 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4180 = io_x[30] ? _GEN4179 : _GEN3304;
wire  _GEN4181 = io_x[26] ? _GEN4180 : _GEN4178;
wire  _GEN4182 = io_x[73] ? _GEN4181 : _GEN4176;
wire  _GEN4183 = io_x[33] ? _GEN4182 : _GEN4171;
wire  _GEN4184 = io_x[28] ? _GEN4183 : _GEN4162;
wire  _GEN4185 = io_x[18] ? _GEN4184 : _GEN4155;
wire  _GEN4186 = io_x[25] ? _GEN4185 : _GEN4142;
wire  _GEN4187 = io_x[29] ? _GEN4186 : _GEN4104;
wire  _GEN4188 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN4189 = io_x[73] ? _GEN4188 : _GEN3308;
wire  _GEN4190 = io_x[33] ? _GEN4189 : _GEN3302;
wire  _GEN4191 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN4192 = io_x[73] ? _GEN3324 : _GEN4191;
wire  _GEN4193 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4194 = io_x[30] ? _GEN4193 : _GEN3304;
wire  _GEN4195 = io_x[26] ? _GEN4194 : _GEN3306;
wire  _GEN4196 = io_x[73] ? _GEN3308 : _GEN4195;
wire  _GEN4197 = io_x[33] ? _GEN4196 : _GEN4192;
wire  _GEN4198 = io_x[28] ? _GEN4197 : _GEN4190;
wire  _GEN4199 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN4200 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4201 = io_x[30] ? _GEN4200 : _GEN3304;
wire  _GEN4202 = io_x[26] ? _GEN3311 : _GEN4201;
wire  _GEN4203 = io_x[73] ? _GEN4202 : _GEN4199;
wire  _GEN4204 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4205 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4206 = io_x[30] ? _GEN4205 : _GEN3304;
wire  _GEN4207 = io_x[26] ? _GEN4206 : _GEN4204;
wire  _GEN4208 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4209 = io_x[30] ? _GEN4208 : _GEN3304;
wire  _GEN4210 = io_x[26] ? _GEN4209 : _GEN3306;
wire  _GEN4211 = io_x[73] ? _GEN4210 : _GEN4207;
wire  _GEN4212 = io_x[33] ? _GEN4211 : _GEN4203;
wire  _GEN4213 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4214 = io_x[26] ? _GEN4213 : _GEN3311;
wire  _GEN4215 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4216 = io_x[30] ? _GEN4215 : _GEN3304;
wire  _GEN4217 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4218 = io_x[30] ? _GEN4217 : _GEN3304;
wire  _GEN4219 = io_x[26] ? _GEN4218 : _GEN4216;
wire  _GEN4220 = io_x[73] ? _GEN4219 : _GEN4214;
wire  _GEN4221 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4222 = io_x[30] ? _GEN3304 : _GEN4221;
wire  _GEN4223 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4224 = io_x[30] ? _GEN4223 : _GEN3304;
wire  _GEN4225 = io_x[26] ? _GEN4224 : _GEN4222;
wire  _GEN4226 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4227 = io_x[30] ? _GEN3303 : _GEN4226;
wire  _GEN4228 = io_x[26] ? _GEN4227 : _GEN3306;
wire  _GEN4229 = io_x[73] ? _GEN4228 : _GEN4225;
wire  _GEN4230 = io_x[33] ? _GEN4229 : _GEN4220;
wire  _GEN4231 = io_x[28] ? _GEN4230 : _GEN4212;
wire  _GEN4232 = io_x[18] ? _GEN4231 : _GEN4198;
wire  _GEN4233 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4234 = io_x[30] ? _GEN3304 : _GEN4233;
wire  _GEN4235 = io_x[26] ? _GEN3306 : _GEN4234;
wire  _GEN4236 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4237 = io_x[30] ? _GEN4236 : _GEN3304;
wire  _GEN4238 = io_x[26] ? _GEN3306 : _GEN4237;
wire  _GEN4239 = io_x[73] ? _GEN4238 : _GEN4235;
wire  _GEN4240 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN4241 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4242 = io_x[30] ? _GEN4241 : _GEN3304;
wire  _GEN4243 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4244 = io_x[30] ? _GEN4243 : _GEN3304;
wire  _GEN4245 = io_x[26] ? _GEN4244 : _GEN4242;
wire  _GEN4246 = io_x[73] ? _GEN4245 : _GEN4240;
wire  _GEN4247 = io_x[33] ? _GEN4246 : _GEN4239;
wire  _GEN4248 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4249 = io_x[30] ? _GEN4248 : _GEN3303;
wire  _GEN4250 = io_x[26] ? _GEN4249 : _GEN3311;
wire  _GEN4251 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4252 = io_x[26] ? _GEN4251 : _GEN3311;
wire  _GEN4253 = io_x[73] ? _GEN4252 : _GEN4250;
wire  _GEN4254 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4255 = io_x[30] ? _GEN4254 : _GEN3303;
wire  _GEN4256 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4257 = io_x[30] ? _GEN4256 : _GEN3303;
wire  _GEN4258 = io_x[26] ? _GEN4257 : _GEN4255;
wire  _GEN4259 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4260 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4261 = io_x[26] ? _GEN4260 : _GEN4259;
wire  _GEN4262 = io_x[73] ? _GEN4261 : _GEN4258;
wire  _GEN4263 = io_x[33] ? _GEN4262 : _GEN4253;
wire  _GEN4264 = io_x[28] ? _GEN4263 : _GEN4247;
wire  _GEN4265 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4266 = io_x[30] ? _GEN4265 : _GEN3304;
wire  _GEN4267 = io_x[26] ? _GEN4266 : _GEN3306;
wire  _GEN4268 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4269 = io_x[30] ? _GEN4268 : _GEN3304;
wire  _GEN4270 = io_x[26] ? _GEN4269 : _GEN3306;
wire  _GEN4271 = io_x[73] ? _GEN4270 : _GEN4267;
wire  _GEN4272 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4273 = io_x[26] ? _GEN4272 : _GEN3306;
wire  _GEN4274 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4275 = io_x[30] ? _GEN4274 : _GEN3303;
wire  _GEN4276 = io_x[26] ? _GEN3311 : _GEN4275;
wire  _GEN4277 = io_x[73] ? _GEN4276 : _GEN4273;
wire  _GEN4278 = io_x[33] ? _GEN4277 : _GEN4271;
wire  _GEN4279 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4280 = io_x[30] ? _GEN4279 : _GEN3304;
wire  _GEN4281 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4282 = io_x[26] ? _GEN4281 : _GEN4280;
wire  _GEN4283 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4284 = io_x[30] ? _GEN3303 : _GEN4283;
wire  _GEN4285 = io_x[26] ? _GEN4284 : _GEN3306;
wire  _GEN4286 = io_x[73] ? _GEN4285 : _GEN4282;
wire  _GEN4287 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4288 = io_x[30] ? _GEN4287 : _GEN3303;
wire  _GEN4289 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4290 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4291 = io_x[30] ? _GEN4290 : _GEN4289;
wire  _GEN4292 = io_x[26] ? _GEN4291 : _GEN4288;
wire  _GEN4293 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4294 = io_x[30] ? _GEN3303 : _GEN4293;
wire  _GEN4295 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4296 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4297 = io_x[30] ? _GEN4296 : _GEN4295;
wire  _GEN4298 = io_x[26] ? _GEN4297 : _GEN4294;
wire  _GEN4299 = io_x[73] ? _GEN4298 : _GEN4292;
wire  _GEN4300 = io_x[33] ? _GEN4299 : _GEN4286;
wire  _GEN4301 = io_x[28] ? _GEN4300 : _GEN4278;
wire  _GEN4302 = io_x[18] ? _GEN4301 : _GEN4264;
wire  _GEN4303 = io_x[25] ? _GEN4302 : _GEN4232;
wire  _GEN4304 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4305 = io_x[30] ? _GEN3303 : _GEN4304;
wire  _GEN4306 = io_x[26] ? _GEN4305 : _GEN3306;
wire  _GEN4307 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4308 = io_x[26] ? _GEN3306 : _GEN4307;
wire  _GEN4309 = io_x[73] ? _GEN4308 : _GEN4306;
wire  _GEN4310 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4311 = io_x[30] ? _GEN4310 : _GEN3304;
wire  _GEN4312 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4313 = io_x[30] ? _GEN3304 : _GEN4312;
wire  _GEN4314 = io_x[26] ? _GEN4313 : _GEN4311;
wire  _GEN4315 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4316 = io_x[26] ? _GEN4315 : _GEN3311;
wire  _GEN4317 = io_x[73] ? _GEN4316 : _GEN4314;
wire  _GEN4318 = io_x[33] ? _GEN4317 : _GEN4309;
wire  _GEN4319 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4320 = io_x[26] ? _GEN4319 : _GEN3306;
wire  _GEN4321 = io_x[73] ? _GEN3308 : _GEN4320;
wire  _GEN4322 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4323 = io_x[30] ? _GEN4322 : _GEN3303;
wire  _GEN4324 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4325 = io_x[30] ? _GEN4324 : _GEN3304;
wire  _GEN4326 = io_x[26] ? _GEN4325 : _GEN4323;
wire  _GEN4327 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4328 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4329 = io_x[26] ? _GEN4328 : _GEN4327;
wire  _GEN4330 = io_x[73] ? _GEN4329 : _GEN4326;
wire  _GEN4331 = io_x[33] ? _GEN4330 : _GEN4321;
wire  _GEN4332 = io_x[28] ? _GEN4331 : _GEN4318;
wire  _GEN4333 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4334 = io_x[26] ? _GEN3306 : _GEN4333;
wire  _GEN4335 = io_x[73] ? _GEN4334 : _GEN3324;
wire  _GEN4336 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4337 = io_x[30] ? _GEN4336 : _GEN3304;
wire  _GEN4338 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4339 = io_x[26] ? _GEN4338 : _GEN4337;
wire  _GEN4340 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4341 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4342 = io_x[26] ? _GEN4341 : _GEN4340;
wire  _GEN4343 = io_x[73] ? _GEN4342 : _GEN4339;
wire  _GEN4344 = io_x[33] ? _GEN4343 : _GEN4335;
wire  _GEN4345 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4346 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4347 = io_x[30] ? _GEN4346 : _GEN4345;
wire  _GEN4348 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4349 = io_x[26] ? _GEN4348 : _GEN4347;
wire  _GEN4350 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN4351 = io_x[73] ? _GEN4350 : _GEN4349;
wire  _GEN4352 = io_x[33] ? _GEN4351 : _GEN3371;
wire  _GEN4353 = io_x[28] ? _GEN4352 : _GEN4344;
wire  _GEN4354 = io_x[18] ? _GEN4353 : _GEN4332;
wire  _GEN4355 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4356 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4357 = io_x[30] ? _GEN4356 : _GEN4355;
wire  _GEN4358 = io_x[26] ? _GEN3306 : _GEN4357;
wire  _GEN4359 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4360 = io_x[30] ? _GEN4359 : _GEN3304;
wire  _GEN4361 = io_x[26] ? _GEN4360 : _GEN3311;
wire  _GEN4362 = io_x[73] ? _GEN4361 : _GEN4358;
wire  _GEN4363 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4364 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4365 = io_x[30] ? _GEN4364 : _GEN4363;
wire  _GEN4366 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4367 = io_x[30] ? _GEN4366 : _GEN3304;
wire  _GEN4368 = io_x[26] ? _GEN4367 : _GEN4365;
wire  _GEN4369 = io_x[73] ? _GEN3324 : _GEN4368;
wire  _GEN4370 = io_x[33] ? _GEN4369 : _GEN4362;
wire  _GEN4371 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4372 = io_x[30] ? _GEN4371 : _GEN3304;
wire  _GEN4373 = io_x[26] ? _GEN4372 : _GEN3311;
wire  _GEN4374 = io_x[73] ? _GEN3308 : _GEN4373;
wire  _GEN4375 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4376 = io_x[30] ? _GEN4375 : _GEN3303;
wire  _GEN4377 = io_x[26] ? _GEN4376 : _GEN3311;
wire  _GEN4378 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4379 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4380 = io_x[30] ? _GEN4379 : _GEN4378;
wire  _GEN4381 = io_x[26] ? _GEN4380 : _GEN3306;
wire  _GEN4382 = io_x[73] ? _GEN4381 : _GEN4377;
wire  _GEN4383 = io_x[33] ? _GEN4382 : _GEN4374;
wire  _GEN4384 = io_x[28] ? _GEN4383 : _GEN4370;
wire  _GEN4385 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4386 = io_x[26] ? _GEN4385 : _GEN3306;
wire  _GEN4387 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4388 = io_x[30] ? _GEN3304 : _GEN4387;
wire  _GEN4389 = io_x[26] ? _GEN3306 : _GEN4388;
wire  _GEN4390 = io_x[73] ? _GEN4389 : _GEN4386;
wire  _GEN4391 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4392 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4393 = io_x[26] ? _GEN4392 : _GEN4391;
wire  _GEN4394 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4395 = io_x[26] ? _GEN4394 : _GEN3306;
wire  _GEN4396 = io_x[73] ? _GEN4395 : _GEN4393;
wire  _GEN4397 = io_x[33] ? _GEN4396 : _GEN4390;
wire  _GEN4398 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4399 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4400 = io_x[30] ? _GEN4399 : _GEN3304;
wire  _GEN4401 = io_x[26] ? _GEN4400 : _GEN4398;
wire  _GEN4402 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4403 = io_x[30] ? _GEN4402 : _GEN3303;
wire  _GEN4404 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4405 = io_x[30] ? _GEN4404 : _GEN3304;
wire  _GEN4406 = io_x[26] ? _GEN4405 : _GEN4403;
wire  _GEN4407 = io_x[73] ? _GEN4406 : _GEN4401;
wire  _GEN4408 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4409 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4410 = io_x[30] ? _GEN4409 : _GEN4408;
wire  _GEN4411 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4412 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4413 = io_x[30] ? _GEN4412 : _GEN4411;
wire  _GEN4414 = io_x[26] ? _GEN4413 : _GEN4410;
wire  _GEN4415 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4416 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4417 = io_x[30] ? _GEN4416 : _GEN4415;
wire  _GEN4418 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4419 = io_x[30] ? _GEN4418 : _GEN3304;
wire  _GEN4420 = io_x[26] ? _GEN4419 : _GEN4417;
wire  _GEN4421 = io_x[73] ? _GEN4420 : _GEN4414;
wire  _GEN4422 = io_x[33] ? _GEN4421 : _GEN4407;
wire  _GEN4423 = io_x[28] ? _GEN4422 : _GEN4397;
wire  _GEN4424 = io_x[18] ? _GEN4423 : _GEN4384;
wire  _GEN4425 = io_x[25] ? _GEN4424 : _GEN4354;
wire  _GEN4426 = io_x[29] ? _GEN4425 : _GEN4303;
wire  _GEN4427 = io_x[23] ? _GEN4426 : _GEN4187;
wire  _GEN4428 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4429 = io_x[26] ? _GEN4428 : _GEN3306;
wire  _GEN4430 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4431 = io_x[26] ? _GEN3306 : _GEN4430;
wire  _GEN4432 = io_x[73] ? _GEN4431 : _GEN4429;
wire  _GEN4433 = io_x[33] ? _GEN4432 : _GEN3302;
wire  _GEN4434 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4435 = io_x[26] ? _GEN4434 : _GEN3306;
wire  _GEN4436 = io_x[73] ? _GEN3308 : _GEN4435;
wire  _GEN4437 = io_x[33] ? _GEN4436 : _GEN3302;
wire  _GEN4438 = io_x[28] ? _GEN4437 : _GEN4433;
wire  _GEN4439 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4440 = io_x[26] ? _GEN4439 : _GEN3306;
wire  _GEN4441 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4442 = io_x[30] ? _GEN4441 : _GEN3304;
wire  _GEN4443 = io_x[26] ? _GEN3306 : _GEN4442;
wire  _GEN4444 = io_x[73] ? _GEN4443 : _GEN4440;
wire  _GEN4445 = io_x[33] ? _GEN4444 : _GEN3371;
wire  _GEN4446 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4447 = io_x[30] ? _GEN4446 : _GEN3304;
wire  _GEN4448 = io_x[26] ? _GEN4447 : _GEN3311;
wire  _GEN4449 = io_x[73] ? _GEN4448 : _GEN3324;
wire  _GEN4450 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4451 = io_x[30] ? _GEN3304 : _GEN4450;
wire  _GEN4452 = io_x[26] ? _GEN3311 : _GEN4451;
wire  _GEN4453 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4454 = io_x[30] ? _GEN4453 : _GEN3303;
wire  _GEN4455 = io_x[26] ? _GEN4454 : _GEN3306;
wire  _GEN4456 = io_x[73] ? _GEN4455 : _GEN4452;
wire  _GEN4457 = io_x[33] ? _GEN4456 : _GEN4449;
wire  _GEN4458 = io_x[28] ? _GEN4457 : _GEN4445;
wire  _GEN4459 = io_x[18] ? _GEN4458 : _GEN4438;
wire  _GEN4460 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4461 = io_x[26] ? _GEN3306 : _GEN4460;
wire  _GEN4462 = io_x[73] ? _GEN3308 : _GEN4461;
wire  _GEN4463 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4464 = io_x[30] ? _GEN4463 : _GEN3304;
wire  _GEN4465 = io_x[26] ? _GEN3306 : _GEN4464;
wire  _GEN4466 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4467 = io_x[26] ? _GEN3311 : _GEN4466;
wire  _GEN4468 = io_x[73] ? _GEN4467 : _GEN4465;
wire  _GEN4469 = io_x[33] ? _GEN4468 : _GEN4462;
wire  _GEN4470 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4471 = io_x[26] ? _GEN3306 : _GEN4470;
wire  _GEN4472 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4473 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4474 = io_x[30] ? _GEN4473 : _GEN3304;
wire  _GEN4475 = io_x[26] ? _GEN4474 : _GEN4472;
wire  _GEN4476 = io_x[73] ? _GEN4475 : _GEN4471;
wire  _GEN4477 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4478 = io_x[30] ? _GEN4477 : _GEN3304;
wire  _GEN4479 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4480 = io_x[30] ? _GEN4479 : _GEN3303;
wire  _GEN4481 = io_x[26] ? _GEN4480 : _GEN4478;
wire  _GEN4482 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4483 = io_x[30] ? _GEN3303 : _GEN4482;
wire  _GEN4484 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4485 = io_x[30] ? _GEN4484 : _GEN3304;
wire  _GEN4486 = io_x[26] ? _GEN4485 : _GEN4483;
wire  _GEN4487 = io_x[73] ? _GEN4486 : _GEN4481;
wire  _GEN4488 = io_x[33] ? _GEN4487 : _GEN4476;
wire  _GEN4489 = io_x[28] ? _GEN4488 : _GEN4469;
wire  _GEN4490 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN4491 = io_x[73] ? _GEN3308 : _GEN4490;
wire  _GEN4492 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4493 = io_x[26] ? _GEN3311 : _GEN4492;
wire  _GEN4494 = io_x[73] ? _GEN4493 : _GEN3308;
wire  _GEN4495 = io_x[33] ? _GEN4494 : _GEN4491;
wire  _GEN4496 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4497 = io_x[30] ? _GEN3304 : _GEN4496;
wire  _GEN4498 = io_x[26] ? _GEN3311 : _GEN4497;
wire  _GEN4499 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4500 = io_x[30] ? _GEN4499 : _GEN3304;
wire  _GEN4501 = io_x[26] ? _GEN4500 : _GEN3306;
wire  _GEN4502 = io_x[73] ? _GEN4501 : _GEN4498;
wire  _GEN4503 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4504 = io_x[26] ? _GEN4503 : _GEN3306;
wire  _GEN4505 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4506 = io_x[30] ? _GEN3304 : _GEN4505;
wire  _GEN4507 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4508 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4509 = io_x[30] ? _GEN4508 : _GEN4507;
wire  _GEN4510 = io_x[26] ? _GEN4509 : _GEN4506;
wire  _GEN4511 = io_x[73] ? _GEN4510 : _GEN4504;
wire  _GEN4512 = io_x[33] ? _GEN4511 : _GEN4502;
wire  _GEN4513 = io_x[28] ? _GEN4512 : _GEN4495;
wire  _GEN4514 = io_x[18] ? _GEN4513 : _GEN4489;
wire  _GEN4515 = io_x[25] ? _GEN4514 : _GEN4459;
wire  _GEN4516 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4517 = io_x[30] ? _GEN4516 : _GEN3303;
wire  _GEN4518 = io_x[26] ? _GEN4517 : _GEN3306;
wire  _GEN4519 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4520 = io_x[30] ? _GEN3304 : _GEN4519;
wire  _GEN4521 = io_x[26] ? _GEN4520 : _GEN3306;
wire  _GEN4522 = io_x[73] ? _GEN4521 : _GEN4518;
wire  _GEN4523 = io_x[33] ? _GEN4522 : _GEN3302;
wire  _GEN4524 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN4525 = io_x[73] ? _GEN3308 : _GEN4524;
wire  _GEN4526 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4527 = io_x[30] ? _GEN4526 : _GEN3303;
wire  _GEN4528 = io_x[26] ? _GEN4527 : _GEN3311;
wire  _GEN4529 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4530 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4531 = io_x[30] ? _GEN4530 : _GEN4529;
wire  _GEN4532 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4533 = io_x[26] ? _GEN4532 : _GEN4531;
wire  _GEN4534 = io_x[73] ? _GEN4533 : _GEN4528;
wire  _GEN4535 = io_x[33] ? _GEN4534 : _GEN4525;
wire  _GEN4536 = io_x[28] ? _GEN4535 : _GEN4523;
wire  _GEN4537 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4538 = io_x[26] ? _GEN4537 : _GEN3306;
wire  _GEN4539 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4540 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4541 = io_x[30] ? _GEN3303 : _GEN4540;
wire  _GEN4542 = io_x[26] ? _GEN4541 : _GEN4539;
wire  _GEN4543 = io_x[73] ? _GEN4542 : _GEN4538;
wire  _GEN4544 = io_x[33] ? _GEN4543 : _GEN3302;
wire  _GEN4545 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4546 = io_x[30] ? _GEN4545 : _GEN3304;
wire  _GEN4547 = io_x[26] ? _GEN4546 : _GEN3311;
wire  _GEN4548 = io_x[73] ? _GEN4547 : _GEN3308;
wire  _GEN4549 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4550 = io_x[30] ? _GEN4549 : _GEN3304;
wire  _GEN4551 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4552 = io_x[30] ? _GEN4551 : _GEN3304;
wire  _GEN4553 = io_x[26] ? _GEN4552 : _GEN4550;
wire  _GEN4554 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4555 = io_x[30] ? _GEN4554 : _GEN3304;
wire  _GEN4556 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4557 = io_x[30] ? _GEN3303 : _GEN4556;
wire  _GEN4558 = io_x[26] ? _GEN4557 : _GEN4555;
wire  _GEN4559 = io_x[73] ? _GEN4558 : _GEN4553;
wire  _GEN4560 = io_x[33] ? _GEN4559 : _GEN4548;
wire  _GEN4561 = io_x[28] ? _GEN4560 : _GEN4544;
wire  _GEN4562 = io_x[18] ? _GEN4561 : _GEN4536;
wire  _GEN4563 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4564 = io_x[30] ? _GEN4563 : _GEN3304;
wire  _GEN4565 = io_x[26] ? _GEN4564 : _GEN3311;
wire  _GEN4566 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4567 = io_x[26] ? _GEN3306 : _GEN4566;
wire  _GEN4568 = io_x[73] ? _GEN4567 : _GEN4565;
wire  _GEN4569 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4570 = io_x[30] ? _GEN3304 : _GEN4569;
wire  _GEN4571 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4572 = io_x[30] ? _GEN4571 : _GEN3304;
wire  _GEN4573 = io_x[26] ? _GEN4572 : _GEN4570;
wire  _GEN4574 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4575 = io_x[30] ? _GEN3304 : _GEN4574;
wire  _GEN4576 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4577 = io_x[26] ? _GEN4576 : _GEN4575;
wire  _GEN4578 = io_x[73] ? _GEN4577 : _GEN4573;
wire  _GEN4579 = io_x[33] ? _GEN4578 : _GEN4568;
wire  _GEN4580 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4581 = io_x[30] ? _GEN4580 : _GEN3304;
wire  _GEN4582 = io_x[26] ? _GEN4581 : _GEN3306;
wire  _GEN4583 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4584 = io_x[30] ? _GEN3304 : _GEN4583;
wire  _GEN4585 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4586 = io_x[26] ? _GEN4585 : _GEN4584;
wire  _GEN4587 = io_x[73] ? _GEN4586 : _GEN4582;
wire  _GEN4588 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4589 = io_x[30] ? _GEN4588 : _GEN3304;
wire  _GEN4590 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4591 = io_x[30] ? _GEN4590 : _GEN3303;
wire  _GEN4592 = io_x[26] ? _GEN4591 : _GEN4589;
wire  _GEN4593 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4594 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4595 = io_x[30] ? _GEN4594 : _GEN4593;
wire  _GEN4596 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4597 = io_x[30] ? _GEN4596 : _GEN3303;
wire  _GEN4598 = io_x[26] ? _GEN4597 : _GEN4595;
wire  _GEN4599 = io_x[73] ? _GEN4598 : _GEN4592;
wire  _GEN4600 = io_x[33] ? _GEN4599 : _GEN4587;
wire  _GEN4601 = io_x[28] ? _GEN4600 : _GEN4579;
wire  _GEN4602 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4603 = io_x[30] ? _GEN3304 : _GEN4602;
wire  _GEN4604 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4605 = io_x[30] ? _GEN4604 : _GEN3304;
wire  _GEN4606 = io_x[26] ? _GEN4605 : _GEN4603;
wire  _GEN4607 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4608 = io_x[30] ? _GEN4607 : _GEN3303;
wire  _GEN4609 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4610 = io_x[30] ? _GEN4609 : _GEN3304;
wire  _GEN4611 = io_x[26] ? _GEN4610 : _GEN4608;
wire  _GEN4612 = io_x[73] ? _GEN4611 : _GEN4606;
wire  _GEN4613 = io_x[33] ? _GEN4612 : _GEN3371;
wire  _GEN4614 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4615 = io_x[30] ? _GEN4614 : _GEN3304;
wire  _GEN4616 = io_x[26] ? _GEN4615 : _GEN3311;
wire  _GEN4617 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4618 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4619 = io_x[30] ? _GEN4618 : _GEN3304;
wire  _GEN4620 = io_x[26] ? _GEN4619 : _GEN4617;
wire  _GEN4621 = io_x[73] ? _GEN4620 : _GEN4616;
wire  _GEN4622 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4623 = io_x[30] ? _GEN4622 : _GEN3303;
wire  _GEN4624 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4625 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4626 = io_x[30] ? _GEN4625 : _GEN4624;
wire  _GEN4627 = io_x[26] ? _GEN4626 : _GEN4623;
wire  _GEN4628 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4629 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4630 = io_x[30] ? _GEN4629 : _GEN4628;
wire  _GEN4631 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4632 = io_x[30] ? _GEN4631 : _GEN3304;
wire  _GEN4633 = io_x[26] ? _GEN4632 : _GEN4630;
wire  _GEN4634 = io_x[73] ? _GEN4633 : _GEN4627;
wire  _GEN4635 = io_x[33] ? _GEN4634 : _GEN4621;
wire  _GEN4636 = io_x[28] ? _GEN4635 : _GEN4613;
wire  _GEN4637 = io_x[18] ? _GEN4636 : _GEN4601;
wire  _GEN4638 = io_x[25] ? _GEN4637 : _GEN4562;
wire  _GEN4639 = io_x[29] ? _GEN4638 : _GEN4515;
wire  _GEN4640 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4641 = io_x[30] ? _GEN3304 : _GEN4640;
wire  _GEN4642 = io_x[26] ? _GEN3311 : _GEN4641;
wire  _GEN4643 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4644 = io_x[30] ? _GEN4643 : _GEN3304;
wire  _GEN4645 = io_x[26] ? _GEN4644 : _GEN3306;
wire  _GEN4646 = io_x[73] ? _GEN4645 : _GEN4642;
wire  _GEN4647 = io_x[33] ? _GEN4646 : _GEN3371;
wire  _GEN4648 = io_x[73] ? _GEN3308 : _GEN3324;
wire  _GEN4649 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4650 = io_x[30] ? _GEN4649 : _GEN3304;
wire  _GEN4651 = io_x[26] ? _GEN4650 : _GEN3311;
wire  _GEN4652 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4653 = io_x[30] ? _GEN3304 : _GEN4652;
wire  _GEN4654 = io_x[26] ? _GEN4653 : _GEN3311;
wire  _GEN4655 = io_x[73] ? _GEN4654 : _GEN4651;
wire  _GEN4656 = io_x[33] ? _GEN4655 : _GEN4648;
wire  _GEN4657 = io_x[28] ? _GEN4656 : _GEN4647;
wire  _GEN4658 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4659 = io_x[26] ? _GEN4658 : _GEN3311;
wire  _GEN4660 = io_x[73] ? _GEN4659 : _GEN3308;
wire  _GEN4661 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4662 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4663 = io_x[30] ? _GEN4662 : _GEN4661;
wire  _GEN4664 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4665 = io_x[26] ? _GEN4664 : _GEN4663;
wire  _GEN4666 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4667 = io_x[26] ? _GEN4666 : _GEN3311;
wire  _GEN4668 = io_x[73] ? _GEN4667 : _GEN4665;
wire  _GEN4669 = io_x[33] ? _GEN4668 : _GEN4660;
wire  _GEN4670 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4671 = io_x[30] ? _GEN4670 : _GEN3304;
wire  _GEN4672 = io_x[26] ? _GEN4671 : _GEN3311;
wire  _GEN4673 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4674 = io_x[26] ? _GEN4673 : _GEN3311;
wire  _GEN4675 = io_x[73] ? _GEN4674 : _GEN4672;
wire  _GEN4676 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4677 = io_x[30] ? _GEN4676 : _GEN3303;
wire  _GEN4678 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4679 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4680 = io_x[30] ? _GEN4679 : _GEN4678;
wire  _GEN4681 = io_x[26] ? _GEN4680 : _GEN4677;
wire  _GEN4682 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4683 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4684 = io_x[30] ? _GEN4683 : _GEN4682;
wire  _GEN4685 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4686 = io_x[26] ? _GEN4685 : _GEN4684;
wire  _GEN4687 = io_x[73] ? _GEN4686 : _GEN4681;
wire  _GEN4688 = io_x[33] ? _GEN4687 : _GEN4675;
wire  _GEN4689 = io_x[28] ? _GEN4688 : _GEN4669;
wire  _GEN4690 = io_x[18] ? _GEN4689 : _GEN4657;
wire  _GEN4691 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4692 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4693 = io_x[30] ? _GEN4692 : _GEN4691;
wire  _GEN4694 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4695 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4696 = io_x[30] ? _GEN4695 : _GEN4694;
wire  _GEN4697 = io_x[26] ? _GEN4696 : _GEN4693;
wire  _GEN4698 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4699 = io_x[30] ? _GEN4698 : _GEN3304;
wire  _GEN4700 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4701 = io_x[26] ? _GEN4700 : _GEN4699;
wire  _GEN4702 = io_x[73] ? _GEN4701 : _GEN4697;
wire  _GEN4703 = io_x[33] ? _GEN4702 : _GEN3371;
wire  _GEN4704 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4705 = io_x[30] ? _GEN3304 : _GEN4704;
wire  _GEN4706 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4707 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4708 = io_x[30] ? _GEN4707 : _GEN4706;
wire  _GEN4709 = io_x[26] ? _GEN4708 : _GEN4705;
wire  _GEN4710 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4711 = io_x[26] ? _GEN4710 : _GEN3306;
wire  _GEN4712 = io_x[73] ? _GEN4711 : _GEN4709;
wire  _GEN4713 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4714 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4715 = io_x[30] ? _GEN4714 : _GEN4713;
wire  _GEN4716 = io_x[26] ? _GEN4715 : _GEN3311;
wire  _GEN4717 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN4718 = io_x[73] ? _GEN4717 : _GEN4716;
wire  _GEN4719 = io_x[33] ? _GEN4718 : _GEN4712;
wire  _GEN4720 = io_x[28] ? _GEN4719 : _GEN4703;
wire  _GEN4721 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4722 = io_x[30] ? _GEN4721 : _GEN3304;
wire  _GEN4723 = io_x[26] ? _GEN4722 : _GEN3311;
wire  _GEN4724 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4725 = io_x[30] ? _GEN4724 : _GEN3304;
wire  _GEN4726 = io_x[26] ? _GEN4725 : _GEN3306;
wire  _GEN4727 = io_x[73] ? _GEN4726 : _GEN4723;
wire  _GEN4728 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4729 = io_x[30] ? _GEN4728 : _GEN3304;
wire  _GEN4730 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4731 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4732 = io_x[30] ? _GEN4731 : _GEN4730;
wire  _GEN4733 = io_x[26] ? _GEN4732 : _GEN4729;
wire  _GEN4734 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4735 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4736 = io_x[30] ? _GEN3303 : _GEN4735;
wire  _GEN4737 = io_x[26] ? _GEN4736 : _GEN4734;
wire  _GEN4738 = io_x[73] ? _GEN4737 : _GEN4733;
wire  _GEN4739 = io_x[33] ? _GEN4738 : _GEN4727;
wire  _GEN4740 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4741 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4742 = io_x[30] ? _GEN4741 : _GEN4740;
wire  _GEN4743 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4744 = io_x[30] ? _GEN4743 : _GEN3304;
wire  _GEN4745 = io_x[26] ? _GEN4744 : _GEN4742;
wire  _GEN4746 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4747 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4748 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4749 = io_x[30] ? _GEN4748 : _GEN4747;
wire  _GEN4750 = io_x[26] ? _GEN4749 : _GEN4746;
wire  _GEN4751 = io_x[73] ? _GEN4750 : _GEN4745;
wire  _GEN4752 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4753 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4754 = io_x[30] ? _GEN4753 : _GEN4752;
wire  _GEN4755 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4756 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4757 = io_x[30] ? _GEN4756 : _GEN4755;
wire  _GEN4758 = io_x[26] ? _GEN4757 : _GEN4754;
wire  _GEN4759 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4760 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4761 = io_x[30] ? _GEN4760 : _GEN4759;
wire  _GEN4762 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4763 = io_x[30] ? _GEN4762 : _GEN3304;
wire  _GEN4764 = io_x[26] ? _GEN4763 : _GEN4761;
wire  _GEN4765 = io_x[73] ? _GEN4764 : _GEN4758;
wire  _GEN4766 = io_x[33] ? _GEN4765 : _GEN4751;
wire  _GEN4767 = io_x[28] ? _GEN4766 : _GEN4739;
wire  _GEN4768 = io_x[18] ? _GEN4767 : _GEN4720;
wire  _GEN4769 = io_x[25] ? _GEN4768 : _GEN4690;
wire  _GEN4770 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4771 = io_x[30] ? _GEN3304 : _GEN4770;
wire  _GEN4772 = io_x[26] ? _GEN4771 : _GEN3306;
wire  _GEN4773 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN4774 = io_x[73] ? _GEN4773 : _GEN4772;
wire  _GEN4775 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4776 = io_x[30] ? _GEN4775 : _GEN3303;
wire  _GEN4777 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4778 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4779 = io_x[30] ? _GEN4778 : _GEN4777;
wire  _GEN4780 = io_x[26] ? _GEN4779 : _GEN4776;
wire  _GEN4781 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4782 = io_x[30] ? _GEN4781 : _GEN3304;
wire  _GEN4783 = io_x[26] ? _GEN4782 : _GEN3311;
wire  _GEN4784 = io_x[73] ? _GEN4783 : _GEN4780;
wire  _GEN4785 = io_x[33] ? _GEN4784 : _GEN4774;
wire  _GEN4786 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4787 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4788 = io_x[30] ? _GEN4787 : _GEN4786;
wire  _GEN4789 = io_x[26] ? _GEN4788 : _GEN3306;
wire  _GEN4790 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4791 = io_x[30] ? _GEN4790 : _GEN3304;
wire  _GEN4792 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4793 = io_x[30] ? _GEN4792 : _GEN3303;
wire  _GEN4794 = io_x[26] ? _GEN4793 : _GEN4791;
wire  _GEN4795 = io_x[73] ? _GEN4794 : _GEN4789;
wire  _GEN4796 = io_x[33] ? _GEN4795 : _GEN3302;
wire  _GEN4797 = io_x[28] ? _GEN4796 : _GEN4785;
wire  _GEN4798 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4799 = io_x[30] ? _GEN3303 : _GEN4798;
wire  _GEN4800 = io_x[26] ? _GEN4799 : _GEN3306;
wire  _GEN4801 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4802 = io_x[30] ? _GEN3304 : _GEN4801;
wire  _GEN4803 = io_x[26] ? _GEN4802 : _GEN3311;
wire  _GEN4804 = io_x[73] ? _GEN4803 : _GEN4800;
wire  _GEN4805 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4806 = io_x[30] ? _GEN4805 : _GEN3303;
wire  _GEN4807 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4808 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4809 = io_x[30] ? _GEN4808 : _GEN4807;
wire  _GEN4810 = io_x[26] ? _GEN4809 : _GEN4806;
wire  _GEN4811 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4812 = io_x[26] ? _GEN3311 : _GEN4811;
wire  _GEN4813 = io_x[73] ? _GEN4812 : _GEN4810;
wire  _GEN4814 = io_x[33] ? _GEN4813 : _GEN4804;
wire  _GEN4815 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4816 = io_x[30] ? _GEN4815 : _GEN3303;
wire  _GEN4817 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4818 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4819 = io_x[30] ? _GEN4818 : _GEN4817;
wire  _GEN4820 = io_x[26] ? _GEN4819 : _GEN4816;
wire  _GEN4821 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4822 = io_x[30] ? _GEN4821 : _GEN3304;
wire  _GEN4823 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4824 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4825 = io_x[30] ? _GEN4824 : _GEN4823;
wire  _GEN4826 = io_x[26] ? _GEN4825 : _GEN4822;
wire  _GEN4827 = io_x[73] ? _GEN4826 : _GEN4820;
wire  _GEN4828 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4829 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4830 = io_x[30] ? _GEN4829 : _GEN4828;
wire  _GEN4831 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4832 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4833 = io_x[30] ? _GEN4832 : _GEN4831;
wire  _GEN4834 = io_x[26] ? _GEN4833 : _GEN4830;
wire  _GEN4835 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4836 = io_x[30] ? _GEN4835 : _GEN3304;
wire  _GEN4837 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4838 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4839 = io_x[30] ? _GEN4838 : _GEN4837;
wire  _GEN4840 = io_x[26] ? _GEN4839 : _GEN4836;
wire  _GEN4841 = io_x[73] ? _GEN4840 : _GEN4834;
wire  _GEN4842 = io_x[33] ? _GEN4841 : _GEN4827;
wire  _GEN4843 = io_x[28] ? _GEN4842 : _GEN4814;
wire  _GEN4844 = io_x[18] ? _GEN4843 : _GEN4797;
wire  _GEN4845 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4846 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4847 = io_x[30] ? _GEN3303 : _GEN4846;
wire  _GEN4848 = io_x[26] ? _GEN4847 : _GEN4845;
wire  _GEN4849 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4850 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4851 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4852 = io_x[30] ? _GEN4851 : _GEN4850;
wire  _GEN4853 = io_x[26] ? _GEN4852 : _GEN4849;
wire  _GEN4854 = io_x[73] ? _GEN4853 : _GEN4848;
wire  _GEN4855 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4856 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4857 = io_x[30] ? _GEN4856 : _GEN4855;
wire  _GEN4858 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4859 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4860 = io_x[30] ? _GEN4859 : _GEN4858;
wire  _GEN4861 = io_x[26] ? _GEN4860 : _GEN4857;
wire  _GEN4862 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4863 = io_x[30] ? _GEN3304 : _GEN4862;
wire  _GEN4864 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4865 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4866 = io_x[30] ? _GEN4865 : _GEN4864;
wire  _GEN4867 = io_x[26] ? _GEN4866 : _GEN4863;
wire  _GEN4868 = io_x[73] ? _GEN4867 : _GEN4861;
wire  _GEN4869 = io_x[33] ? _GEN4868 : _GEN4854;
wire  _GEN4870 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4871 = io_x[30] ? _GEN4870 : _GEN3303;
wire  _GEN4872 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4873 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4874 = io_x[30] ? _GEN4873 : _GEN4872;
wire  _GEN4875 = io_x[26] ? _GEN4874 : _GEN4871;
wire  _GEN4876 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4877 = io_x[30] ? _GEN3304 : _GEN4876;
wire  _GEN4878 = io_x[26] ? _GEN4877 : _GEN3311;
wire  _GEN4879 = io_x[73] ? _GEN4878 : _GEN4875;
wire  _GEN4880 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4881 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4882 = io_x[30] ? _GEN4881 : _GEN4880;
wire  _GEN4883 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4884 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4885 = io_x[30] ? _GEN4884 : _GEN4883;
wire  _GEN4886 = io_x[26] ? _GEN4885 : _GEN4882;
wire  _GEN4887 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4888 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4889 = io_x[30] ? _GEN4888 : _GEN4887;
wire  _GEN4890 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4891 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4892 = io_x[30] ? _GEN4891 : _GEN4890;
wire  _GEN4893 = io_x[26] ? _GEN4892 : _GEN4889;
wire  _GEN4894 = io_x[73] ? _GEN4893 : _GEN4886;
wire  _GEN4895 = io_x[33] ? _GEN4894 : _GEN4879;
wire  _GEN4896 = io_x[28] ? _GEN4895 : _GEN4869;
wire  _GEN4897 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4898 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4899 = io_x[30] ? _GEN4898 : _GEN4897;
wire  _GEN4900 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4901 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4902 = io_x[30] ? _GEN4901 : _GEN4900;
wire  _GEN4903 = io_x[26] ? _GEN4902 : _GEN4899;
wire  _GEN4904 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4905 = io_x[30] ? _GEN3303 : _GEN4904;
wire  _GEN4906 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4907 = io_x[30] ? _GEN4906 : _GEN3304;
wire  _GEN4908 = io_x[26] ? _GEN4907 : _GEN4905;
wire  _GEN4909 = io_x[73] ? _GEN4908 : _GEN4903;
wire  _GEN4910 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4911 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4912 = io_x[30] ? _GEN4911 : _GEN4910;
wire  _GEN4913 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4914 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4915 = io_x[30] ? _GEN4914 : _GEN4913;
wire  _GEN4916 = io_x[26] ? _GEN4915 : _GEN4912;
wire  _GEN4917 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4918 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4919 = io_x[30] ? _GEN4918 : _GEN4917;
wire  _GEN4920 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4921 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4922 = io_x[30] ? _GEN4921 : _GEN4920;
wire  _GEN4923 = io_x[26] ? _GEN4922 : _GEN4919;
wire  _GEN4924 = io_x[73] ? _GEN4923 : _GEN4916;
wire  _GEN4925 = io_x[33] ? _GEN4924 : _GEN4909;
wire  _GEN4926 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4927 = io_x[30] ? _GEN4926 : _GEN3304;
wire  _GEN4928 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4929 = io_x[30] ? _GEN4928 : _GEN3304;
wire  _GEN4930 = io_x[26] ? _GEN4929 : _GEN4927;
wire  _GEN4931 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4932 = io_x[30] ? _GEN4931 : _GEN3304;
wire  _GEN4933 = io_x[26] ? _GEN4932 : _GEN3306;
wire  _GEN4934 = io_x[73] ? _GEN4933 : _GEN4930;
wire  _GEN4935 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4936 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4937 = io_x[30] ? _GEN4936 : _GEN4935;
wire  _GEN4938 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4939 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4940 = io_x[30] ? _GEN4939 : _GEN4938;
wire  _GEN4941 = io_x[26] ? _GEN4940 : _GEN4937;
wire  _GEN4942 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4943 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4944 = io_x[30] ? _GEN4943 : _GEN4942;
wire  _GEN4945 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4946 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4947 = io_x[30] ? _GEN4946 : _GEN4945;
wire  _GEN4948 = io_x[26] ? _GEN4947 : _GEN4944;
wire  _GEN4949 = io_x[73] ? _GEN4948 : _GEN4941;
wire  _GEN4950 = io_x[33] ? _GEN4949 : _GEN4934;
wire  _GEN4951 = io_x[28] ? _GEN4950 : _GEN4925;
wire  _GEN4952 = io_x[18] ? _GEN4951 : _GEN4896;
wire  _GEN4953 = io_x[25] ? _GEN4952 : _GEN4844;
wire  _GEN4954 = io_x[29] ? _GEN4953 : _GEN4769;
wire  _GEN4955 = io_x[23] ? _GEN4954 : _GEN4639;
wire  _GEN4956 = io_x[31] ? _GEN4955 : _GEN4427;
wire  _GEN4957 = io_x[19] ? _GEN4956 : _GEN4031;
wire  _GEN4958 = io_x[73] ? _GEN3308 : _GEN3324;
wire  _GEN4959 = io_x[33] ? _GEN4958 : _GEN3302;
wire  _GEN4960 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4961 = io_x[26] ? _GEN3311 : _GEN4960;
wire  _GEN4962 = io_x[73] ? _GEN4961 : _GEN3324;
wire  _GEN4963 = io_x[73] ? _GEN3308 : _GEN3324;
wire  _GEN4964 = io_x[33] ? _GEN4963 : _GEN4962;
wire  _GEN4965 = io_x[28] ? _GEN4964 : _GEN4959;
wire  _GEN4966 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN4967 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4968 = io_x[30] ? _GEN4967 : _GEN3304;
wire  _GEN4969 = io_x[26] ? _GEN4968 : _GEN3306;
wire  _GEN4970 = io_x[73] ? _GEN4969 : _GEN4966;
wire  _GEN4971 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN4972 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4973 = io_x[30] ? _GEN4972 : _GEN3304;
wire  _GEN4974 = io_x[26] ? _GEN4973 : _GEN4971;
wire  _GEN4975 = io_x[73] ? _GEN4974 : _GEN3308;
wire  _GEN4976 = io_x[33] ? _GEN4975 : _GEN4970;
wire  _GEN4977 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4978 = io_x[30] ? _GEN4977 : _GEN3304;
wire  _GEN4979 = io_x[26] ? _GEN4978 : _GEN3311;
wire  _GEN4980 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN4981 = io_x[73] ? _GEN4980 : _GEN4979;
wire  _GEN4982 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN4983 = io_x[30] ? _GEN4982 : _GEN3304;
wire  _GEN4984 = io_x[26] ? _GEN4983 : _GEN3311;
wire  _GEN4985 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN4986 = io_x[73] ? _GEN4985 : _GEN4984;
wire  _GEN4987 = io_x[33] ? _GEN4986 : _GEN4981;
wire  _GEN4988 = io_x[28] ? _GEN4987 : _GEN4976;
wire  _GEN4989 = io_x[18] ? _GEN4988 : _GEN4965;
wire  _GEN4990 = io_x[73] ? _GEN3324 : _GEN3308;
wire  _GEN4991 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN4992 = io_x[30] ? _GEN4991 : _GEN3304;
wire  _GEN4993 = io_x[26] ? _GEN4992 : _GEN3306;
wire  _GEN4994 = io_x[73] ? _GEN4993 : _GEN3308;
wire  _GEN4995 = io_x[33] ? _GEN4994 : _GEN4990;
wire  _GEN4996 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN4997 = io_x[26] ? _GEN4996 : _GEN3311;
wire  _GEN4998 = io_x[73] ? _GEN4997 : _GEN3308;
wire  _GEN4999 = io_x[33] ? _GEN4998 : _GEN3371;
wire  _GEN5000 = io_x[28] ? _GEN4999 : _GEN4995;
wire  _GEN5001 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5002 = io_x[73] ? _GEN3324 : _GEN5001;
wire  _GEN5003 = io_x[33] ? _GEN5002 : _GEN3371;
wire  _GEN5004 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5005 = io_x[30] ? _GEN3304 : _GEN5004;
wire  _GEN5006 = io_x[26] ? _GEN5005 : _GEN3311;
wire  _GEN5007 = io_x[73] ? _GEN3308 : _GEN5006;
wire  _GEN5008 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5009 = io_x[30] ? _GEN5008 : _GEN3304;
wire  _GEN5010 = io_x[26] ? _GEN5009 : _GEN3306;
wire  _GEN5011 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5012 = io_x[30] ? _GEN5011 : _GEN3303;
wire  _GEN5013 = io_x[26] ? _GEN5012 : _GEN3311;
wire  _GEN5014 = io_x[73] ? _GEN5013 : _GEN5010;
wire  _GEN5015 = io_x[33] ? _GEN5014 : _GEN5007;
wire  _GEN5016 = io_x[28] ? _GEN5015 : _GEN5003;
wire  _GEN5017 = io_x[18] ? _GEN5016 : _GEN5000;
wire  _GEN5018 = io_x[25] ? _GEN5017 : _GEN4989;
wire  _GEN5019 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5020 = io_x[30] ? _GEN5019 : _GEN3304;
wire  _GEN5021 = io_x[26] ? _GEN3306 : _GEN5020;
wire  _GEN5022 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5023 = io_x[73] ? _GEN5022 : _GEN5021;
wire  _GEN5024 = io_x[33] ? _GEN5023 : _GEN3302;
wire  _GEN5025 = io_x[28] ? _GEN4086 : _GEN5024;
wire  _GEN5026 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5027 = io_x[26] ? _GEN5026 : _GEN3306;
wire  _GEN5028 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5029 = io_x[26] ? _GEN5028 : _GEN3306;
wire  _GEN5030 = io_x[73] ? _GEN5029 : _GEN5027;
wire  _GEN5031 = io_x[33] ? _GEN5030 : _GEN3371;
wire  _GEN5032 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5033 = io_x[26] ? _GEN5032 : _GEN3306;
wire  _GEN5034 = io_x[73] ? _GEN3308 : _GEN5033;
wire  _GEN5035 = io_x[33] ? _GEN3302 : _GEN5034;
wire  _GEN5036 = io_x[28] ? _GEN5035 : _GEN5031;
wire  _GEN5037 = io_x[18] ? _GEN5036 : _GEN5025;
wire  _GEN5038 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5039 = io_x[26] ? _GEN5038 : _GEN3306;
wire  _GEN5040 = io_x[73] ? _GEN3324 : _GEN5039;
wire  _GEN5041 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5042 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5043 = io_x[73] ? _GEN5042 : _GEN5041;
wire  _GEN5044 = io_x[33] ? _GEN5043 : _GEN5040;
wire  _GEN5045 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5046 = io_x[73] ? _GEN3308 : _GEN5045;
wire  _GEN5047 = io_x[33] ? _GEN5046 : _GEN3302;
wire  _GEN5048 = io_x[28] ? _GEN5047 : _GEN5044;
wire  _GEN5049 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5050 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5051 = io_x[30] ? _GEN5050 : _GEN5049;
wire  _GEN5052 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5053 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5054 = io_x[30] ? _GEN5053 : _GEN5052;
wire  _GEN5055 = io_x[26] ? _GEN5054 : _GEN5051;
wire  _GEN5056 = io_x[73] ? _GEN3324 : _GEN5055;
wire  _GEN5057 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5058 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5059 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5060 = io_x[30] ? _GEN5059 : _GEN5058;
wire  _GEN5061 = io_x[26] ? _GEN5060 : _GEN5057;
wire  _GEN5062 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5063 = io_x[30] ? _GEN3304 : _GEN5062;
wire  _GEN5064 = io_x[26] ? _GEN5063 : _GEN3311;
wire  _GEN5065 = io_x[73] ? _GEN5064 : _GEN5061;
wire  _GEN5066 = io_x[33] ? _GEN5065 : _GEN5056;
wire  _GEN5067 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5068 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5069 = io_x[73] ? _GEN5068 : _GEN5067;
wire  _GEN5070 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5071 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5072 = io_x[30] ? _GEN3304 : _GEN5071;
wire  _GEN5073 = io_x[26] ? _GEN5072 : _GEN3311;
wire  _GEN5074 = io_x[73] ? _GEN5073 : _GEN5070;
wire  _GEN5075 = io_x[33] ? _GEN5074 : _GEN5069;
wire  _GEN5076 = io_x[28] ? _GEN5075 : _GEN5066;
wire  _GEN5077 = io_x[18] ? _GEN5076 : _GEN5048;
wire  _GEN5078 = io_x[25] ? _GEN5077 : _GEN5037;
wire  _GEN5079 = io_x[29] ? _GEN5078 : _GEN5018;
wire  _GEN5080 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5081 = io_x[30] ? _GEN5080 : _GEN3304;
wire  _GEN5082 = io_x[26] ? _GEN5081 : _GEN3306;
wire  _GEN5083 = io_x[73] ? _GEN3324 : _GEN5082;
wire  _GEN5084 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5085 = io_x[26] ? _GEN5084 : _GEN3311;
wire  _GEN5086 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5087 = io_x[73] ? _GEN5086 : _GEN5085;
wire  _GEN5088 = io_x[33] ? _GEN5087 : _GEN5083;
wire  _GEN5089 = io_x[28] ? _GEN5088 : _GEN3498;
wire  _GEN5090 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5091 = io_x[30] ? _GEN5090 : _GEN3303;
wire  _GEN5092 = io_x[26] ? _GEN3311 : _GEN5091;
wire  _GEN5093 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5094 = io_x[73] ? _GEN5093 : _GEN5092;
wire  _GEN5095 = io_x[33] ? _GEN5094 : _GEN3371;
wire  _GEN5096 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5097 = io_x[30] ? _GEN5096 : _GEN3304;
wire  _GEN5098 = io_x[26] ? _GEN5097 : _GEN3306;
wire  _GEN5099 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5100 = io_x[30] ? _GEN5099 : _GEN3304;
wire  _GEN5101 = io_x[26] ? _GEN5100 : _GEN3306;
wire  _GEN5102 = io_x[73] ? _GEN5101 : _GEN5098;
wire  _GEN5103 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5104 = io_x[30] ? _GEN5103 : _GEN3304;
wire  _GEN5105 = io_x[26] ? _GEN5104 : _GEN3311;
wire  _GEN5106 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5107 = io_x[30] ? _GEN5106 : _GEN3304;
wire  _GEN5108 = io_x[26] ? _GEN5107 : _GEN3306;
wire  _GEN5109 = io_x[73] ? _GEN5108 : _GEN5105;
wire  _GEN5110 = io_x[33] ? _GEN5109 : _GEN5102;
wire  _GEN5111 = io_x[28] ? _GEN5110 : _GEN5095;
wire  _GEN5112 = io_x[18] ? _GEN5111 : _GEN5089;
wire  _GEN5113 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5114 = io_x[26] ? _GEN3311 : _GEN5113;
wire  _GEN5115 = io_x[73] ? _GEN5114 : _GEN3324;
wire  _GEN5116 = io_x[33] ? _GEN5115 : _GEN3371;
wire  _GEN5117 = io_x[28] ? _GEN5116 : _GEN4086;
wire  _GEN5118 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5119 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5120 = io_x[30] ? _GEN5119 : _GEN3304;
wire  _GEN5121 = io_x[26] ? _GEN5120 : _GEN5118;
wire  _GEN5122 = io_x[73] ? _GEN3308 : _GEN5121;
wire  _GEN5123 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5124 = io_x[73] ? _GEN3308 : _GEN5123;
wire  _GEN5125 = io_x[33] ? _GEN5124 : _GEN5122;
wire  _GEN5126 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5127 = io_x[30] ? _GEN5126 : _GEN3303;
wire  _GEN5128 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5129 = io_x[30] ? _GEN5128 : _GEN3304;
wire  _GEN5130 = io_x[26] ? _GEN5129 : _GEN5127;
wire  _GEN5131 = io_x[73] ? _GEN3308 : _GEN5130;
wire  _GEN5132 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5133 = io_x[30] ? _GEN5132 : _GEN3303;
wire  _GEN5134 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5135 = io_x[30] ? _GEN5134 : _GEN3304;
wire  _GEN5136 = io_x[26] ? _GEN5135 : _GEN5133;
wire  _GEN5137 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5138 = io_x[30] ? _GEN5137 : _GEN3303;
wire  _GEN5139 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5140 = io_x[30] ? _GEN5139 : _GEN3304;
wire  _GEN5141 = io_x[26] ? _GEN5140 : _GEN5138;
wire  _GEN5142 = io_x[73] ? _GEN5141 : _GEN5136;
wire  _GEN5143 = io_x[33] ? _GEN5142 : _GEN5131;
wire  _GEN5144 = io_x[28] ? _GEN5143 : _GEN5125;
wire  _GEN5145 = io_x[18] ? _GEN5144 : _GEN5117;
wire  _GEN5146 = io_x[25] ? _GEN5145 : _GEN5112;
wire  _GEN5147 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5148 = io_x[30] ? _GEN3304 : _GEN5147;
wire  _GEN5149 = io_x[26] ? _GEN5148 : _GEN3306;
wire  _GEN5150 = io_x[73] ? _GEN3324 : _GEN5149;
wire  _GEN5151 = io_x[33] ? _GEN5150 : _GEN3371;
wire  _GEN5152 = io_x[28] ? _GEN3498 : _GEN5151;
wire  _GEN5153 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5154 = io_x[30] ? _GEN3304 : _GEN5153;
wire  _GEN5155 = io_x[26] ? _GEN5154 : _GEN3306;
wire  _GEN5156 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5157 = io_x[26] ? _GEN5156 : _GEN3306;
wire  _GEN5158 = io_x[73] ? _GEN5157 : _GEN5155;
wire  _GEN5159 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5160 = io_x[30] ? _GEN3304 : _GEN5159;
wire  _GEN5161 = io_x[26] ? _GEN5160 : _GEN3306;
wire  _GEN5162 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5163 = io_x[30] ? _GEN3304 : _GEN5162;
wire  _GEN5164 = io_x[26] ? _GEN5163 : _GEN3306;
wire  _GEN5165 = io_x[73] ? _GEN5164 : _GEN5161;
wire  _GEN5166 = io_x[33] ? _GEN5165 : _GEN5158;
wire  _GEN5167 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5168 = io_x[30] ? _GEN5167 : _GEN3304;
wire  _GEN5169 = io_x[26] ? _GEN3311 : _GEN5168;
wire  _GEN5170 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5171 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5172 = io_x[30] ? _GEN5171 : _GEN3304;
wire  _GEN5173 = io_x[26] ? _GEN5172 : _GEN5170;
wire  _GEN5174 = io_x[73] ? _GEN5173 : _GEN5169;
wire  _GEN5175 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5176 = io_x[30] ? _GEN3304 : _GEN5175;
wire  _GEN5177 = io_x[26] ? _GEN3311 : _GEN5176;
wire  _GEN5178 = io_x[73] ? _GEN5177 : _GEN3308;
wire  _GEN5179 = io_x[33] ? _GEN5178 : _GEN5174;
wire  _GEN5180 = io_x[28] ? _GEN5179 : _GEN5166;
wire  _GEN5181 = io_x[18] ? _GEN5180 : _GEN5152;
wire  _GEN5182 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5183 = io_x[30] ? _GEN5182 : _GEN3304;
wire  _GEN5184 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5185 = io_x[30] ? _GEN5184 : _GEN3304;
wire  _GEN5186 = io_x[26] ? _GEN5185 : _GEN5183;
wire  _GEN5187 = io_x[73] ? _GEN3324 : _GEN5186;
wire  _GEN5188 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5189 = io_x[30] ? _GEN5188 : _GEN3304;
wire  _GEN5190 = io_x[26] ? _GEN3306 : _GEN5189;
wire  _GEN5191 = io_x[73] ? _GEN3324 : _GEN5190;
wire  _GEN5192 = io_x[33] ? _GEN5191 : _GEN5187;
wire  _GEN5193 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5194 = io_x[26] ? _GEN3306 : _GEN5193;
wire  _GEN5195 = io_x[73] ? _GEN3308 : _GEN5194;
wire  _GEN5196 = io_x[73] ? _GEN3324 : _GEN3308;
wire  _GEN5197 = io_x[33] ? _GEN5196 : _GEN5195;
wire  _GEN5198 = io_x[28] ? _GEN5197 : _GEN5192;
wire  _GEN5199 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5200 = io_x[26] ? _GEN3306 : _GEN5199;
wire  _GEN5201 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5202 = io_x[30] ? _GEN5201 : _GEN3304;
wire  _GEN5203 = io_x[26] ? _GEN3306 : _GEN5202;
wire  _GEN5204 = io_x[73] ? _GEN5203 : _GEN5200;
wire  _GEN5205 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5206 = io_x[30] ? _GEN5205 : _GEN3304;
wire  _GEN5207 = io_x[26] ? _GEN3306 : _GEN5206;
wire  _GEN5208 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5209 = io_x[30] ? _GEN5208 : _GEN3304;
wire  _GEN5210 = io_x[26] ? _GEN3306 : _GEN5209;
wire  _GEN5211 = io_x[73] ? _GEN5210 : _GEN5207;
wire  _GEN5212 = io_x[33] ? _GEN5211 : _GEN5204;
wire  _GEN5213 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5214 = io_x[30] ? _GEN5213 : _GEN3304;
wire  _GEN5215 = io_x[26] ? _GEN5214 : _GEN3311;
wire  _GEN5216 = io_x[73] ? _GEN3324 : _GEN5215;
wire  _GEN5217 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5218 = io_x[30] ? _GEN5217 : _GEN3303;
wire  _GEN5219 = io_x[26] ? _GEN5218 : _GEN3311;
wire  _GEN5220 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5221 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5222 = io_x[30] ? _GEN5221 : _GEN3304;
wire  _GEN5223 = io_x[26] ? _GEN5222 : _GEN5220;
wire  _GEN5224 = io_x[73] ? _GEN5223 : _GEN5219;
wire  _GEN5225 = io_x[33] ? _GEN5224 : _GEN5216;
wire  _GEN5226 = io_x[28] ? _GEN5225 : _GEN5212;
wire  _GEN5227 = io_x[18] ? _GEN5226 : _GEN5198;
wire  _GEN5228 = io_x[25] ? _GEN5227 : _GEN5181;
wire  _GEN5229 = io_x[29] ? _GEN5228 : _GEN5146;
wire  _GEN5230 = io_x[23] ? _GEN5229 : _GEN5079;
wire  _GEN5231 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5232 = io_x[30] ? _GEN3304 : _GEN5231;
wire  _GEN5233 = io_x[26] ? _GEN5232 : _GEN3306;
wire  _GEN5234 = io_x[73] ? _GEN5233 : _GEN3308;
wire  _GEN5235 = io_x[33] ? _GEN5234 : _GEN3302;
wire  _GEN5236 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5237 = io_x[26] ? _GEN5236 : _GEN3306;
wire  _GEN5238 = io_x[73] ? _GEN3308 : _GEN5237;
wire  _GEN5239 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5240 = io_x[26] ? _GEN5239 : _GEN3306;
wire  _GEN5241 = io_x[73] ? _GEN3308 : _GEN5240;
wire  _GEN5242 = io_x[33] ? _GEN5241 : _GEN5238;
wire  _GEN5243 = io_x[28] ? _GEN5242 : _GEN5235;
wire  _GEN5244 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5245 = io_x[26] ? _GEN5244 : _GEN3306;
wire  _GEN5246 = io_x[73] ? _GEN3308 : _GEN5245;
wire  _GEN5247 = io_x[33] ? _GEN5246 : _GEN3302;
wire  _GEN5248 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5249 = io_x[26] ? _GEN5248 : _GEN3306;
wire  _GEN5250 = io_x[73] ? _GEN5249 : _GEN3324;
wire  _GEN5251 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5252 = io_x[30] ? _GEN5251 : _GEN3303;
wire  _GEN5253 = io_x[26] ? _GEN5252 : _GEN3306;
wire  _GEN5254 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5255 = io_x[30] ? _GEN5254 : _GEN3303;
wire  _GEN5256 = io_x[26] ? _GEN5255 : _GEN3306;
wire  _GEN5257 = io_x[73] ? _GEN5256 : _GEN5253;
wire  _GEN5258 = io_x[33] ? _GEN5257 : _GEN5250;
wire  _GEN5259 = io_x[28] ? _GEN5258 : _GEN5247;
wire  _GEN5260 = io_x[18] ? _GEN5259 : _GEN5243;
wire  _GEN5261 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5262 = io_x[30] ? _GEN5261 : _GEN3304;
wire  _GEN5263 = io_x[26] ? _GEN5262 : _GEN3306;
wire  _GEN5264 = io_x[73] ? _GEN5263 : _GEN3308;
wire  _GEN5265 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5266 = io_x[30] ? _GEN5265 : _GEN3303;
wire  _GEN5267 = io_x[26] ? _GEN5266 : _GEN3306;
wire  _GEN5268 = io_x[73] ? _GEN5267 : _GEN3308;
wire  _GEN5269 = io_x[33] ? _GEN5268 : _GEN5264;
wire  _GEN5270 = io_x[28] ? _GEN4086 : _GEN5269;
wire  _GEN5271 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5272 = io_x[30] ? _GEN5271 : _GEN3303;
wire  _GEN5273 = io_x[26] ? _GEN3306 : _GEN5272;
wire  _GEN5274 = io_x[73] ? _GEN3324 : _GEN5273;
wire  _GEN5275 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5276 = io_x[73] ? _GEN3308 : _GEN5275;
wire  _GEN5277 = io_x[33] ? _GEN5276 : _GEN5274;
wire  _GEN5278 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5279 = io_x[30] ? _GEN3304 : _GEN5278;
wire  _GEN5280 = io_x[26] ? _GEN3311 : _GEN5279;
wire  _GEN5281 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5282 = io_x[30] ? _GEN3303 : _GEN5281;
wire  _GEN5283 = io_x[26] ? _GEN3306 : _GEN5282;
wire  _GEN5284 = io_x[73] ? _GEN5283 : _GEN5280;
wire  _GEN5285 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5286 = io_x[30] ? _GEN3303 : _GEN5285;
wire  _GEN5287 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5288 = io_x[30] ? _GEN5287 : _GEN3303;
wire  _GEN5289 = io_x[26] ? _GEN5288 : _GEN5286;
wire  _GEN5290 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5291 = io_x[30] ? _GEN5290 : _GEN3304;
wire  _GEN5292 = io_x[26] ? _GEN5291 : _GEN3311;
wire  _GEN5293 = io_x[73] ? _GEN5292 : _GEN5289;
wire  _GEN5294 = io_x[33] ? _GEN5293 : _GEN5284;
wire  _GEN5295 = io_x[28] ? _GEN5294 : _GEN5277;
wire  _GEN5296 = io_x[18] ? _GEN5295 : _GEN5270;
wire  _GEN5297 = io_x[25] ? _GEN5296 : _GEN5260;
wire  _GEN5298 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5299 = io_x[26] ? _GEN5298 : _GEN3311;
wire  _GEN5300 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5301 = io_x[30] ? _GEN5300 : _GEN3304;
wire  _GEN5302 = io_x[26] ? _GEN5301 : _GEN3306;
wire  _GEN5303 = io_x[73] ? _GEN5302 : _GEN5299;
wire  _GEN5304 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5305 = io_x[26] ? _GEN5304 : _GEN3311;
wire  _GEN5306 = io_x[73] ? _GEN3308 : _GEN5305;
wire  _GEN5307 = io_x[33] ? _GEN5306 : _GEN5303;
wire  _GEN5308 = io_x[73] ? _GEN3324 : _GEN3308;
wire  _GEN5309 = io_x[33] ? _GEN3302 : _GEN5308;
wire  _GEN5310 = io_x[28] ? _GEN5309 : _GEN5307;
wire  _GEN5311 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5312 = io_x[26] ? _GEN5311 : _GEN3311;
wire  _GEN5313 = io_x[73] ? _GEN3308 : _GEN5312;
wire  _GEN5314 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5315 = io_x[30] ? _GEN5314 : _GEN3304;
wire  _GEN5316 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5317 = io_x[26] ? _GEN5316 : _GEN5315;
wire  _GEN5318 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5319 = io_x[30] ? _GEN5318 : _GEN3303;
wire  _GEN5320 = io_x[26] ? _GEN5319 : _GEN3306;
wire  _GEN5321 = io_x[73] ? _GEN5320 : _GEN5317;
wire  _GEN5322 = io_x[33] ? _GEN5321 : _GEN5313;
wire  _GEN5323 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5324 = io_x[30] ? _GEN3304 : _GEN5323;
wire  _GEN5325 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5326 = io_x[26] ? _GEN5325 : _GEN5324;
wire  _GEN5327 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5328 = io_x[73] ? _GEN5327 : _GEN5326;
wire  _GEN5329 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5330 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5331 = io_x[30] ? _GEN5330 : _GEN5329;
wire  _GEN5332 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5333 = io_x[26] ? _GEN5332 : _GEN5331;
wire  _GEN5334 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5335 = io_x[30] ? _GEN3304 : _GEN5334;
wire  _GEN5336 = io_x[26] ? _GEN3311 : _GEN5335;
wire  _GEN5337 = io_x[73] ? _GEN5336 : _GEN5333;
wire  _GEN5338 = io_x[33] ? _GEN5337 : _GEN5328;
wire  _GEN5339 = io_x[28] ? _GEN5338 : _GEN5322;
wire  _GEN5340 = io_x[18] ? _GEN5339 : _GEN5310;
wire  _GEN5341 = io_x[73] ? _GEN3324 : _GEN3308;
wire  _GEN5342 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5343 = io_x[30] ? _GEN5342 : _GEN3304;
wire  _GEN5344 = io_x[26] ? _GEN5343 : _GEN3306;
wire  _GEN5345 = io_x[73] ? _GEN3308 : _GEN5344;
wire  _GEN5346 = io_x[33] ? _GEN5345 : _GEN5341;
wire  _GEN5347 = io_x[73] ? _GEN3308 : _GEN3324;
wire  _GEN5348 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5349 = io_x[30] ? _GEN5348 : _GEN3303;
wire  _GEN5350 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5351 = io_x[30] ? _GEN5350 : _GEN3304;
wire  _GEN5352 = io_x[26] ? _GEN5351 : _GEN5349;
wire  _GEN5353 = io_x[73] ? _GEN5352 : _GEN3324;
wire  _GEN5354 = io_x[33] ? _GEN5353 : _GEN5347;
wire  _GEN5355 = io_x[28] ? _GEN5354 : _GEN5346;
wire  _GEN5356 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5357 = io_x[30] ? _GEN3303 : _GEN5356;
wire  _GEN5358 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5359 = io_x[30] ? _GEN5358 : _GEN3304;
wire  _GEN5360 = io_x[26] ? _GEN5359 : _GEN5357;
wire  _GEN5361 = io_x[73] ? _GEN3308 : _GEN5360;
wire  _GEN5362 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5363 = io_x[30] ? _GEN5362 : _GEN3304;
wire  _GEN5364 = io_x[26] ? _GEN5363 : _GEN3306;
wire  _GEN5365 = io_x[73] ? _GEN3324 : _GEN5364;
wire  _GEN5366 = io_x[33] ? _GEN5365 : _GEN5361;
wire  _GEN5367 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5368 = io_x[26] ? _GEN3306 : _GEN5367;
wire  _GEN5369 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5370 = io_x[73] ? _GEN5369 : _GEN5368;
wire  _GEN5371 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5372 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5373 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5374 = io_x[30] ? _GEN5373 : _GEN5372;
wire  _GEN5375 = io_x[26] ? _GEN5374 : _GEN5371;
wire  _GEN5376 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5377 = io_x[30] ? _GEN5376 : _GEN3304;
wire  _GEN5378 = io_x[26] ? _GEN5377 : _GEN3311;
wire  _GEN5379 = io_x[73] ? _GEN5378 : _GEN5375;
wire  _GEN5380 = io_x[33] ? _GEN5379 : _GEN5370;
wire  _GEN5381 = io_x[28] ? _GEN5380 : _GEN5366;
wire  _GEN5382 = io_x[18] ? _GEN5381 : _GEN5355;
wire  _GEN5383 = io_x[25] ? _GEN5382 : _GEN5340;
wire  _GEN5384 = io_x[29] ? _GEN5383 : _GEN5297;
wire  _GEN5385 = io_x[33] ? _GEN3371 : _GEN3302;
wire  _GEN5386 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5387 = io_x[30] ? _GEN5386 : _GEN3304;
wire  _GEN5388 = io_x[26] ? _GEN3306 : _GEN5387;
wire  _GEN5389 = io_x[73] ? _GEN3324 : _GEN5388;
wire  _GEN5390 = io_x[33] ? _GEN3302 : _GEN5389;
wire  _GEN5391 = io_x[28] ? _GEN5390 : _GEN5385;
wire  _GEN5392 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5393 = io_x[26] ? _GEN3306 : _GEN5392;
wire  _GEN5394 = io_x[73] ? _GEN3308 : _GEN5393;
wire  _GEN5395 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5396 = io_x[26] ? _GEN3306 : _GEN5395;
wire  _GEN5397 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5398 = io_x[30] ? _GEN5397 : _GEN3303;
wire  _GEN5399 = io_x[26] ? _GEN5398 : _GEN3311;
wire  _GEN5400 = io_x[73] ? _GEN5399 : _GEN5396;
wire  _GEN5401 = io_x[33] ? _GEN5400 : _GEN5394;
wire  _GEN5402 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5403 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5404 = io_x[30] ? _GEN5403 : _GEN5402;
wire  _GEN5405 = io_x[26] ? _GEN5404 : _GEN3306;
wire  _GEN5406 = io_x[73] ? _GEN5405 : _GEN3324;
wire  _GEN5407 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5408 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5409 = io_x[30] ? _GEN5408 : _GEN5407;
wire  _GEN5410 = io_x[26] ? _GEN5409 : _GEN3306;
wire  _GEN5411 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5412 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5413 = io_x[30] ? _GEN5412 : _GEN5411;
wire  _GEN5414 = io_x[26] ? _GEN5413 : _GEN3311;
wire  _GEN5415 = io_x[73] ? _GEN5414 : _GEN5410;
wire  _GEN5416 = io_x[33] ? _GEN5415 : _GEN5406;
wire  _GEN5417 = io_x[28] ? _GEN5416 : _GEN5401;
wire  _GEN5418 = io_x[18] ? _GEN5417 : _GEN5391;
wire  _GEN5419 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5420 = io_x[30] ? _GEN5419 : _GEN3303;
wire  _GEN5421 = io_x[26] ? _GEN5420 : _GEN3311;
wire  _GEN5422 = io_x[73] ? _GEN3324 : _GEN5421;
wire  _GEN5423 = io_x[33] ? _GEN5422 : _GEN3371;
wire  _GEN5424 = io_x[28] ? _GEN5423 : _GEN3498;
wire  _GEN5425 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5426 = io_x[73] ? _GEN3308 : _GEN5425;
wire  _GEN5427 = io_x[33] ? _GEN3302 : _GEN5426;
wire  _GEN5428 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5429 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5430 = io_x[30] ? _GEN5429 : _GEN5428;
wire  _GEN5431 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5432 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5433 = io_x[30] ? _GEN5432 : _GEN5431;
wire  _GEN5434 = io_x[26] ? _GEN5433 : _GEN5430;
wire  _GEN5435 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5436 = io_x[30] ? _GEN5435 : _GEN3304;
wire  _GEN5437 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5438 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5439 = io_x[30] ? _GEN5438 : _GEN5437;
wire  _GEN5440 = io_x[26] ? _GEN5439 : _GEN5436;
wire  _GEN5441 = io_x[73] ? _GEN5440 : _GEN5434;
wire  _GEN5442 = io_x[33] ? _GEN5441 : _GEN3302;
wire  _GEN5443 = io_x[28] ? _GEN5442 : _GEN5427;
wire  _GEN5444 = io_x[18] ? _GEN5443 : _GEN5424;
wire  _GEN5445 = io_x[25] ? _GEN5444 : _GEN5418;
wire  _GEN5446 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5447 = io_x[30] ? _GEN5446 : _GEN3304;
wire  _GEN5448 = io_x[26] ? _GEN5447 : _GEN3306;
wire  _GEN5449 = io_x[73] ? _GEN5448 : _GEN3308;
wire  _GEN5450 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5451 = io_x[30] ? _GEN5450 : _GEN3303;
wire  _GEN5452 = io_x[26] ? _GEN5451 : _GEN3306;
wire  _GEN5453 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5454 = io_x[30] ? _GEN5453 : _GEN3303;
wire  _GEN5455 = io_x[26] ? _GEN5454 : _GEN3306;
wire  _GEN5456 = io_x[73] ? _GEN5455 : _GEN5452;
wire  _GEN5457 = io_x[33] ? _GEN5456 : _GEN5449;
wire  _GEN5458 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5459 = io_x[26] ? _GEN5458 : _GEN3306;
wire  _GEN5460 = io_x[73] ? _GEN3324 : _GEN5459;
wire  _GEN5461 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5462 = io_x[30] ? _GEN3304 : _GEN5461;
wire  _GEN5463 = io_x[26] ? _GEN5462 : _GEN3306;
wire  _GEN5464 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5465 = io_x[30] ? _GEN3304 : _GEN5464;
wire  _GEN5466 = io_x[26] ? _GEN5465 : _GEN3306;
wire  _GEN5467 = io_x[73] ? _GEN5466 : _GEN5463;
wire  _GEN5468 = io_x[33] ? _GEN5467 : _GEN5460;
wire  _GEN5469 = io_x[28] ? _GEN5468 : _GEN5457;
wire  _GEN5470 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5471 = io_x[26] ? _GEN5470 : _GEN3306;
wire  _GEN5472 = io_x[73] ? _GEN3324 : _GEN5471;
wire  _GEN5473 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5474 = io_x[30] ? _GEN5473 : _GEN3304;
wire  _GEN5475 = io_x[26] ? _GEN5474 : _GEN3311;
wire  _GEN5476 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5477 = io_x[30] ? _GEN5476 : _GEN3303;
wire  _GEN5478 = io_x[26] ? _GEN5477 : _GEN3306;
wire  _GEN5479 = io_x[73] ? _GEN5478 : _GEN5475;
wire  _GEN5480 = io_x[33] ? _GEN5479 : _GEN5472;
wire  _GEN5481 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5482 = io_x[30] ? _GEN3304 : _GEN5481;
wire  _GEN5483 = io_x[26] ? _GEN5482 : _GEN3306;
wire  _GEN5484 = io_x[73] ? _GEN3324 : _GEN5483;
wire  _GEN5485 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5486 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5487 = io_x[30] ? _GEN5486 : _GEN5485;
wire  _GEN5488 = io_x[26] ? _GEN5487 : _GEN3306;
wire  _GEN5489 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5490 = io_x[30] ? _GEN3303 : _GEN5489;
wire  _GEN5491 = io_x[26] ? _GEN5490 : _GEN3306;
wire  _GEN5492 = io_x[73] ? _GEN5491 : _GEN5488;
wire  _GEN5493 = io_x[33] ? _GEN5492 : _GEN5484;
wire  _GEN5494 = io_x[28] ? _GEN5493 : _GEN5480;
wire  _GEN5495 = io_x[18] ? _GEN5494 : _GEN5469;
wire  _GEN5496 = io_x[73] ? _GEN3324 : _GEN3308;
wire  _GEN5497 = io_x[73] ? _GEN3324 : _GEN3308;
wire  _GEN5498 = io_x[33] ? _GEN5497 : _GEN5496;
wire  _GEN5499 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5500 = io_x[30] ? _GEN5499 : _GEN3304;
wire  _GEN5501 = io_x[26] ? _GEN5500 : _GEN3306;
wire  _GEN5502 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5503 = io_x[30] ? _GEN5502 : _GEN3304;
wire  _GEN5504 = io_x[26] ? _GEN5503 : _GEN3311;
wire  _GEN5505 = io_x[73] ? _GEN5504 : _GEN5501;
wire  _GEN5506 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5507 = io_x[26] ? _GEN3306 : _GEN5506;
wire  _GEN5508 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5509 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5510 = io_x[30] ? _GEN5509 : _GEN3304;
wire  _GEN5511 = io_x[26] ? _GEN5510 : _GEN5508;
wire  _GEN5512 = io_x[73] ? _GEN5511 : _GEN5507;
wire  _GEN5513 = io_x[33] ? _GEN5512 : _GEN5505;
wire  _GEN5514 = io_x[28] ? _GEN5513 : _GEN5498;
wire  _GEN5515 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5516 = io_x[30] ? _GEN3304 : _GEN5515;
wire  _GEN5517 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5518 = io_x[26] ? _GEN5517 : _GEN5516;
wire  _GEN5519 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5520 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5521 = io_x[30] ? _GEN5520 : _GEN5519;
wire  _GEN5522 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5523 = io_x[26] ? _GEN5522 : _GEN5521;
wire  _GEN5524 = io_x[73] ? _GEN5523 : _GEN5518;
wire  _GEN5525 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5526 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5527 = io_x[30] ? _GEN5526 : _GEN5525;
wire  _GEN5528 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5529 = io_x[26] ? _GEN5528 : _GEN5527;
wire  _GEN5530 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5531 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5532 = io_x[30] ? _GEN5531 : _GEN5530;
wire  _GEN5533 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5534 = io_x[26] ? _GEN5533 : _GEN5532;
wire  _GEN5535 = io_x[73] ? _GEN5534 : _GEN5529;
wire  _GEN5536 = io_x[33] ? _GEN5535 : _GEN5524;
wire  _GEN5537 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5538 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5539 = io_x[30] ? _GEN5538 : _GEN5537;
wire  _GEN5540 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5541 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5542 = io_x[30] ? _GEN5541 : _GEN5540;
wire  _GEN5543 = io_x[26] ? _GEN5542 : _GEN5539;
wire  _GEN5544 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5545 = io_x[30] ? _GEN5544 : _GEN3304;
wire  _GEN5546 = io_x[26] ? _GEN5545 : _GEN3311;
wire  _GEN5547 = io_x[73] ? _GEN5546 : _GEN5543;
wire  _GEN5548 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5549 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5550 = io_x[30] ? _GEN5549 : _GEN5548;
wire  _GEN5551 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5552 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5553 = io_x[30] ? _GEN5552 : _GEN5551;
wire  _GEN5554 = io_x[26] ? _GEN5553 : _GEN5550;
wire  _GEN5555 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5556 = io_x[30] ? _GEN3303 : _GEN5555;
wire  _GEN5557 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5558 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5559 = io_x[30] ? _GEN5558 : _GEN5557;
wire  _GEN5560 = io_x[26] ? _GEN5559 : _GEN5556;
wire  _GEN5561 = io_x[73] ? _GEN5560 : _GEN5554;
wire  _GEN5562 = io_x[33] ? _GEN5561 : _GEN5547;
wire  _GEN5563 = io_x[28] ? _GEN5562 : _GEN5536;
wire  _GEN5564 = io_x[18] ? _GEN5563 : _GEN5514;
wire  _GEN5565 = io_x[25] ? _GEN5564 : _GEN5495;
wire  _GEN5566 = io_x[29] ? _GEN5565 : _GEN5445;
wire  _GEN5567 = io_x[23] ? _GEN5566 : _GEN5384;
wire  _GEN5568 = io_x[31] ? _GEN5567 : _GEN5230;
wire  _GEN5569 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5570 = io_x[73] ? _GEN3308 : _GEN5569;
wire  _GEN5571 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5572 = io_x[30] ? _GEN5571 : _GEN3303;
wire  _GEN5573 = io_x[26] ? _GEN3306 : _GEN5572;
wire  _GEN5574 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5575 = io_x[30] ? _GEN5574 : _GEN3304;
wire  _GEN5576 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5577 = io_x[26] ? _GEN5576 : _GEN5575;
wire  _GEN5578 = io_x[73] ? _GEN5577 : _GEN5573;
wire  _GEN5579 = io_x[33] ? _GEN5578 : _GEN5570;
wire  _GEN5580 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5581 = io_x[30] ? _GEN5580 : _GEN3303;
wire  _GEN5582 = io_x[26] ? _GEN5581 : _GEN3306;
wire  _GEN5583 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5584 = io_x[73] ? _GEN5583 : _GEN5582;
wire  _GEN5585 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5586 = io_x[30] ? _GEN5585 : _GEN3303;
wire  _GEN5587 = io_x[26] ? _GEN5586 : _GEN3306;
wire  _GEN5588 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5589 = io_x[73] ? _GEN5588 : _GEN5587;
wire  _GEN5590 = io_x[33] ? _GEN5589 : _GEN5584;
wire  _GEN5591 = io_x[28] ? _GEN5590 : _GEN5579;
wire  _GEN5592 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5593 = io_x[30] ? _GEN5592 : _GEN3304;
wire  _GEN5594 = io_x[26] ? _GEN3306 : _GEN5593;
wire  _GEN5595 = io_x[73] ? _GEN3308 : _GEN5594;
wire  _GEN5596 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5597 = io_x[30] ? _GEN5596 : _GEN3303;
wire  _GEN5598 = io_x[26] ? _GEN3306 : _GEN5597;
wire  _GEN5599 = io_x[73] ? _GEN3308 : _GEN5598;
wire  _GEN5600 = io_x[33] ? _GEN5599 : _GEN5595;
wire  _GEN5601 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5602 = io_x[30] ? _GEN5601 : _GEN3304;
wire  _GEN5603 = io_x[26] ? _GEN5602 : _GEN3311;
wire  _GEN5604 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5605 = io_x[30] ? _GEN5604 : _GEN3304;
wire  _GEN5606 = io_x[26] ? _GEN3306 : _GEN5605;
wire  _GEN5607 = io_x[73] ? _GEN5606 : _GEN5603;
wire  _GEN5608 = io_x[33] ? _GEN5607 : _GEN3302;
wire  _GEN5609 = io_x[28] ? _GEN5608 : _GEN5600;
wire  _GEN5610 = io_x[18] ? _GEN5609 : _GEN5591;
wire  _GEN5611 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5612 = io_x[26] ? _GEN5611 : _GEN3306;
wire  _GEN5613 = io_x[73] ? _GEN5612 : _GEN3324;
wire  _GEN5614 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5615 = io_x[26] ? _GEN5614 : _GEN3306;
wire  _GEN5616 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5617 = io_x[30] ? _GEN5616 : _GEN3304;
wire  _GEN5618 = io_x[26] ? _GEN5617 : _GEN3311;
wire  _GEN5619 = io_x[73] ? _GEN5618 : _GEN5615;
wire  _GEN5620 = io_x[33] ? _GEN5619 : _GEN5613;
wire  _GEN5621 = io_x[28] ? _GEN5620 : _GEN3498;
wire  _GEN5622 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5623 = io_x[30] ? _GEN5622 : _GEN3304;
wire  _GEN5624 = io_x[26] ? _GEN5623 : _GEN3306;
wire  _GEN5625 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5626 = io_x[26] ? _GEN5625 : _GEN3306;
wire  _GEN5627 = io_x[73] ? _GEN5626 : _GEN5624;
wire  _GEN5628 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5629 = io_x[30] ? _GEN5628 : _GEN3304;
wire  _GEN5630 = io_x[26] ? _GEN5629 : _GEN3311;
wire  _GEN5631 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5632 = io_x[73] ? _GEN5631 : _GEN5630;
wire  _GEN5633 = io_x[33] ? _GEN5632 : _GEN5627;
wire  _GEN5634 = io_x[28] ? _GEN5633 : _GEN4086;
wire  _GEN5635 = io_x[18] ? _GEN5634 : _GEN5621;
wire  _GEN5636 = io_x[25] ? _GEN5635 : _GEN5610;
wire  _GEN5637 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5638 = io_x[26] ? _GEN5637 : _GEN3306;
wire  _GEN5639 = io_x[73] ? _GEN5638 : _GEN3308;
wire  _GEN5640 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5641 = io_x[30] ? _GEN5640 : _GEN3304;
wire  _GEN5642 = io_x[26] ? _GEN5641 : _GEN3306;
wire  _GEN5643 = io_x[73] ? _GEN3308 : _GEN5642;
wire  _GEN5644 = io_x[33] ? _GEN5643 : _GEN5639;
wire  _GEN5645 = io_x[73] ? _GEN3324 : _GEN3308;
wire  _GEN5646 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5647 = io_x[30] ? _GEN5646 : _GEN3303;
wire  _GEN5648 = io_x[26] ? _GEN3311 : _GEN5647;
wire  _GEN5649 = io_x[73] ? _GEN5648 : _GEN3308;
wire  _GEN5650 = io_x[33] ? _GEN5649 : _GEN5645;
wire  _GEN5651 = io_x[28] ? _GEN5650 : _GEN5644;
wire  _GEN5652 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5653 = io_x[30] ? _GEN3304 : _GEN5652;
wire  _GEN5654 = io_x[26] ? _GEN5653 : _GEN3306;
wire  _GEN5655 = io_x[73] ? _GEN3324 : _GEN5654;
wire  _GEN5656 = io_x[33] ? _GEN5655 : _GEN3371;
wire  _GEN5657 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5658 = io_x[26] ? _GEN5657 : _GEN3306;
wire  _GEN5659 = io_x[73] ? _GEN3308 : _GEN5658;
wire  _GEN5660 = io_x[33] ? _GEN5659 : _GEN3302;
wire  _GEN5661 = io_x[28] ? _GEN5660 : _GEN5656;
wire  _GEN5662 = io_x[18] ? _GEN5661 : _GEN5651;
wire  _GEN5663 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5664 = io_x[26] ? _GEN5663 : _GEN3306;
wire  _GEN5665 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5666 = io_x[26] ? _GEN5665 : _GEN3306;
wire  _GEN5667 = io_x[73] ? _GEN5666 : _GEN5664;
wire  _GEN5668 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5669 = io_x[30] ? _GEN5668 : _GEN3304;
wire  _GEN5670 = io_x[26] ? _GEN5669 : _GEN3306;
wire  _GEN5671 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5672 = io_x[30] ? _GEN5671 : _GEN3304;
wire  _GEN5673 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5674 = io_x[30] ? _GEN3303 : _GEN5673;
wire  _GEN5675 = io_x[26] ? _GEN5674 : _GEN5672;
wire  _GEN5676 = io_x[73] ? _GEN5675 : _GEN5670;
wire  _GEN5677 = io_x[33] ? _GEN5676 : _GEN5667;
wire  _GEN5678 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5679 = io_x[30] ? _GEN5678 : _GEN3303;
wire  _GEN5680 = io_x[26] ? _GEN5679 : _GEN3306;
wire  _GEN5681 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5682 = io_x[30] ? _GEN5681 : _GEN3304;
wire  _GEN5683 = io_x[26] ? _GEN5682 : _GEN3306;
wire  _GEN5684 = io_x[73] ? _GEN5683 : _GEN5680;
wire  _GEN5685 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5686 = io_x[30] ? _GEN5685 : _GEN3303;
wire  _GEN5687 = io_x[26] ? _GEN5686 : _GEN3306;
wire  _GEN5688 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5689 = io_x[30] ? _GEN5688 : _GEN3304;
wire  _GEN5690 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5691 = io_x[30] ? _GEN5690 : _GEN3304;
wire  _GEN5692 = io_x[26] ? _GEN5691 : _GEN5689;
wire  _GEN5693 = io_x[73] ? _GEN5692 : _GEN5687;
wire  _GEN5694 = io_x[33] ? _GEN5693 : _GEN5684;
wire  _GEN5695 = io_x[28] ? _GEN5694 : _GEN5677;
wire  _GEN5696 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5697 = io_x[30] ? _GEN3304 : _GEN5696;
wire  _GEN5698 = io_x[26] ? _GEN5697 : _GEN3306;
wire  _GEN5699 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5700 = io_x[30] ? _GEN5699 : _GEN3303;
wire  _GEN5701 = io_x[26] ? _GEN3306 : _GEN5700;
wire  _GEN5702 = io_x[73] ? _GEN5701 : _GEN5698;
wire  _GEN5703 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5704 = io_x[30] ? _GEN3304 : _GEN5703;
wire  _GEN5705 = io_x[26] ? _GEN5704 : _GEN3311;
wire  _GEN5706 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5707 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5708 = io_x[30] ? _GEN5707 : _GEN5706;
wire  _GEN5709 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5710 = io_x[30] ? _GEN3304 : _GEN5709;
wire  _GEN5711 = io_x[26] ? _GEN5710 : _GEN5708;
wire  _GEN5712 = io_x[73] ? _GEN5711 : _GEN5705;
wire  _GEN5713 = io_x[33] ? _GEN5712 : _GEN5702;
wire  _GEN5714 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5715 = io_x[73] ? _GEN3308 : _GEN5714;
wire  _GEN5716 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5717 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5718 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5719 = io_x[30] ? _GEN5718 : _GEN3304;
wire  _GEN5720 = io_x[26] ? _GEN5719 : _GEN5717;
wire  _GEN5721 = io_x[73] ? _GEN5720 : _GEN5716;
wire  _GEN5722 = io_x[33] ? _GEN5721 : _GEN5715;
wire  _GEN5723 = io_x[28] ? _GEN5722 : _GEN5713;
wire  _GEN5724 = io_x[18] ? _GEN5723 : _GEN5695;
wire  _GEN5725 = io_x[25] ? _GEN5724 : _GEN5662;
wire  _GEN5726 = io_x[29] ? _GEN5725 : _GEN5636;
wire  _GEN5727 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5728 = io_x[30] ? _GEN5727 : _GEN3304;
wire  _GEN5729 = io_x[26] ? _GEN5728 : _GEN3306;
wire  _GEN5730 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5731 = io_x[30] ? _GEN5730 : _GEN3304;
wire  _GEN5732 = io_x[26] ? _GEN5731 : _GEN3306;
wire  _GEN5733 = io_x[73] ? _GEN5732 : _GEN5729;
wire  _GEN5734 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5735 = io_x[30] ? _GEN5734 : _GEN3304;
wire  _GEN5736 = io_x[26] ? _GEN5735 : _GEN3306;
wire  _GEN5737 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5738 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5739 = io_x[30] ? _GEN5738 : _GEN3304;
wire  _GEN5740 = io_x[26] ? _GEN5739 : _GEN5737;
wire  _GEN5741 = io_x[73] ? _GEN5740 : _GEN5736;
wire  _GEN5742 = io_x[33] ? _GEN5741 : _GEN5733;
wire  _GEN5743 = io_x[28] ? _GEN5742 : _GEN4086;
wire  _GEN5744 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5745 = io_x[30] ? _GEN5744 : _GEN3304;
wire  _GEN5746 = io_x[26] ? _GEN5745 : _GEN3311;
wire  _GEN5747 = io_x[73] ? _GEN3308 : _GEN5746;
wire  _GEN5748 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5749 = io_x[30] ? _GEN5748 : _GEN3303;
wire  _GEN5750 = io_x[26] ? _GEN5749 : _GEN3306;
wire  _GEN5751 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5752 = io_x[30] ? _GEN5751 : _GEN3304;
wire  _GEN5753 = io_x[26] ? _GEN5752 : _GEN3306;
wire  _GEN5754 = io_x[73] ? _GEN5753 : _GEN5750;
wire  _GEN5755 = io_x[33] ? _GEN5754 : _GEN5747;
wire  _GEN5756 = io_x[28] ? _GEN5755 : _GEN4086;
wire  _GEN5757 = io_x[18] ? _GEN5756 : _GEN5743;
wire  _GEN5758 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5759 = io_x[30] ? _GEN5758 : _GEN3304;
wire  _GEN5760 = io_x[26] ? _GEN3306 : _GEN5759;
wire  _GEN5761 = io_x[73] ? _GEN5760 : _GEN3308;
wire  _GEN5762 = io_x[33] ? _GEN3302 : _GEN5761;
wire  _GEN5763 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5764 = io_x[73] ? _GEN5763 : _GEN3324;
wire  _GEN5765 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5766 = io_x[30] ? _GEN5765 : _GEN3304;
wire  _GEN5767 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5768 = io_x[30] ? _GEN5767 : _GEN3304;
wire  _GEN5769 = io_x[26] ? _GEN5768 : _GEN5766;
wire  _GEN5770 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5771 = io_x[30] ? _GEN5770 : _GEN3303;
wire  _GEN5772 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5773 = io_x[26] ? _GEN5772 : _GEN5771;
wire  _GEN5774 = io_x[73] ? _GEN5773 : _GEN5769;
wire  _GEN5775 = io_x[33] ? _GEN5774 : _GEN5764;
wire  _GEN5776 = io_x[28] ? _GEN5775 : _GEN5762;
wire  _GEN5777 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5778 = io_x[30] ? _GEN5777 : _GEN3304;
wire  _GEN5779 = io_x[26] ? _GEN5778 : _GEN3311;
wire  _GEN5780 = io_x[73] ? _GEN3308 : _GEN5779;
wire  _GEN5781 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5782 = io_x[30] ? _GEN5781 : _GEN3304;
wire  _GEN5783 = io_x[26] ? _GEN5782 : _GEN3306;
wire  _GEN5784 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5785 = io_x[30] ? _GEN5784 : _GEN3304;
wire  _GEN5786 = io_x[26] ? _GEN3306 : _GEN5785;
wire  _GEN5787 = io_x[73] ? _GEN5786 : _GEN5783;
wire  _GEN5788 = io_x[33] ? _GEN5787 : _GEN5780;
wire  _GEN5789 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5790 = io_x[30] ? _GEN5789 : _GEN3304;
wire  _GEN5791 = io_x[26] ? _GEN3306 : _GEN5790;
wire  _GEN5792 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5793 = io_x[73] ? _GEN5792 : _GEN5791;
wire  _GEN5794 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5795 = io_x[30] ? _GEN5794 : _GEN3304;
wire  _GEN5796 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5797 = io_x[26] ? _GEN5796 : _GEN5795;
wire  _GEN5798 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5799 = io_x[30] ? _GEN5798 : _GEN3304;
wire  _GEN5800 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5801 = io_x[30] ? _GEN5800 : _GEN3304;
wire  _GEN5802 = io_x[26] ? _GEN5801 : _GEN5799;
wire  _GEN5803 = io_x[73] ? _GEN5802 : _GEN5797;
wire  _GEN5804 = io_x[33] ? _GEN5803 : _GEN5793;
wire  _GEN5805 = io_x[28] ? _GEN5804 : _GEN5788;
wire  _GEN5806 = io_x[18] ? _GEN5805 : _GEN5776;
wire  _GEN5807 = io_x[25] ? _GEN5806 : _GEN5757;
wire  _GEN5808 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5809 = io_x[30] ? _GEN3304 : _GEN5808;
wire  _GEN5810 = io_x[26] ? _GEN5809 : _GEN3306;
wire  _GEN5811 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5812 = io_x[30] ? _GEN3304 : _GEN5811;
wire  _GEN5813 = io_x[26] ? _GEN5812 : _GEN3306;
wire  _GEN5814 = io_x[73] ? _GEN5813 : _GEN5810;
wire  _GEN5815 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5816 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5817 = io_x[30] ? _GEN5816 : _GEN5815;
wire  _GEN5818 = io_x[26] ? _GEN5817 : _GEN3306;
wire  _GEN5819 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5820 = io_x[30] ? _GEN3304 : _GEN5819;
wire  _GEN5821 = io_x[26] ? _GEN5820 : _GEN3306;
wire  _GEN5822 = io_x[73] ? _GEN5821 : _GEN5818;
wire  _GEN5823 = io_x[33] ? _GEN5822 : _GEN5814;
wire  _GEN5824 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5825 = io_x[30] ? _GEN5824 : _GEN3304;
wire  _GEN5826 = io_x[26] ? _GEN3311 : _GEN5825;
wire  _GEN5827 = io_x[73] ? _GEN3324 : _GEN5826;
wire  _GEN5828 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5829 = io_x[73] ? _GEN3324 : _GEN5828;
wire  _GEN5830 = io_x[33] ? _GEN5829 : _GEN5827;
wire  _GEN5831 = io_x[28] ? _GEN5830 : _GEN5823;
wire  _GEN5832 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5833 = io_x[30] ? _GEN3304 : _GEN5832;
wire  _GEN5834 = io_x[26] ? _GEN5833 : _GEN3306;
wire  _GEN5835 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5836 = io_x[73] ? _GEN5835 : _GEN5834;
wire  _GEN5837 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5838 = io_x[30] ? _GEN3304 : _GEN5837;
wire  _GEN5839 = io_x[26] ? _GEN5838 : _GEN3311;
wire  _GEN5840 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5841 = io_x[73] ? _GEN5840 : _GEN5839;
wire  _GEN5842 = io_x[33] ? _GEN5841 : _GEN5836;
wire  _GEN5843 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN5844 = io_x[73] ? _GEN5843 : _GEN3308;
wire  _GEN5845 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5846 = io_x[26] ? _GEN3306 : _GEN5845;
wire  _GEN5847 = io_x[73] ? _GEN5846 : _GEN3308;
wire  _GEN5848 = io_x[33] ? _GEN5847 : _GEN5844;
wire  _GEN5849 = io_x[28] ? _GEN5848 : _GEN5842;
wire  _GEN5850 = io_x[18] ? _GEN5849 : _GEN5831;
wire  _GEN5851 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5852 = io_x[30] ? _GEN5851 : _GEN3303;
wire  _GEN5853 = io_x[26] ? _GEN3306 : _GEN5852;
wire  _GEN5854 = io_x[73] ? _GEN5853 : _GEN3308;
wire  _GEN5855 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5856 = io_x[30] ? _GEN5855 : _GEN3304;
wire  _GEN5857 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5858 = io_x[30] ? _GEN3303 : _GEN5857;
wire  _GEN5859 = io_x[26] ? _GEN5858 : _GEN5856;
wire  _GEN5860 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5861 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5862 = io_x[30] ? _GEN5861 : _GEN5860;
wire  _GEN5863 = io_x[26] ? _GEN3306 : _GEN5862;
wire  _GEN5864 = io_x[73] ? _GEN5863 : _GEN5859;
wire  _GEN5865 = io_x[33] ? _GEN5864 : _GEN5854;
wire  _GEN5866 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5867 = io_x[30] ? _GEN5866 : _GEN3304;
wire  _GEN5868 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5869 = io_x[30] ? _GEN5868 : _GEN3304;
wire  _GEN5870 = io_x[26] ? _GEN5869 : _GEN5867;
wire  _GEN5871 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5872 = io_x[30] ? _GEN5871 : _GEN3304;
wire  _GEN5873 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5874 = io_x[30] ? _GEN5873 : _GEN3303;
wire  _GEN5875 = io_x[26] ? _GEN5874 : _GEN5872;
wire  _GEN5876 = io_x[73] ? _GEN5875 : _GEN5870;
wire  _GEN5877 = io_x[33] ? _GEN5876 : _GEN3302;
wire  _GEN5878 = io_x[28] ? _GEN5877 : _GEN5865;
wire  _GEN5879 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5880 = io_x[30] ? _GEN5879 : _GEN3304;
wire  _GEN5881 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5882 = io_x[30] ? _GEN3304 : _GEN5881;
wire  _GEN5883 = io_x[26] ? _GEN5882 : _GEN5880;
wire  _GEN5884 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5885 = io_x[26] ? _GEN3311 : _GEN5884;
wire  _GEN5886 = io_x[73] ? _GEN5885 : _GEN5883;
wire  _GEN5887 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5888 = io_x[30] ? _GEN5887 : _GEN3303;
wire  _GEN5889 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5890 = io_x[26] ? _GEN5889 : _GEN5888;
wire  _GEN5891 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5892 = io_x[30] ? _GEN5891 : _GEN3304;
wire  _GEN5893 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5894 = io_x[26] ? _GEN5893 : _GEN5892;
wire  _GEN5895 = io_x[73] ? _GEN5894 : _GEN5890;
wire  _GEN5896 = io_x[33] ? _GEN5895 : _GEN5886;
wire  _GEN5897 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5898 = io_x[30] ? _GEN3303 : _GEN5897;
wire  _GEN5899 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5900 = io_x[30] ? _GEN5899 : _GEN3304;
wire  _GEN5901 = io_x[26] ? _GEN5900 : _GEN5898;
wire  _GEN5902 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5903 = io_x[30] ? _GEN5902 : _GEN3304;
wire  _GEN5904 = io_x[26] ? _GEN5903 : _GEN3306;
wire  _GEN5905 = io_x[73] ? _GEN5904 : _GEN5901;
wire  _GEN5906 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5907 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5908 = io_x[30] ? _GEN5907 : _GEN5906;
wire  _GEN5909 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5910 = io_x[30] ? _GEN5909 : _GEN3303;
wire  _GEN5911 = io_x[26] ? _GEN5910 : _GEN5908;
wire  _GEN5912 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5913 = io_x[30] ? _GEN5912 : _GEN3304;
wire  _GEN5914 = io_x[26] ? _GEN5913 : _GEN3311;
wire  _GEN5915 = io_x[73] ? _GEN5914 : _GEN5911;
wire  _GEN5916 = io_x[33] ? _GEN5915 : _GEN5905;
wire  _GEN5917 = io_x[28] ? _GEN5916 : _GEN5896;
wire  _GEN5918 = io_x[18] ? _GEN5917 : _GEN5878;
wire  _GEN5919 = io_x[25] ? _GEN5918 : _GEN5850;
wire  _GEN5920 = io_x[29] ? _GEN5919 : _GEN5807;
wire  _GEN5921 = io_x[23] ? _GEN5920 : _GEN5726;
wire  _GEN5922 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5923 = io_x[30] ? _GEN5922 : _GEN3304;
wire  _GEN5924 = io_x[26] ? _GEN3306 : _GEN5923;
wire  _GEN5925 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5926 = io_x[30] ? _GEN5925 : _GEN3304;
wire  _GEN5927 = io_x[26] ? _GEN3306 : _GEN5926;
wire  _GEN5928 = io_x[73] ? _GEN5927 : _GEN5924;
wire  _GEN5929 = io_x[33] ? _GEN5928 : _GEN3302;
wire  _GEN5930 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5931 = io_x[30] ? _GEN3304 : _GEN5930;
wire  _GEN5932 = io_x[26] ? _GEN5931 : _GEN3306;
wire  _GEN5933 = io_x[73] ? _GEN3324 : _GEN5932;
wire  _GEN5934 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5935 = io_x[30] ? _GEN3304 : _GEN5934;
wire  _GEN5936 = io_x[26] ? _GEN5935 : _GEN3306;
wire  _GEN5937 = io_x[73] ? _GEN3324 : _GEN5936;
wire  _GEN5938 = io_x[33] ? _GEN5937 : _GEN5933;
wire  _GEN5939 = io_x[28] ? _GEN5938 : _GEN5929;
wire  _GEN5940 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5941 = io_x[30] ? _GEN5940 : _GEN3304;
wire  _GEN5942 = io_x[26] ? _GEN3306 : _GEN5941;
wire  _GEN5943 = io_x[73] ? _GEN3308 : _GEN5942;
wire  _GEN5944 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5945 = io_x[30] ? _GEN5944 : _GEN3304;
wire  _GEN5946 = io_x[26] ? _GEN3306 : _GEN5945;
wire  _GEN5947 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN5948 = io_x[73] ? _GEN5947 : _GEN5946;
wire  _GEN5949 = io_x[33] ? _GEN5948 : _GEN5943;
wire  _GEN5950 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5951 = io_x[30] ? _GEN3304 : _GEN5950;
wire  _GEN5952 = io_x[26] ? _GEN5951 : _GEN3306;
wire  _GEN5953 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5954 = io_x[26] ? _GEN5953 : _GEN3306;
wire  _GEN5955 = io_x[73] ? _GEN5954 : _GEN5952;
wire  _GEN5956 = io_x[33] ? _GEN5955 : _GEN3302;
wire  _GEN5957 = io_x[28] ? _GEN5956 : _GEN5949;
wire  _GEN5958 = io_x[18] ? _GEN5957 : _GEN5939;
wire  _GEN5959 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5960 = io_x[26] ? _GEN3306 : _GEN5959;
wire  _GEN5961 = io_x[73] ? _GEN5960 : _GEN3308;
wire  _GEN5962 = io_x[33] ? _GEN5961 : _GEN3302;
wire  _GEN5963 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN5964 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5965 = io_x[26] ? _GEN5964 : _GEN5963;
wire  _GEN5966 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5967 = io_x[26] ? _GEN5966 : _GEN3311;
wire  _GEN5968 = io_x[73] ? _GEN5967 : _GEN5965;
wire  _GEN5969 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5970 = io_x[30] ? _GEN5969 : _GEN3304;
wire  _GEN5971 = io_x[26] ? _GEN5970 : _GEN3311;
wire  _GEN5972 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5973 = io_x[30] ? _GEN5972 : _GEN3303;
wire  _GEN5974 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5975 = io_x[26] ? _GEN5974 : _GEN5973;
wire  _GEN5976 = io_x[73] ? _GEN5975 : _GEN5971;
wire  _GEN5977 = io_x[33] ? _GEN5976 : _GEN5968;
wire  _GEN5978 = io_x[28] ? _GEN5977 : _GEN5962;
wire  _GEN5979 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5980 = io_x[30] ? _GEN5979 : _GEN3303;
wire  _GEN5981 = io_x[26] ? _GEN3306 : _GEN5980;
wire  _GEN5982 = io_x[73] ? _GEN5981 : _GEN3324;
wire  _GEN5983 = io_x[33] ? _GEN5982 : _GEN3371;
wire  _GEN5984 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5985 = io_x[30] ? _GEN5984 : _GEN3303;
wire  _GEN5986 = io_x[26] ? _GEN5985 : _GEN3306;
wire  _GEN5987 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5988 = io_x[26] ? _GEN3311 : _GEN5987;
wire  _GEN5989 = io_x[73] ? _GEN5988 : _GEN5986;
wire  _GEN5990 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN5991 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN5992 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN5993 = io_x[30] ? _GEN5992 : _GEN5991;
wire  _GEN5994 = io_x[26] ? _GEN5993 : _GEN5990;
wire  _GEN5995 = io_x[73] ? _GEN3308 : _GEN5994;
wire  _GEN5996 = io_x[33] ? _GEN5995 : _GEN5989;
wire  _GEN5997 = io_x[28] ? _GEN5996 : _GEN5983;
wire  _GEN5998 = io_x[18] ? _GEN5997 : _GEN5978;
wire  _GEN5999 = io_x[25] ? _GEN5998 : _GEN5958;
wire  _GEN6000 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6001 = io_x[30] ? _GEN3303 : _GEN6000;
wire  _GEN6002 = io_x[26] ? _GEN6001 : _GEN3306;
wire  _GEN6003 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN6004 = io_x[26] ? _GEN6003 : _GEN3311;
wire  _GEN6005 = io_x[73] ? _GEN6004 : _GEN6002;
wire  _GEN6006 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6007 = io_x[30] ? _GEN3303 : _GEN6006;
wire  _GEN6008 = io_x[26] ? _GEN6007 : _GEN3306;
wire  _GEN6009 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN6010 = io_x[26] ? _GEN6009 : _GEN3311;
wire  _GEN6011 = io_x[73] ? _GEN6010 : _GEN6008;
wire  _GEN6012 = io_x[33] ? _GEN6011 : _GEN6005;
wire  _GEN6013 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6014 = io_x[30] ? _GEN3304 : _GEN6013;
wire  _GEN6015 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN6016 = io_x[26] ? _GEN6015 : _GEN6014;
wire  _GEN6017 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6018 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6019 = io_x[30] ? _GEN6018 : _GEN6017;
wire  _GEN6020 = io_x[26] ? _GEN3306 : _GEN6019;
wire  _GEN6021 = io_x[73] ? _GEN6020 : _GEN6016;
wire  _GEN6022 = io_x[33] ? _GEN6021 : _GEN3371;
wire  _GEN6023 = io_x[28] ? _GEN6022 : _GEN6012;
wire  _GEN6024 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN6025 = io_x[26] ? _GEN6024 : _GEN3306;
wire  _GEN6026 = io_x[73] ? _GEN3308 : _GEN6025;
wire  _GEN6027 = io_x[33] ? _GEN6026 : _GEN3371;
wire  _GEN6028 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6029 = io_x[30] ? _GEN3303 : _GEN6028;
wire  _GEN6030 = io_x[26] ? _GEN3311 : _GEN6029;
wire  _GEN6031 = io_x[73] ? _GEN3324 : _GEN6030;
wire  _GEN6032 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6033 = io_x[30] ? _GEN3303 : _GEN6032;
wire  _GEN6034 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN6035 = io_x[26] ? _GEN6034 : _GEN6033;
wire  _GEN6036 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6037 = io_x[30] ? _GEN6036 : _GEN3304;
wire  _GEN6038 = io_x[26] ? _GEN3311 : _GEN6037;
wire  _GEN6039 = io_x[73] ? _GEN6038 : _GEN6035;
wire  _GEN6040 = io_x[33] ? _GEN6039 : _GEN6031;
wire  _GEN6041 = io_x[28] ? _GEN6040 : _GEN6027;
wire  _GEN6042 = io_x[18] ? _GEN6041 : _GEN6023;
wire  _GEN6043 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN6044 = io_x[26] ? _GEN3306 : _GEN6043;
wire  _GEN6045 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6046 = io_x[30] ? _GEN3304 : _GEN6045;
wire  _GEN6047 = io_x[26] ? _GEN6046 : _GEN3311;
wire  _GEN6048 = io_x[73] ? _GEN6047 : _GEN6044;
wire  _GEN6049 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6050 = io_x[30] ? _GEN6049 : _GEN3304;
wire  _GEN6051 = io_x[26] ? _GEN6050 : _GEN3306;
wire  _GEN6052 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6053 = io_x[30] ? _GEN3303 : _GEN6052;
wire  _GEN6054 = io_x[26] ? _GEN6053 : _GEN3311;
wire  _GEN6055 = io_x[73] ? _GEN6054 : _GEN6051;
wire  _GEN6056 = io_x[33] ? _GEN6055 : _GEN6048;
wire  _GEN6057 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6058 = io_x[30] ? _GEN3304 : _GEN6057;
wire  _GEN6059 = io_x[26] ? _GEN6058 : _GEN3306;
wire  _GEN6060 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN6061 = io_x[26] ? _GEN6060 : _GEN3306;
wire  _GEN6062 = io_x[73] ? _GEN6061 : _GEN6059;
wire  _GEN6063 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6064 = io_x[30] ? _GEN6063 : _GEN3303;
wire  _GEN6065 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6066 = io_x[30] ? _GEN6065 : _GEN3304;
wire  _GEN6067 = io_x[26] ? _GEN6066 : _GEN6064;
wire  _GEN6068 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN6069 = io_x[26] ? _GEN6068 : _GEN3306;
wire  _GEN6070 = io_x[73] ? _GEN6069 : _GEN6067;
wire  _GEN6071 = io_x[33] ? _GEN6070 : _GEN6062;
wire  _GEN6072 = io_x[28] ? _GEN6071 : _GEN6056;
wire  _GEN6073 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6074 = io_x[30] ? _GEN6073 : _GEN3303;
wire  _GEN6075 = io_x[26] ? _GEN6074 : _GEN3306;
wire  _GEN6076 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6077 = io_x[30] ? _GEN3304 : _GEN6076;
wire  _GEN6078 = io_x[26] ? _GEN3311 : _GEN6077;
wire  _GEN6079 = io_x[73] ? _GEN6078 : _GEN6075;
wire  _GEN6080 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6081 = io_x[30] ? _GEN6080 : _GEN3303;
wire  _GEN6082 = io_x[26] ? _GEN6081 : _GEN3311;
wire  _GEN6083 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6084 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6085 = io_x[30] ? _GEN6084 : _GEN6083;
wire  _GEN6086 = io_x[26] ? _GEN3311 : _GEN6085;
wire  _GEN6087 = io_x[73] ? _GEN6086 : _GEN6082;
wire  _GEN6088 = io_x[33] ? _GEN6087 : _GEN6079;
wire  _GEN6089 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN6090 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6091 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6092 = io_x[30] ? _GEN6091 : _GEN6090;
wire  _GEN6093 = io_x[26] ? _GEN6092 : _GEN6089;
wire  _GEN6094 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6095 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6096 = io_x[30] ? _GEN6095 : _GEN6094;
wire  _GEN6097 = io_x[26] ? _GEN6096 : _GEN3306;
wire  _GEN6098 = io_x[73] ? _GEN6097 : _GEN6093;
wire  _GEN6099 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN6100 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6101 = io_x[30] ? _GEN6100 : _GEN3304;
wire  _GEN6102 = io_x[26] ? _GEN6101 : _GEN6099;
wire  _GEN6103 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6104 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6105 = io_x[30] ? _GEN6104 : _GEN6103;
wire  _GEN6106 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6107 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6108 = io_x[30] ? _GEN6107 : _GEN6106;
wire  _GEN6109 = io_x[26] ? _GEN6108 : _GEN6105;
wire  _GEN6110 = io_x[73] ? _GEN6109 : _GEN6102;
wire  _GEN6111 = io_x[33] ? _GEN6110 : _GEN6098;
wire  _GEN6112 = io_x[28] ? _GEN6111 : _GEN6088;
wire  _GEN6113 = io_x[18] ? _GEN6112 : _GEN6072;
wire  _GEN6114 = io_x[25] ? _GEN6113 : _GEN6042;
wire  _GEN6115 = io_x[29] ? _GEN6114 : _GEN5999;
wire  _GEN6116 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6117 = io_x[30] ? _GEN6116 : _GEN3304;
wire  _GEN6118 = io_x[26] ? _GEN6117 : _GEN3306;
wire  _GEN6119 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN6120 = io_x[73] ? _GEN6119 : _GEN6118;
wire  _GEN6121 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6122 = io_x[30] ? _GEN6121 : _GEN3304;
wire  _GEN6123 = io_x[26] ? _GEN6122 : _GEN3311;
wire  _GEN6124 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6125 = io_x[30] ? _GEN6124 : _GEN3304;
wire  _GEN6126 = io_x[26] ? _GEN6125 : _GEN3311;
wire  _GEN6127 = io_x[73] ? _GEN6126 : _GEN6123;
wire  _GEN6128 = io_x[33] ? _GEN6127 : _GEN6120;
wire  _GEN6129 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6130 = io_x[30] ? _GEN6129 : _GEN3304;
wire  _GEN6131 = io_x[26] ? _GEN6130 : _GEN3311;
wire  _GEN6132 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6133 = io_x[30] ? _GEN6132 : _GEN3304;
wire  _GEN6134 = io_x[26] ? _GEN6133 : _GEN3306;
wire  _GEN6135 = io_x[73] ? _GEN6134 : _GEN6131;
wire  _GEN6136 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6137 = io_x[30] ? _GEN6136 : _GEN3303;
wire  _GEN6138 = io_x[26] ? _GEN6137 : _GEN3311;
wire  _GEN6139 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6140 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6141 = io_x[30] ? _GEN6140 : _GEN6139;
wire  _GEN6142 = io_x[26] ? _GEN6141 : _GEN3306;
wire  _GEN6143 = io_x[73] ? _GEN6142 : _GEN6138;
wire  _GEN6144 = io_x[33] ? _GEN6143 : _GEN6135;
wire  _GEN6145 = io_x[28] ? _GEN6144 : _GEN6128;
wire  _GEN6146 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6147 = io_x[30] ? _GEN6146 : _GEN3303;
wire  _GEN6148 = io_x[26] ? _GEN6147 : _GEN3311;
wire  _GEN6149 = io_x[73] ? _GEN6148 : _GEN3308;
wire  _GEN6150 = io_x[33] ? _GEN6149 : _GEN3371;
wire  _GEN6151 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6152 = io_x[30] ? _GEN6151 : _GEN3304;
wire  _GEN6153 = io_x[26] ? _GEN6152 : _GEN3306;
wire  _GEN6154 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN6155 = io_x[73] ? _GEN6154 : _GEN6153;
wire  _GEN6156 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6157 = io_x[30] ? _GEN3304 : _GEN6156;
wire  _GEN6158 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6159 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6160 = io_x[30] ? _GEN6159 : _GEN6158;
wire  _GEN6161 = io_x[26] ? _GEN6160 : _GEN6157;
wire  _GEN6162 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6163 = io_x[30] ? _GEN6162 : _GEN3303;
wire  _GEN6164 = io_x[26] ? _GEN6163 : _GEN3311;
wire  _GEN6165 = io_x[73] ? _GEN6164 : _GEN6161;
wire  _GEN6166 = io_x[33] ? _GEN6165 : _GEN6155;
wire  _GEN6167 = io_x[28] ? _GEN6166 : _GEN6150;
wire  _GEN6168 = io_x[18] ? _GEN6167 : _GEN6145;
wire  _GEN6169 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6170 = io_x[30] ? _GEN6169 : _GEN3303;
wire  _GEN6171 = io_x[26] ? _GEN3306 : _GEN6170;
wire  _GEN6172 = io_x[73] ? _GEN3308 : _GEN6171;
wire  _GEN6173 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6174 = io_x[30] ? _GEN6173 : _GEN3303;
wire  _GEN6175 = io_x[26] ? _GEN3306 : _GEN6174;
wire  _GEN6176 = io_x[73] ? _GEN3308 : _GEN6175;
wire  _GEN6177 = io_x[33] ? _GEN6176 : _GEN6172;
wire  _GEN6178 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6179 = io_x[30] ? _GEN3304 : _GEN6178;
wire  _GEN6180 = io_x[26] ? _GEN3311 : _GEN6179;
wire  _GEN6181 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6182 = io_x[30] ? _GEN6181 : _GEN3304;
wire  _GEN6183 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6184 = io_x[30] ? _GEN6183 : _GEN3303;
wire  _GEN6185 = io_x[26] ? _GEN6184 : _GEN6182;
wire  _GEN6186 = io_x[73] ? _GEN6185 : _GEN6180;
wire  _GEN6187 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN6188 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6189 = io_x[30] ? _GEN3303 : _GEN6188;
wire  _GEN6190 = io_x[26] ? _GEN6189 : _GEN6187;
wire  _GEN6191 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN6192 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN6193 = io_x[26] ? _GEN6192 : _GEN6191;
wire  _GEN6194 = io_x[73] ? _GEN6193 : _GEN6190;
wire  _GEN6195 = io_x[33] ? _GEN6194 : _GEN6186;
wire  _GEN6196 = io_x[28] ? _GEN6195 : _GEN6177;
wire  _GEN6197 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6198 = io_x[30] ? _GEN6197 : _GEN3304;
wire  _GEN6199 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6200 = io_x[30] ? _GEN6199 : _GEN3304;
wire  _GEN6201 = io_x[26] ? _GEN6200 : _GEN6198;
wire  _GEN6202 = io_x[73] ? _GEN3308 : _GEN6201;
wire  _GEN6203 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6204 = io_x[30] ? _GEN6203 : _GEN3304;
wire  _GEN6205 = io_x[30] ? _GEN3304 : _GEN3303;
wire  _GEN6206 = io_x[26] ? _GEN6205 : _GEN6204;
wire  _GEN6207 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6208 = io_x[30] ? _GEN6207 : _GEN3304;
wire  _GEN6209 = io_x[26] ? _GEN3311 : _GEN6208;
wire  _GEN6210 = io_x[73] ? _GEN6209 : _GEN6206;
wire  _GEN6211 = io_x[33] ? _GEN6210 : _GEN6202;
wire  _GEN6212 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6213 = io_x[30] ? _GEN6212 : _GEN3303;
wire  _GEN6214 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6215 = io_x[30] ? _GEN3304 : _GEN6214;
wire  _GEN6216 = io_x[26] ? _GEN6215 : _GEN6213;
wire  _GEN6217 = io_x[73] ? _GEN3324 : _GEN6216;
wire  _GEN6218 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6219 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6220 = io_x[30] ? _GEN6219 : _GEN6218;
wire  _GEN6221 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6222 = io_x[30] ? _GEN3304 : _GEN6221;
wire  _GEN6223 = io_x[26] ? _GEN6222 : _GEN6220;
wire  _GEN6224 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6225 = io_x[30] ? _GEN3303 : _GEN6224;
wire  _GEN6226 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6227 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6228 = io_x[30] ? _GEN6227 : _GEN6226;
wire  _GEN6229 = io_x[26] ? _GEN6228 : _GEN6225;
wire  _GEN6230 = io_x[73] ? _GEN6229 : _GEN6223;
wire  _GEN6231 = io_x[33] ? _GEN6230 : _GEN6217;
wire  _GEN6232 = io_x[28] ? _GEN6231 : _GEN6211;
wire  _GEN6233 = io_x[18] ? _GEN6232 : _GEN6196;
wire  _GEN6234 = io_x[25] ? _GEN6233 : _GEN6168;
wire  _GEN6235 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6236 = io_x[30] ? _GEN6235 : _GEN3303;
wire  _GEN6237 = io_x[26] ? _GEN6236 : _GEN3306;
wire  _GEN6238 = io_x[73] ? _GEN6237 : _GEN3324;
wire  _GEN6239 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6240 = io_x[30] ? _GEN6239 : _GEN3303;
wire  _GEN6241 = io_x[26] ? _GEN6240 : _GEN3306;
wire  _GEN6242 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6243 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6244 = io_x[30] ? _GEN6243 : _GEN6242;
wire  _GEN6245 = io_x[26] ? _GEN6244 : _GEN3311;
wire  _GEN6246 = io_x[73] ? _GEN6245 : _GEN6241;
wire  _GEN6247 = io_x[33] ? _GEN6246 : _GEN6238;
wire  _GEN6248 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6249 = io_x[30] ? _GEN3304 : _GEN6248;
wire  _GEN6250 = io_x[26] ? _GEN6249 : _GEN3306;
wire  _GEN6251 = io_x[73] ? _GEN6250 : _GEN3308;
wire  _GEN6252 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6253 = io_x[30] ? _GEN3303 : _GEN6252;
wire  _GEN6254 = io_x[26] ? _GEN6253 : _GEN3306;
wire  _GEN6255 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6256 = io_x[30] ? _GEN3304 : _GEN6255;
wire  _GEN6257 = io_x[26] ? _GEN6256 : _GEN3306;
wire  _GEN6258 = io_x[73] ? _GEN6257 : _GEN6254;
wire  _GEN6259 = io_x[33] ? _GEN6258 : _GEN6251;
wire  _GEN6260 = io_x[28] ? _GEN6259 : _GEN6247;
wire  _GEN6261 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6262 = io_x[30] ? _GEN6261 : _GEN3304;
wire  _GEN6263 = io_x[26] ? _GEN6262 : _GEN3306;
wire  _GEN6264 = io_x[26] ? _GEN3306 : _GEN3311;
wire  _GEN6265 = io_x[73] ? _GEN6264 : _GEN6263;
wire  _GEN6266 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6267 = io_x[30] ? _GEN3304 : _GEN6266;
wire  _GEN6268 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6269 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6270 = io_x[30] ? _GEN6269 : _GEN6268;
wire  _GEN6271 = io_x[26] ? _GEN6270 : _GEN6267;
wire  _GEN6272 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6273 = io_x[30] ? _GEN6272 : _GEN3304;
wire  _GEN6274 = io_x[26] ? _GEN6273 : _GEN3306;
wire  _GEN6275 = io_x[73] ? _GEN6274 : _GEN6271;
wire  _GEN6276 = io_x[33] ? _GEN6275 : _GEN6265;
wire  _GEN6277 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6278 = io_x[30] ? _GEN6277 : _GEN3304;
wire  _GEN6279 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6280 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6281 = io_x[30] ? _GEN6280 : _GEN6279;
wire  _GEN6282 = io_x[26] ? _GEN6281 : _GEN6278;
wire  _GEN6283 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6284 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6285 = io_x[30] ? _GEN6284 : _GEN6283;
wire  _GEN6286 = io_x[26] ? _GEN6285 : _GEN3306;
wire  _GEN6287 = io_x[73] ? _GEN6286 : _GEN6282;
wire  _GEN6288 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN6289 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6290 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6291 = io_x[30] ? _GEN6290 : _GEN6289;
wire  _GEN6292 = io_x[26] ? _GEN6291 : _GEN6288;
wire  _GEN6293 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6294 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6295 = io_x[30] ? _GEN6294 : _GEN6293;
wire  _GEN6296 = io_x[26] ? _GEN6295 : _GEN3311;
wire  _GEN6297 = io_x[73] ? _GEN6296 : _GEN6292;
wire  _GEN6298 = io_x[33] ? _GEN6297 : _GEN6287;
wire  _GEN6299 = io_x[28] ? _GEN6298 : _GEN6276;
wire  _GEN6300 = io_x[18] ? _GEN6299 : _GEN6260;
wire  _GEN6301 = io_x[30] ? _GEN3303 : _GEN3304;
wire  _GEN6302 = io_x[26] ? _GEN3311 : _GEN6301;
wire  _GEN6303 = io_x[73] ? _GEN6302 : _GEN3324;
wire  _GEN6304 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6305 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6306 = io_x[30] ? _GEN6305 : _GEN6304;
wire  _GEN6307 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6308 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6309 = io_x[30] ? _GEN6308 : _GEN6307;
wire  _GEN6310 = io_x[26] ? _GEN6309 : _GEN6306;
wire  _GEN6311 = io_x[26] ? _GEN3311 : _GEN3306;
wire  _GEN6312 = io_x[73] ? _GEN6311 : _GEN6310;
wire  _GEN6313 = io_x[33] ? _GEN6312 : _GEN6303;
wire  _GEN6314 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6315 = io_x[30] ? _GEN6314 : _GEN3304;
wire  _GEN6316 = io_x[26] ? _GEN6315 : _GEN3311;
wire  _GEN6317 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6318 = io_x[30] ? _GEN3304 : _GEN6317;
wire  _GEN6319 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6320 = io_x[30] ? _GEN6319 : _GEN3303;
wire  _GEN6321 = io_x[26] ? _GEN6320 : _GEN6318;
wire  _GEN6322 = io_x[73] ? _GEN6321 : _GEN6316;
wire  _GEN6323 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6324 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6325 = io_x[30] ? _GEN6324 : _GEN6323;
wire  _GEN6326 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6327 = io_x[30] ? _GEN6326 : _GEN3304;
wire  _GEN6328 = io_x[26] ? _GEN6327 : _GEN6325;
wire  _GEN6329 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6330 = io_x[30] ? _GEN3303 : _GEN6329;
wire  _GEN6331 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6332 = io_x[30] ? _GEN6331 : _GEN3303;
wire  _GEN6333 = io_x[26] ? _GEN6332 : _GEN6330;
wire  _GEN6334 = io_x[73] ? _GEN6333 : _GEN6328;
wire  _GEN6335 = io_x[33] ? _GEN6334 : _GEN6322;
wire  _GEN6336 = io_x[28] ? _GEN6335 : _GEN6313;
wire  _GEN6337 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6338 = io_x[30] ? _GEN6337 : _GEN3303;
wire  _GEN6339 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6340 = io_x[30] ? _GEN6339 : _GEN3304;
wire  _GEN6341 = io_x[26] ? _GEN6340 : _GEN6338;
wire  _GEN6342 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6343 = io_x[30] ? _GEN3303 : _GEN6342;
wire  _GEN6344 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6345 = io_x[30] ? _GEN3304 : _GEN6344;
wire  _GEN6346 = io_x[26] ? _GEN6345 : _GEN6343;
wire  _GEN6347 = io_x[73] ? _GEN6346 : _GEN6341;
wire  _GEN6348 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6349 = io_x[30] ? _GEN3304 : _GEN6348;
wire  _GEN6350 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6351 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6352 = io_x[30] ? _GEN6351 : _GEN6350;
wire  _GEN6353 = io_x[26] ? _GEN6352 : _GEN6349;
wire  _GEN6354 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6355 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6356 = io_x[30] ? _GEN6355 : _GEN6354;
wire  _GEN6357 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6358 = io_x[30] ? _GEN6357 : _GEN3304;
wire  _GEN6359 = io_x[26] ? _GEN6358 : _GEN6356;
wire  _GEN6360 = io_x[73] ? _GEN6359 : _GEN6353;
wire  _GEN6361 = io_x[33] ? _GEN6360 : _GEN6347;
wire  _GEN6362 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6363 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6364 = io_x[30] ? _GEN6363 : _GEN6362;
wire  _GEN6365 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6366 = io_x[30] ? _GEN6365 : _GEN3303;
wire  _GEN6367 = io_x[26] ? _GEN6366 : _GEN6364;
wire  _GEN6368 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6369 = io_x[30] ? _GEN3303 : _GEN6368;
wire  _GEN6370 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6371 = io_x[30] ? _GEN6370 : _GEN3303;
wire  _GEN6372 = io_x[26] ? _GEN6371 : _GEN6369;
wire  _GEN6373 = io_x[73] ? _GEN6372 : _GEN6367;
wire  _GEN6374 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6375 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6376 = io_x[30] ? _GEN6375 : _GEN6374;
wire  _GEN6377 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6378 = io_x[30] ? _GEN6377 : _GEN3303;
wire  _GEN6379 = io_x[26] ? _GEN6378 : _GEN6376;
wire  _GEN6380 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6381 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6382 = io_x[30] ? _GEN6381 : _GEN6380;
wire  _GEN6383 = io_x[22] ? _GEN3312 : _GEN3313;
wire  _GEN6384 = io_x[22] ? _GEN3313 : _GEN3312;
wire  _GEN6385 = io_x[30] ? _GEN6384 : _GEN6383;
wire  _GEN6386 = io_x[26] ? _GEN6385 : _GEN6382;
wire  _GEN6387 = io_x[73] ? _GEN6386 : _GEN6379;
wire  _GEN6388 = io_x[33] ? _GEN6387 : _GEN6373;
wire  _GEN6389 = io_x[28] ? _GEN6388 : _GEN6361;
wire  _GEN6390 = io_x[18] ? _GEN6389 : _GEN6336;
wire  _GEN6391 = io_x[25] ? _GEN6390 : _GEN6300;
wire  _GEN6392 = io_x[29] ? _GEN6391 : _GEN6234;
wire  _GEN6393 = io_x[23] ? _GEN6392 : _GEN6115;
wire  _GEN6394 = io_x[31] ? _GEN6393 : _GEN5921;
wire  _GEN6395 = io_x[19] ? _GEN6394 : _GEN5568;
wire  _GEN6396 = io_x[76] ? _GEN6395 : _GEN4957;
assign io_y[17] = _GEN6396;
wire  _GEN6397 = 1'b0;
wire  _GEN6398 = 1'b1;
wire  _GEN6399 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6400 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6401 = io_x[25] ? _GEN6400 : _GEN6399;
wire  _GEN6402 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6403 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6404 = io_x[25] ? _GEN6403 : _GEN6402;
wire  _GEN6405 = io_x[73] ? _GEN6404 : _GEN6401;
wire  _GEN6406 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6407 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6408 = io_x[25] ? _GEN6407 : _GEN6406;
wire  _GEN6409 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6410 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6411 = io_x[25] ? _GEN6410 : _GEN6409;
wire  _GEN6412 = io_x[73] ? _GEN6411 : _GEN6408;
wire  _GEN6413 = io_x[75] ? _GEN6412 : _GEN6405;
wire  _GEN6414 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6415 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6416 = io_x[25] ? _GEN6415 : _GEN6414;
wire  _GEN6417 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6418 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6419 = io_x[25] ? _GEN6418 : _GEN6417;
wire  _GEN6420 = io_x[73] ? _GEN6419 : _GEN6416;
wire  _GEN6421 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6422 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6423 = io_x[25] ? _GEN6422 : _GEN6421;
wire  _GEN6424 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6425 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6426 = io_x[25] ? _GEN6425 : _GEN6424;
wire  _GEN6427 = io_x[73] ? _GEN6426 : _GEN6423;
wire  _GEN6428 = io_x[75] ? _GEN6427 : _GEN6420;
wire  _GEN6429 = io_x[21] ? _GEN6428 : _GEN6413;
wire  _GEN6430 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6431 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6432 = io_x[25] ? _GEN6431 : _GEN6430;
wire  _GEN6433 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6434 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6435 = io_x[25] ? _GEN6434 : _GEN6433;
wire  _GEN6436 = io_x[73] ? _GEN6435 : _GEN6432;
wire  _GEN6437 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6438 = 1'b1;
wire  _GEN6439 = io_x[25] ? _GEN6438 : _GEN6437;
wire  _GEN6440 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6441 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6442 = io_x[25] ? _GEN6441 : _GEN6440;
wire  _GEN6443 = io_x[73] ? _GEN6442 : _GEN6439;
wire  _GEN6444 = io_x[75] ? _GEN6443 : _GEN6436;
wire  _GEN6445 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6446 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6447 = io_x[25] ? _GEN6446 : _GEN6445;
wire  _GEN6448 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6449 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6450 = io_x[25] ? _GEN6449 : _GEN6448;
wire  _GEN6451 = io_x[73] ? _GEN6450 : _GEN6447;
wire  _GEN6452 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6453 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6454 = io_x[25] ? _GEN6453 : _GEN6452;
wire  _GEN6455 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6456 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6457 = io_x[25] ? _GEN6456 : _GEN6455;
wire  _GEN6458 = io_x[73] ? _GEN6457 : _GEN6454;
wire  _GEN6459 = io_x[75] ? _GEN6458 : _GEN6451;
wire  _GEN6460 = io_x[21] ? _GEN6459 : _GEN6444;
wire  _GEN6461 = io_x[71] ? _GEN6460 : _GEN6429;
wire  _GEN6462 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6463 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6464 = io_x[25] ? _GEN6463 : _GEN6462;
wire  _GEN6465 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6466 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6467 = io_x[25] ? _GEN6466 : _GEN6465;
wire  _GEN6468 = io_x[73] ? _GEN6467 : _GEN6464;
wire  _GEN6469 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6470 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6471 = io_x[25] ? _GEN6470 : _GEN6469;
wire  _GEN6472 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6473 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6474 = io_x[25] ? _GEN6473 : _GEN6472;
wire  _GEN6475 = io_x[73] ? _GEN6474 : _GEN6471;
wire  _GEN6476 = io_x[75] ? _GEN6475 : _GEN6468;
wire  _GEN6477 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6478 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6479 = io_x[25] ? _GEN6478 : _GEN6477;
wire  _GEN6480 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6481 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6482 = io_x[25] ? _GEN6481 : _GEN6480;
wire  _GEN6483 = io_x[73] ? _GEN6482 : _GEN6479;
wire  _GEN6484 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6485 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6486 = io_x[25] ? _GEN6485 : _GEN6484;
wire  _GEN6487 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6488 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6489 = io_x[25] ? _GEN6488 : _GEN6487;
wire  _GEN6490 = io_x[73] ? _GEN6489 : _GEN6486;
wire  _GEN6491 = io_x[75] ? _GEN6490 : _GEN6483;
wire  _GEN6492 = io_x[21] ? _GEN6491 : _GEN6476;
wire  _GEN6493 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6494 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6495 = io_x[25] ? _GEN6494 : _GEN6493;
wire  _GEN6496 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6497 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6498 = io_x[25] ? _GEN6497 : _GEN6496;
wire  _GEN6499 = io_x[73] ? _GEN6498 : _GEN6495;
wire  _GEN6500 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6501 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6502 = io_x[25] ? _GEN6501 : _GEN6500;
wire  _GEN6503 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6504 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6505 = io_x[25] ? _GEN6504 : _GEN6503;
wire  _GEN6506 = io_x[73] ? _GEN6505 : _GEN6502;
wire  _GEN6507 = io_x[75] ? _GEN6506 : _GEN6499;
wire  _GEN6508 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6509 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6510 = io_x[25] ? _GEN6509 : _GEN6508;
wire  _GEN6511 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6512 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6513 = io_x[25] ? _GEN6512 : _GEN6511;
wire  _GEN6514 = io_x[73] ? _GEN6513 : _GEN6510;
wire  _GEN6515 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6516 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6517 = io_x[25] ? _GEN6516 : _GEN6515;
wire  _GEN6518 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6519 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6520 = io_x[25] ? _GEN6519 : _GEN6518;
wire  _GEN6521 = io_x[73] ? _GEN6520 : _GEN6517;
wire  _GEN6522 = io_x[75] ? _GEN6521 : _GEN6514;
wire  _GEN6523 = io_x[21] ? _GEN6522 : _GEN6507;
wire  _GEN6524 = io_x[71] ? _GEN6523 : _GEN6492;
wire  _GEN6525 = io_x[29] ? _GEN6524 : _GEN6461;
wire  _GEN6526 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6527 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6528 = io_x[25] ? _GEN6527 : _GEN6526;
wire  _GEN6529 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6530 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6531 = io_x[25] ? _GEN6530 : _GEN6529;
wire  _GEN6532 = io_x[73] ? _GEN6531 : _GEN6528;
wire  _GEN6533 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6534 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6535 = io_x[25] ? _GEN6534 : _GEN6533;
wire  _GEN6536 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6537 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6538 = io_x[25] ? _GEN6537 : _GEN6536;
wire  _GEN6539 = io_x[73] ? _GEN6538 : _GEN6535;
wire  _GEN6540 = io_x[75] ? _GEN6539 : _GEN6532;
wire  _GEN6541 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6542 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6543 = io_x[25] ? _GEN6542 : _GEN6541;
wire  _GEN6544 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6545 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6546 = io_x[25] ? _GEN6545 : _GEN6544;
wire  _GEN6547 = io_x[73] ? _GEN6546 : _GEN6543;
wire  _GEN6548 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6549 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6550 = io_x[25] ? _GEN6549 : _GEN6548;
wire  _GEN6551 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6552 = io_x[25] ? _GEN6551 : _GEN6438;
wire  _GEN6553 = io_x[73] ? _GEN6552 : _GEN6550;
wire  _GEN6554 = io_x[75] ? _GEN6553 : _GEN6547;
wire  _GEN6555 = io_x[21] ? _GEN6554 : _GEN6540;
wire  _GEN6556 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6557 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6558 = io_x[25] ? _GEN6557 : _GEN6556;
wire  _GEN6559 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6560 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6561 = io_x[25] ? _GEN6560 : _GEN6559;
wire  _GEN6562 = io_x[73] ? _GEN6561 : _GEN6558;
wire  _GEN6563 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6564 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6565 = io_x[25] ? _GEN6564 : _GEN6563;
wire  _GEN6566 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6567 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6568 = io_x[25] ? _GEN6567 : _GEN6566;
wire  _GEN6569 = io_x[73] ? _GEN6568 : _GEN6565;
wire  _GEN6570 = io_x[75] ? _GEN6569 : _GEN6562;
wire  _GEN6571 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6572 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6573 = io_x[25] ? _GEN6572 : _GEN6571;
wire  _GEN6574 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6575 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6576 = io_x[25] ? _GEN6575 : _GEN6574;
wire  _GEN6577 = io_x[73] ? _GEN6576 : _GEN6573;
wire  _GEN6578 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6579 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6580 = io_x[25] ? _GEN6579 : _GEN6578;
wire  _GEN6581 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6582 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6583 = io_x[25] ? _GEN6582 : _GEN6581;
wire  _GEN6584 = io_x[73] ? _GEN6583 : _GEN6580;
wire  _GEN6585 = io_x[75] ? _GEN6584 : _GEN6577;
wire  _GEN6586 = io_x[21] ? _GEN6585 : _GEN6570;
wire  _GEN6587 = io_x[71] ? _GEN6586 : _GEN6555;
wire  _GEN6588 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6589 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6590 = io_x[25] ? _GEN6589 : _GEN6588;
wire  _GEN6591 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6592 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6593 = io_x[25] ? _GEN6592 : _GEN6591;
wire  _GEN6594 = io_x[73] ? _GEN6593 : _GEN6590;
wire  _GEN6595 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6596 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6597 = io_x[25] ? _GEN6596 : _GEN6595;
wire  _GEN6598 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6599 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6600 = io_x[25] ? _GEN6599 : _GEN6598;
wire  _GEN6601 = io_x[73] ? _GEN6600 : _GEN6597;
wire  _GEN6602 = io_x[75] ? _GEN6601 : _GEN6594;
wire  _GEN6603 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6604 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6605 = io_x[25] ? _GEN6604 : _GEN6603;
wire  _GEN6606 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6607 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6608 = io_x[25] ? _GEN6607 : _GEN6606;
wire  _GEN6609 = io_x[73] ? _GEN6608 : _GEN6605;
wire  _GEN6610 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6611 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6612 = io_x[25] ? _GEN6611 : _GEN6610;
wire  _GEN6613 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6614 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6615 = io_x[25] ? _GEN6614 : _GEN6613;
wire  _GEN6616 = io_x[73] ? _GEN6615 : _GEN6612;
wire  _GEN6617 = io_x[75] ? _GEN6616 : _GEN6609;
wire  _GEN6618 = io_x[21] ? _GEN6617 : _GEN6602;
wire  _GEN6619 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6620 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6621 = io_x[25] ? _GEN6620 : _GEN6619;
wire  _GEN6622 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6623 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6624 = io_x[25] ? _GEN6623 : _GEN6622;
wire  _GEN6625 = io_x[73] ? _GEN6624 : _GEN6621;
wire  _GEN6626 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6627 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6628 = io_x[25] ? _GEN6627 : _GEN6626;
wire  _GEN6629 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6630 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6631 = io_x[25] ? _GEN6630 : _GEN6629;
wire  _GEN6632 = io_x[73] ? _GEN6631 : _GEN6628;
wire  _GEN6633 = io_x[75] ? _GEN6632 : _GEN6625;
wire  _GEN6634 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6635 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6636 = io_x[25] ? _GEN6635 : _GEN6634;
wire  _GEN6637 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6638 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6639 = io_x[25] ? _GEN6638 : _GEN6637;
wire  _GEN6640 = io_x[73] ? _GEN6639 : _GEN6636;
wire  _GEN6641 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6642 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6643 = io_x[25] ? _GEN6642 : _GEN6641;
wire  _GEN6644 = io_x[17] ? _GEN6397 : _GEN6398;
wire  _GEN6645 = io_x[17] ? _GEN6398 : _GEN6397;
wire  _GEN6646 = io_x[25] ? _GEN6645 : _GEN6644;
wire  _GEN6647 = io_x[73] ? _GEN6646 : _GEN6643;
wire  _GEN6648 = io_x[75] ? _GEN6647 : _GEN6640;
wire  _GEN6649 = io_x[21] ? _GEN6648 : _GEN6633;
wire  _GEN6650 = io_x[71] ? _GEN6649 : _GEN6618;
wire  _GEN6651 = io_x[29] ? _GEN6650 : _GEN6587;
wire  _GEN6652 = io_x[79] ? _GEN6651 : _GEN6525;
assign io_y[16] = _GEN6652;
wire  _GEN6653 = 1'b0;
wire  _GEN6654 = 1'b1;
wire  _GEN6655 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6656 = 1'b0;
wire  _GEN6657 = io_x[24] ? _GEN6656 : _GEN6655;
wire  _GEN6658 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6659 = io_x[24] ? _GEN6658 : _GEN6656;
wire  _GEN6660 = io_x[74] ? _GEN6659 : _GEN6657;
wire  _GEN6661 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6662 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6663 = io_x[24] ? _GEN6662 : _GEN6661;
wire  _GEN6664 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6665 = io_x[24] ? _GEN6664 : _GEN6656;
wire  _GEN6666 = io_x[74] ? _GEN6665 : _GEN6663;
wire  _GEN6667 = io_x[19] ? _GEN6666 : _GEN6660;
wire  _GEN6668 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6669 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6670 = io_x[24] ? _GEN6669 : _GEN6668;
wire  _GEN6671 = 1'b1;
wire  _GEN6672 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6673 = io_x[24] ? _GEN6672 : _GEN6671;
wire  _GEN6674 = io_x[74] ? _GEN6673 : _GEN6670;
wire  _GEN6675 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6676 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6677 = io_x[24] ? _GEN6676 : _GEN6675;
wire  _GEN6678 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6679 = io_x[24] ? _GEN6678 : _GEN6671;
wire  _GEN6680 = io_x[74] ? _GEN6679 : _GEN6677;
wire  _GEN6681 = io_x[19] ? _GEN6680 : _GEN6674;
wire  _GEN6682 = io_x[21] ? _GEN6681 : _GEN6667;
wire  _GEN6683 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6684 = io_x[24] ? _GEN6656 : _GEN6683;
wire  _GEN6685 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6686 = io_x[24] ? _GEN6671 : _GEN6685;
wire  _GEN6687 = io_x[74] ? _GEN6686 : _GEN6684;
wire  _GEN6688 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6689 = io_x[24] ? _GEN6688 : _GEN6656;
wire  _GEN6690 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6691 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6692 = io_x[24] ? _GEN6691 : _GEN6690;
wire  _GEN6693 = io_x[74] ? _GEN6692 : _GEN6689;
wire  _GEN6694 = io_x[19] ? _GEN6693 : _GEN6687;
wire  _GEN6695 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6696 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6697 = io_x[24] ? _GEN6696 : _GEN6695;
wire  _GEN6698 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6699 = io_x[24] ? _GEN6656 : _GEN6698;
wire  _GEN6700 = io_x[74] ? _GEN6699 : _GEN6697;
wire  _GEN6701 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6702 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6703 = io_x[24] ? _GEN6702 : _GEN6701;
wire  _GEN6704 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6705 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6706 = io_x[24] ? _GEN6705 : _GEN6704;
wire  _GEN6707 = io_x[74] ? _GEN6706 : _GEN6703;
wire  _GEN6708 = io_x[19] ? _GEN6707 : _GEN6700;
wire  _GEN6709 = io_x[21] ? _GEN6708 : _GEN6694;
wire  _GEN6710 = io_x[23] ? _GEN6709 : _GEN6682;
wire  _GEN6711 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6712 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6713 = io_x[24] ? _GEN6712 : _GEN6711;
wire  _GEN6714 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6715 = io_x[24] ? _GEN6671 : _GEN6714;
wire  _GEN6716 = io_x[74] ? _GEN6715 : _GEN6713;
wire  _GEN6717 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6718 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6719 = io_x[24] ? _GEN6718 : _GEN6717;
wire  _GEN6720 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6721 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6722 = io_x[24] ? _GEN6721 : _GEN6720;
wire  _GEN6723 = io_x[74] ? _GEN6722 : _GEN6719;
wire  _GEN6724 = io_x[19] ? _GEN6723 : _GEN6716;
wire  _GEN6725 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6726 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6727 = io_x[24] ? _GEN6726 : _GEN6725;
wire  _GEN6728 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6729 = io_x[24] ? _GEN6728 : _GEN6671;
wire  _GEN6730 = io_x[74] ? _GEN6729 : _GEN6727;
wire  _GEN6731 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6732 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6733 = io_x[24] ? _GEN6732 : _GEN6731;
wire  _GEN6734 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6735 = io_x[24] ? _GEN6734 : _GEN6671;
wire  _GEN6736 = io_x[74] ? _GEN6735 : _GEN6733;
wire  _GEN6737 = io_x[19] ? _GEN6736 : _GEN6730;
wire  _GEN6738 = io_x[21] ? _GEN6737 : _GEN6724;
wire  _GEN6739 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6740 = io_x[24] ? _GEN6739 : _GEN6656;
wire  _GEN6741 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6742 = io_x[24] ? _GEN6671 : _GEN6741;
wire  _GEN6743 = io_x[74] ? _GEN6742 : _GEN6740;
wire  _GEN6744 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6745 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6746 = io_x[24] ? _GEN6745 : _GEN6744;
wire  _GEN6747 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6748 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6749 = io_x[24] ? _GEN6748 : _GEN6747;
wire  _GEN6750 = io_x[74] ? _GEN6749 : _GEN6746;
wire  _GEN6751 = io_x[19] ? _GEN6750 : _GEN6743;
wire  _GEN6752 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6753 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6754 = io_x[24] ? _GEN6753 : _GEN6752;
wire  _GEN6755 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6756 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6757 = io_x[24] ? _GEN6756 : _GEN6755;
wire  _GEN6758 = io_x[74] ? _GEN6757 : _GEN6754;
wire  _GEN6759 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6760 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6761 = io_x[24] ? _GEN6760 : _GEN6759;
wire  _GEN6762 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6763 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6764 = io_x[24] ? _GEN6763 : _GEN6762;
wire  _GEN6765 = io_x[74] ? _GEN6764 : _GEN6761;
wire  _GEN6766 = io_x[19] ? _GEN6765 : _GEN6758;
wire  _GEN6767 = io_x[21] ? _GEN6766 : _GEN6751;
wire  _GEN6768 = io_x[23] ? _GEN6767 : _GEN6738;
wire  _GEN6769 = io_x[25] ? _GEN6768 : _GEN6710;
wire  _GEN6770 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6771 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6772 = io_x[24] ? _GEN6771 : _GEN6770;
wire  _GEN6773 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6774 = io_x[24] ? _GEN6656 : _GEN6773;
wire  _GEN6775 = io_x[74] ? _GEN6774 : _GEN6772;
wire  _GEN6776 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6777 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6778 = io_x[24] ? _GEN6777 : _GEN6776;
wire  _GEN6779 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6780 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6781 = io_x[24] ? _GEN6780 : _GEN6779;
wire  _GEN6782 = io_x[74] ? _GEN6781 : _GEN6778;
wire  _GEN6783 = io_x[19] ? _GEN6782 : _GEN6775;
wire  _GEN6784 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6785 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6786 = io_x[24] ? _GEN6785 : _GEN6784;
wire  _GEN6787 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6788 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6789 = io_x[24] ? _GEN6788 : _GEN6787;
wire  _GEN6790 = io_x[74] ? _GEN6789 : _GEN6786;
wire  _GEN6791 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6792 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6793 = io_x[24] ? _GEN6792 : _GEN6791;
wire  _GEN6794 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6795 = io_x[24] ? _GEN6794 : _GEN6671;
wire  _GEN6796 = io_x[74] ? _GEN6795 : _GEN6793;
wire  _GEN6797 = io_x[19] ? _GEN6796 : _GEN6790;
wire  _GEN6798 = io_x[21] ? _GEN6797 : _GEN6783;
wire  _GEN6799 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6800 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6801 = io_x[24] ? _GEN6800 : _GEN6799;
wire  _GEN6802 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6803 = io_x[24] ? _GEN6656 : _GEN6802;
wire  _GEN6804 = io_x[74] ? _GEN6803 : _GEN6801;
wire  _GEN6805 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6806 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6807 = io_x[24] ? _GEN6806 : _GEN6805;
wire  _GEN6808 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6809 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6810 = io_x[24] ? _GEN6809 : _GEN6808;
wire  _GEN6811 = io_x[74] ? _GEN6810 : _GEN6807;
wire  _GEN6812 = io_x[19] ? _GEN6811 : _GEN6804;
wire  _GEN6813 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6814 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6815 = io_x[24] ? _GEN6814 : _GEN6813;
wire  _GEN6816 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6817 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6818 = io_x[24] ? _GEN6817 : _GEN6816;
wire  _GEN6819 = io_x[74] ? _GEN6818 : _GEN6815;
wire  _GEN6820 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6821 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6822 = io_x[24] ? _GEN6821 : _GEN6820;
wire  _GEN6823 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6824 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6825 = io_x[24] ? _GEN6824 : _GEN6823;
wire  _GEN6826 = io_x[74] ? _GEN6825 : _GEN6822;
wire  _GEN6827 = io_x[19] ? _GEN6826 : _GEN6819;
wire  _GEN6828 = io_x[21] ? _GEN6827 : _GEN6812;
wire  _GEN6829 = io_x[23] ? _GEN6828 : _GEN6798;
wire  _GEN6830 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6831 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6832 = io_x[24] ? _GEN6831 : _GEN6830;
wire  _GEN6833 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6834 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6835 = io_x[24] ? _GEN6834 : _GEN6833;
wire  _GEN6836 = io_x[74] ? _GEN6835 : _GEN6832;
wire  _GEN6837 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6838 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6839 = io_x[24] ? _GEN6838 : _GEN6837;
wire  _GEN6840 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6841 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6842 = io_x[24] ? _GEN6841 : _GEN6840;
wire  _GEN6843 = io_x[74] ? _GEN6842 : _GEN6839;
wire  _GEN6844 = io_x[19] ? _GEN6843 : _GEN6836;
wire  _GEN6845 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6846 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6847 = io_x[24] ? _GEN6846 : _GEN6845;
wire  _GEN6848 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6849 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6850 = io_x[24] ? _GEN6849 : _GEN6848;
wire  _GEN6851 = io_x[74] ? _GEN6850 : _GEN6847;
wire  _GEN6852 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6853 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6854 = io_x[24] ? _GEN6853 : _GEN6852;
wire  _GEN6855 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6856 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6857 = io_x[24] ? _GEN6856 : _GEN6855;
wire  _GEN6858 = io_x[74] ? _GEN6857 : _GEN6854;
wire  _GEN6859 = io_x[19] ? _GEN6858 : _GEN6851;
wire  _GEN6860 = io_x[21] ? _GEN6859 : _GEN6844;
wire  _GEN6861 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6862 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6863 = io_x[24] ? _GEN6862 : _GEN6861;
wire  _GEN6864 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6865 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6866 = io_x[24] ? _GEN6865 : _GEN6864;
wire  _GEN6867 = io_x[74] ? _GEN6866 : _GEN6863;
wire  _GEN6868 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6869 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6870 = io_x[24] ? _GEN6869 : _GEN6868;
wire  _GEN6871 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6872 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6873 = io_x[24] ? _GEN6872 : _GEN6871;
wire  _GEN6874 = io_x[74] ? _GEN6873 : _GEN6870;
wire  _GEN6875 = io_x[19] ? _GEN6874 : _GEN6867;
wire  _GEN6876 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6877 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6878 = io_x[24] ? _GEN6877 : _GEN6876;
wire  _GEN6879 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6880 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6881 = io_x[24] ? _GEN6880 : _GEN6879;
wire  _GEN6882 = io_x[74] ? _GEN6881 : _GEN6878;
wire  _GEN6883 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6884 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6885 = io_x[24] ? _GEN6884 : _GEN6883;
wire  _GEN6886 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6887 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6888 = io_x[24] ? _GEN6887 : _GEN6886;
wire  _GEN6889 = io_x[74] ? _GEN6888 : _GEN6885;
wire  _GEN6890 = io_x[19] ? _GEN6889 : _GEN6882;
wire  _GEN6891 = io_x[21] ? _GEN6890 : _GEN6875;
wire  _GEN6892 = io_x[23] ? _GEN6891 : _GEN6860;
wire  _GEN6893 = io_x[25] ? _GEN6892 : _GEN6829;
wire  _GEN6894 = io_x[16] ? _GEN6893 : _GEN6769;
wire  _GEN6895 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6896 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6897 = io_x[24] ? _GEN6896 : _GEN6895;
wire  _GEN6898 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6899 = io_x[24] ? _GEN6898 : _GEN6671;
wire  _GEN6900 = io_x[74] ? _GEN6899 : _GEN6897;
wire  _GEN6901 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6902 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6903 = io_x[24] ? _GEN6902 : _GEN6901;
wire  _GEN6904 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6905 = io_x[24] ? _GEN6904 : _GEN6671;
wire  _GEN6906 = io_x[74] ? _GEN6905 : _GEN6903;
wire  _GEN6907 = io_x[19] ? _GEN6906 : _GEN6900;
wire  _GEN6908 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6909 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6910 = io_x[24] ? _GEN6909 : _GEN6908;
wire  _GEN6911 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6912 = io_x[24] ? _GEN6911 : _GEN6671;
wire  _GEN6913 = io_x[74] ? _GEN6912 : _GEN6910;
wire  _GEN6914 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6915 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6916 = io_x[24] ? _GEN6915 : _GEN6914;
wire  _GEN6917 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6918 = io_x[24] ? _GEN6917 : _GEN6671;
wire  _GEN6919 = io_x[74] ? _GEN6918 : _GEN6916;
wire  _GEN6920 = io_x[19] ? _GEN6919 : _GEN6913;
wire  _GEN6921 = io_x[21] ? _GEN6920 : _GEN6907;
wire  _GEN6922 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6923 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6924 = io_x[24] ? _GEN6923 : _GEN6922;
wire  _GEN6925 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6926 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6927 = io_x[24] ? _GEN6926 : _GEN6925;
wire  _GEN6928 = io_x[74] ? _GEN6927 : _GEN6924;
wire  _GEN6929 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6930 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6931 = io_x[24] ? _GEN6930 : _GEN6929;
wire  _GEN6932 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6933 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6934 = io_x[24] ? _GEN6933 : _GEN6932;
wire  _GEN6935 = io_x[74] ? _GEN6934 : _GEN6931;
wire  _GEN6936 = io_x[19] ? _GEN6935 : _GEN6928;
wire  _GEN6937 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6938 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6939 = io_x[24] ? _GEN6938 : _GEN6937;
wire  _GEN6940 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6941 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6942 = io_x[24] ? _GEN6941 : _GEN6940;
wire  _GEN6943 = io_x[74] ? _GEN6942 : _GEN6939;
wire  _GEN6944 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6945 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6946 = io_x[24] ? _GEN6945 : _GEN6944;
wire  _GEN6947 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6948 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6949 = io_x[24] ? _GEN6948 : _GEN6947;
wire  _GEN6950 = io_x[74] ? _GEN6949 : _GEN6946;
wire  _GEN6951 = io_x[19] ? _GEN6950 : _GEN6943;
wire  _GEN6952 = io_x[21] ? _GEN6951 : _GEN6936;
wire  _GEN6953 = io_x[23] ? _GEN6952 : _GEN6921;
wire  _GEN6954 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6955 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6956 = io_x[24] ? _GEN6955 : _GEN6954;
wire  _GEN6957 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6958 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6959 = io_x[24] ? _GEN6958 : _GEN6957;
wire  _GEN6960 = io_x[74] ? _GEN6959 : _GEN6956;
wire  _GEN6961 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6962 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6963 = io_x[24] ? _GEN6962 : _GEN6961;
wire  _GEN6964 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6965 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6966 = io_x[24] ? _GEN6965 : _GEN6964;
wire  _GEN6967 = io_x[74] ? _GEN6966 : _GEN6963;
wire  _GEN6968 = io_x[19] ? _GEN6967 : _GEN6960;
wire  _GEN6969 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6970 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6971 = io_x[24] ? _GEN6970 : _GEN6969;
wire  _GEN6972 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6973 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6974 = io_x[24] ? _GEN6973 : _GEN6972;
wire  _GEN6975 = io_x[74] ? _GEN6974 : _GEN6971;
wire  _GEN6976 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6977 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6978 = io_x[24] ? _GEN6977 : _GEN6976;
wire  _GEN6979 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6980 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6981 = io_x[24] ? _GEN6980 : _GEN6979;
wire  _GEN6982 = io_x[74] ? _GEN6981 : _GEN6978;
wire  _GEN6983 = io_x[19] ? _GEN6982 : _GEN6975;
wire  _GEN6984 = io_x[21] ? _GEN6983 : _GEN6968;
wire  _GEN6985 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6986 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6987 = io_x[24] ? _GEN6986 : _GEN6985;
wire  _GEN6988 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6989 = io_x[24] ? _GEN6988 : _GEN6671;
wire  _GEN6990 = io_x[74] ? _GEN6989 : _GEN6987;
wire  _GEN6991 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6992 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6993 = io_x[24] ? _GEN6992 : _GEN6991;
wire  _GEN6994 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN6995 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN6996 = io_x[24] ? _GEN6995 : _GEN6994;
wire  _GEN6997 = io_x[74] ? _GEN6996 : _GEN6993;
wire  _GEN6998 = io_x[19] ? _GEN6997 : _GEN6990;
wire  _GEN6999 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7000 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7001 = io_x[24] ? _GEN7000 : _GEN6999;
wire  _GEN7002 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7003 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7004 = io_x[24] ? _GEN7003 : _GEN7002;
wire  _GEN7005 = io_x[74] ? _GEN7004 : _GEN7001;
wire  _GEN7006 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7007 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7008 = io_x[24] ? _GEN7007 : _GEN7006;
wire  _GEN7009 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7010 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7011 = io_x[24] ? _GEN7010 : _GEN7009;
wire  _GEN7012 = io_x[74] ? _GEN7011 : _GEN7008;
wire  _GEN7013 = io_x[19] ? _GEN7012 : _GEN7005;
wire  _GEN7014 = io_x[21] ? _GEN7013 : _GEN6998;
wire  _GEN7015 = io_x[23] ? _GEN7014 : _GEN6984;
wire  _GEN7016 = io_x[25] ? _GEN7015 : _GEN6953;
wire  _GEN7017 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7018 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7019 = io_x[24] ? _GEN7018 : _GEN7017;
wire  _GEN7020 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7021 = io_x[24] ? _GEN7020 : _GEN6656;
wire  _GEN7022 = io_x[74] ? _GEN7021 : _GEN7019;
wire  _GEN7023 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7024 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7025 = io_x[24] ? _GEN7024 : _GEN7023;
wire  _GEN7026 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7027 = io_x[24] ? _GEN7026 : _GEN6671;
wire  _GEN7028 = io_x[74] ? _GEN7027 : _GEN7025;
wire  _GEN7029 = io_x[19] ? _GEN7028 : _GEN7022;
wire  _GEN7030 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7031 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7032 = io_x[24] ? _GEN7031 : _GEN7030;
wire  _GEN7033 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7034 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7035 = io_x[24] ? _GEN7034 : _GEN7033;
wire  _GEN7036 = io_x[74] ? _GEN7035 : _GEN7032;
wire  _GEN7037 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7038 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7039 = io_x[24] ? _GEN7038 : _GEN7037;
wire  _GEN7040 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7041 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7042 = io_x[24] ? _GEN7041 : _GEN7040;
wire  _GEN7043 = io_x[74] ? _GEN7042 : _GEN7039;
wire  _GEN7044 = io_x[19] ? _GEN7043 : _GEN7036;
wire  _GEN7045 = io_x[21] ? _GEN7044 : _GEN7029;
wire  _GEN7046 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7047 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7048 = io_x[24] ? _GEN7047 : _GEN7046;
wire  _GEN7049 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7050 = io_x[24] ? _GEN6671 : _GEN7049;
wire  _GEN7051 = io_x[74] ? _GEN7050 : _GEN7048;
wire  _GEN7052 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7053 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7054 = io_x[24] ? _GEN7053 : _GEN7052;
wire  _GEN7055 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7056 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7057 = io_x[24] ? _GEN7056 : _GEN7055;
wire  _GEN7058 = io_x[74] ? _GEN7057 : _GEN7054;
wire  _GEN7059 = io_x[19] ? _GEN7058 : _GEN7051;
wire  _GEN7060 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7061 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7062 = io_x[24] ? _GEN7061 : _GEN7060;
wire  _GEN7063 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7064 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7065 = io_x[24] ? _GEN7064 : _GEN7063;
wire  _GEN7066 = io_x[74] ? _GEN7065 : _GEN7062;
wire  _GEN7067 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7068 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7069 = io_x[24] ? _GEN7068 : _GEN7067;
wire  _GEN7070 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7071 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7072 = io_x[24] ? _GEN7071 : _GEN7070;
wire  _GEN7073 = io_x[74] ? _GEN7072 : _GEN7069;
wire  _GEN7074 = io_x[19] ? _GEN7073 : _GEN7066;
wire  _GEN7075 = io_x[21] ? _GEN7074 : _GEN7059;
wire  _GEN7076 = io_x[23] ? _GEN7075 : _GEN7045;
wire  _GEN7077 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7078 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7079 = io_x[24] ? _GEN7078 : _GEN7077;
wire  _GEN7080 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7081 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7082 = io_x[24] ? _GEN7081 : _GEN7080;
wire  _GEN7083 = io_x[74] ? _GEN7082 : _GEN7079;
wire  _GEN7084 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7085 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7086 = io_x[24] ? _GEN7085 : _GEN7084;
wire  _GEN7087 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7088 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7089 = io_x[24] ? _GEN7088 : _GEN7087;
wire  _GEN7090 = io_x[74] ? _GEN7089 : _GEN7086;
wire  _GEN7091 = io_x[19] ? _GEN7090 : _GEN7083;
wire  _GEN7092 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7093 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7094 = io_x[24] ? _GEN7093 : _GEN7092;
wire  _GEN7095 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7096 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7097 = io_x[24] ? _GEN7096 : _GEN7095;
wire  _GEN7098 = io_x[74] ? _GEN7097 : _GEN7094;
wire  _GEN7099 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7100 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7101 = io_x[24] ? _GEN7100 : _GEN7099;
wire  _GEN7102 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7103 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7104 = io_x[24] ? _GEN7103 : _GEN7102;
wire  _GEN7105 = io_x[74] ? _GEN7104 : _GEN7101;
wire  _GEN7106 = io_x[19] ? _GEN7105 : _GEN7098;
wire  _GEN7107 = io_x[21] ? _GEN7106 : _GEN7091;
wire  _GEN7108 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7109 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7110 = io_x[24] ? _GEN7109 : _GEN7108;
wire  _GEN7111 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7112 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7113 = io_x[24] ? _GEN7112 : _GEN7111;
wire  _GEN7114 = io_x[74] ? _GEN7113 : _GEN7110;
wire  _GEN7115 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7116 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7117 = io_x[24] ? _GEN7116 : _GEN7115;
wire  _GEN7118 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7119 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7120 = io_x[24] ? _GEN7119 : _GEN7118;
wire  _GEN7121 = io_x[74] ? _GEN7120 : _GEN7117;
wire  _GEN7122 = io_x[19] ? _GEN7121 : _GEN7114;
wire  _GEN7123 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7124 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7125 = io_x[24] ? _GEN7124 : _GEN7123;
wire  _GEN7126 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7127 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7128 = io_x[24] ? _GEN7127 : _GEN7126;
wire  _GEN7129 = io_x[74] ? _GEN7128 : _GEN7125;
wire  _GEN7130 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7131 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7132 = io_x[24] ? _GEN7131 : _GEN7130;
wire  _GEN7133 = io_x[20] ? _GEN6653 : _GEN6654;
wire  _GEN7134 = io_x[20] ? _GEN6654 : _GEN6653;
wire  _GEN7135 = io_x[24] ? _GEN7134 : _GEN7133;
wire  _GEN7136 = io_x[74] ? _GEN7135 : _GEN7132;
wire  _GEN7137 = io_x[19] ? _GEN7136 : _GEN7129;
wire  _GEN7138 = io_x[21] ? _GEN7137 : _GEN7122;
wire  _GEN7139 = io_x[23] ? _GEN7138 : _GEN7107;
wire  _GEN7140 = io_x[25] ? _GEN7139 : _GEN7076;
wire  _GEN7141 = io_x[16] ? _GEN7140 : _GEN7016;
wire  _GEN7142 = io_x[28] ? _GEN7141 : _GEN6894;
assign io_y[15] = _GEN7142;
wire  _GEN7143 = 1'b0;
wire  _GEN7144 = 1'b1;
wire  _GEN7145 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7146 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7147 = io_x[71] ? _GEN7146 : _GEN7145;
wire  _GEN7148 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7149 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7150 = io_x[71] ? _GEN7149 : _GEN7148;
wire  _GEN7151 = io_x[77] ? _GEN7150 : _GEN7147;
wire  _GEN7152 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7153 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7154 = io_x[71] ? _GEN7153 : _GEN7152;
wire  _GEN7155 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7156 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7157 = io_x[71] ? _GEN7156 : _GEN7155;
wire  _GEN7158 = io_x[77] ? _GEN7157 : _GEN7154;
wire  _GEN7159 = io_x[33] ? _GEN7158 : _GEN7151;
wire  _GEN7160 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7161 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7162 = io_x[71] ? _GEN7161 : _GEN7160;
wire  _GEN7163 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7164 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7165 = io_x[71] ? _GEN7164 : _GEN7163;
wire  _GEN7166 = io_x[77] ? _GEN7165 : _GEN7162;
wire  _GEN7167 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7168 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7169 = io_x[71] ? _GEN7168 : _GEN7167;
wire  _GEN7170 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7171 = io_x[73] ? _GEN7144 : _GEN7143;
wire  _GEN7172 = io_x[71] ? _GEN7171 : _GEN7170;
wire  _GEN7173 = io_x[77] ? _GEN7172 : _GEN7169;
wire  _GEN7174 = io_x[33] ? _GEN7173 : _GEN7166;
wire  _GEN7175 = io_x[72] ? _GEN7174 : _GEN7159;
assign io_y[14] = _GEN7175;
wire  _GEN7176 = 1'b0;
wire  _GEN7177 = 1'b1;
wire  _GEN7178 = io_x[72] ? _GEN7177 : _GEN7176;
wire  _GEN7179 = io_x[72] ? _GEN7177 : _GEN7176;
wire  _GEN7180 = io_x[32] ? _GEN7179 : _GEN7178;
assign io_y[13] = _GEN7180;
wire  _GEN7181 = 1'b0;
wire  _GEN7182 = 1'b1;
wire  _GEN7183 = io_x[71] ? _GEN7182 : _GEN7181;
assign io_y[12] = _GEN7183;
wire  _GEN7184 = 1'b0;
wire  _GEN7185 = 1'b1;
wire  _GEN7186 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7187 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7188 = io_x[71] ? _GEN7187 : _GEN7186;
wire  _GEN7189 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7190 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7191 = io_x[71] ? _GEN7190 : _GEN7189;
wire  _GEN7192 = io_x[21] ? _GEN7191 : _GEN7188;
wire  _GEN7193 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7194 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7195 = io_x[71] ? _GEN7194 : _GEN7193;
wire  _GEN7196 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7197 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7198 = io_x[71] ? _GEN7197 : _GEN7196;
wire  _GEN7199 = io_x[21] ? _GEN7198 : _GEN7195;
wire  _GEN7200 = io_x[19] ? _GEN7199 : _GEN7192;
wire  _GEN7201 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7202 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7203 = io_x[71] ? _GEN7202 : _GEN7201;
wire  _GEN7204 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7205 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7206 = io_x[71] ? _GEN7205 : _GEN7204;
wire  _GEN7207 = io_x[21] ? _GEN7206 : _GEN7203;
wire  _GEN7208 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7209 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7210 = io_x[71] ? _GEN7209 : _GEN7208;
wire  _GEN7211 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7212 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7213 = io_x[71] ? _GEN7212 : _GEN7211;
wire  _GEN7214 = io_x[21] ? _GEN7213 : _GEN7210;
wire  _GEN7215 = io_x[19] ? _GEN7214 : _GEN7207;
wire  _GEN7216 = io_x[79] ? _GEN7215 : _GEN7200;
wire  _GEN7217 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7218 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7219 = io_x[71] ? _GEN7218 : _GEN7217;
wire  _GEN7220 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7221 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7222 = io_x[71] ? _GEN7221 : _GEN7220;
wire  _GEN7223 = io_x[21] ? _GEN7222 : _GEN7219;
wire  _GEN7224 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7225 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7226 = io_x[71] ? _GEN7225 : _GEN7224;
wire  _GEN7227 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7228 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7229 = io_x[71] ? _GEN7228 : _GEN7227;
wire  _GEN7230 = io_x[21] ? _GEN7229 : _GEN7226;
wire  _GEN7231 = io_x[19] ? _GEN7230 : _GEN7223;
wire  _GEN7232 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7233 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7234 = io_x[71] ? _GEN7233 : _GEN7232;
wire  _GEN7235 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7236 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7237 = io_x[71] ? _GEN7236 : _GEN7235;
wire  _GEN7238 = io_x[21] ? _GEN7237 : _GEN7234;
wire  _GEN7239 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7240 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7241 = io_x[71] ? _GEN7240 : _GEN7239;
wire  _GEN7242 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7243 = io_x[70] ? _GEN7185 : _GEN7184;
wire  _GEN7244 = io_x[71] ? _GEN7243 : _GEN7242;
wire  _GEN7245 = io_x[21] ? _GEN7244 : _GEN7241;
wire  _GEN7246 = io_x[19] ? _GEN7245 : _GEN7238;
wire  _GEN7247 = io_x[79] ? _GEN7246 : _GEN7231;
wire  _GEN7248 = io_x[33] ? _GEN7247 : _GEN7216;
assign io_y[11] = _GEN7248;
wire  _GEN7249 = 1'b0;
wire  _GEN7250 = 1'b1;
wire  _GEN7251 = io_x[69] ? _GEN7250 : _GEN7249;
wire  _GEN7252 = io_x[69] ? _GEN7250 : _GEN7249;
wire  _GEN7253 = io_x[17] ? _GEN7252 : _GEN7251;
wire  _GEN7254 = io_x[69] ? _GEN7250 : _GEN7249;
wire  _GEN7255 = io_x[69] ? _GEN7250 : _GEN7249;
wire  _GEN7256 = io_x[17] ? _GEN7255 : _GEN7254;
wire  _GEN7257 = io_x[71] ? _GEN7256 : _GEN7253;
wire  _GEN7258 = io_x[69] ? _GEN7250 : _GEN7249;
wire  _GEN7259 = io_x[69] ? _GEN7250 : _GEN7249;
wire  _GEN7260 = io_x[17] ? _GEN7259 : _GEN7258;
wire  _GEN7261 = io_x[69] ? _GEN7250 : _GEN7249;
wire  _GEN7262 = io_x[69] ? _GEN7250 : _GEN7249;
wire  _GEN7263 = io_x[17] ? _GEN7262 : _GEN7261;
wire  _GEN7264 = io_x[71] ? _GEN7263 : _GEN7260;
wire  _GEN7265 = io_x[79] ? _GEN7264 : _GEN7257;
assign io_y[10] = _GEN7265;
wire  _GEN7266 = 1'b0;
wire  _GEN7267 = 1'b1;
wire  _GEN7268 = 1'b1;
wire  _GEN7269 = 1'b0;
wire  _GEN7270 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7271 = 1'b0;
wire  _GEN7272 = io_x[27] ? _GEN7271 : _GEN7270;
wire  _GEN7273 = 1'b0;
wire  _GEN7274 = io_x[19] ? _GEN7273 : _GEN7272;
wire  _GEN7275 = io_x[23] ? _GEN7274 : _GEN7267;
wire  _GEN7276 = io_x[18] ? _GEN7275 : _GEN7266;
wire  _GEN7277 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7278 = 1'b1;
wire  _GEN7279 = io_x[27] ? _GEN7278 : _GEN7277;
wire  _GEN7280 = 1'b1;
wire  _GEN7281 = io_x[19] ? _GEN7280 : _GEN7279;
wire  _GEN7282 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7283 = io_x[27] ? _GEN7282 : _GEN7271;
wire  _GEN7284 = io_x[19] ? _GEN7283 : _GEN7280;
wire  _GEN7285 = io_x[23] ? _GEN7284 : _GEN7281;
wire  _GEN7286 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7287 = io_x[27] ? _GEN7286 : _GEN7278;
wire  _GEN7288 = io_x[19] ? _GEN7287 : _GEN7280;
wire  _GEN7289 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7290 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7291 = io_x[27] ? _GEN7290 : _GEN7289;
wire  _GEN7292 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7293 = io_x[19] ? _GEN7292 : _GEN7291;
wire  _GEN7294 = io_x[23] ? _GEN7293 : _GEN7288;
wire  _GEN7295 = io_x[18] ? _GEN7294 : _GEN7285;
wire  _GEN7296 = io_x[33] ? _GEN7295 : _GEN7276;
wire  _GEN7297 = 1'b1;
wire  _GEN7298 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7299 = io_x[27] ? _GEN7298 : _GEN7278;
wire  _GEN7300 = io_x[19] ? _GEN7280 : _GEN7299;
wire  _GEN7301 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7302 = io_x[19] ? _GEN7280 : _GEN7301;
wire  _GEN7303 = io_x[23] ? _GEN7302 : _GEN7300;
wire  _GEN7304 = io_x[18] ? _GEN7303 : _GEN7297;
wire  _GEN7305 = 1'b0;
wire  _GEN7306 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7307 = io_x[27] ? _GEN7306 : _GEN7278;
wire  _GEN7308 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7309 = io_x[27] ? _GEN7308 : _GEN7278;
wire  _GEN7310 = io_x[19] ? _GEN7309 : _GEN7307;
wire  _GEN7311 = io_x[23] ? _GEN7310 : _GEN7305;
wire  _GEN7312 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7313 = io_x[27] ? _GEN7312 : _GEN7271;
wire  _GEN7314 = io_x[19] ? _GEN7280 : _GEN7313;
wire  _GEN7315 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7316 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7317 = io_x[27] ? _GEN7316 : _GEN7315;
wire  _GEN7318 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7319 = io_x[27] ? _GEN7318 : _GEN7271;
wire  _GEN7320 = io_x[19] ? _GEN7319 : _GEN7317;
wire  _GEN7321 = io_x[23] ? _GEN7320 : _GEN7314;
wire  _GEN7322 = io_x[18] ? _GEN7321 : _GEN7311;
wire  _GEN7323 = io_x[33] ? _GEN7322 : _GEN7304;
wire  _GEN7324 = io_x[31] ? _GEN7323 : _GEN7296;
wire  _GEN7325 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7326 = io_x[27] ? _GEN7325 : _GEN7278;
wire  _GEN7327 = io_x[19] ? _GEN7273 : _GEN7326;
wire  _GEN7328 = io_x[23] ? _GEN7327 : _GEN7305;
wire  _GEN7329 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7330 = io_x[19] ? _GEN7273 : _GEN7329;
wire  _GEN7331 = io_x[23] ? _GEN7330 : _GEN7267;
wire  _GEN7332 = io_x[18] ? _GEN7331 : _GEN7328;
wire  _GEN7333 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN7334 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7335 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7336 = io_x[27] ? _GEN7335 : _GEN7278;
wire  _GEN7337 = io_x[19] ? _GEN7336 : _GEN7334;
wire  _GEN7338 = io_x[23] ? _GEN7337 : _GEN7305;
wire  _GEN7339 = io_x[18] ? _GEN7338 : _GEN7333;
wire  _GEN7340 = io_x[33] ? _GEN7339 : _GEN7332;
wire  _GEN7341 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7342 = io_x[27] ? _GEN7278 : _GEN7341;
wire  _GEN7343 = io_x[19] ? _GEN7342 : _GEN7280;
wire  _GEN7344 = io_x[23] ? _GEN7343 : _GEN7267;
wire  _GEN7345 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN7346 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7347 = io_x[19] ? _GEN7346 : _GEN7280;
wire  _GEN7348 = io_x[23] ? _GEN7347 : _GEN7345;
wire  _GEN7349 = io_x[18] ? _GEN7348 : _GEN7344;
wire  _GEN7350 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7351 = io_x[19] ? _GEN7350 : _GEN7280;
wire  _GEN7352 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7353 = io_x[27] ? _GEN7278 : _GEN7352;
wire  _GEN7354 = io_x[19] ? _GEN7353 : _GEN7280;
wire  _GEN7355 = io_x[23] ? _GEN7354 : _GEN7351;
wire  _GEN7356 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7357 = io_x[19] ? _GEN7280 : _GEN7356;
wire  _GEN7358 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7359 = io_x[27] ? _GEN7358 : _GEN7278;
wire  _GEN7360 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7361 = io_x[27] ? _GEN7360 : _GEN7271;
wire  _GEN7362 = io_x[19] ? _GEN7361 : _GEN7359;
wire  _GEN7363 = io_x[23] ? _GEN7362 : _GEN7357;
wire  _GEN7364 = io_x[18] ? _GEN7363 : _GEN7355;
wire  _GEN7365 = io_x[33] ? _GEN7364 : _GEN7349;
wire  _GEN7366 = io_x[31] ? _GEN7365 : _GEN7340;
wire  _GEN7367 = io_x[28] ? _GEN7366 : _GEN7324;
wire  _GEN7368 = io_x[23] ? _GEN7267 : _GEN7305;
wire  _GEN7369 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7370 = io_x[19] ? _GEN7369 : _GEN7273;
wire  _GEN7371 = io_x[23] ? _GEN7370 : _GEN7267;
wire  _GEN7372 = io_x[18] ? _GEN7371 : _GEN7368;
wire  _GEN7373 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN7374 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7375 = io_x[19] ? _GEN7374 : _GEN7280;
wire  _GEN7376 = io_x[23] ? _GEN7375 : _GEN7373;
wire  _GEN7377 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7378 = io_x[27] ? _GEN7377 : _GEN7278;
wire  _GEN7379 = io_x[19] ? _GEN7378 : _GEN7280;
wire  _GEN7380 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7381 = io_x[27] ? _GEN7380 : _GEN7278;
wire  _GEN7382 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7383 = io_x[19] ? _GEN7382 : _GEN7381;
wire  _GEN7384 = io_x[23] ? _GEN7383 : _GEN7379;
wire  _GEN7385 = io_x[18] ? _GEN7384 : _GEN7376;
wire  _GEN7386 = io_x[33] ? _GEN7385 : _GEN7372;
wire  _GEN7387 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7388 = io_x[19] ? _GEN7280 : _GEN7387;
wire  _GEN7389 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7390 = io_x[27] ? _GEN7389 : _GEN7271;
wire  _GEN7391 = io_x[19] ? _GEN7390 : _GEN7273;
wire  _GEN7392 = io_x[23] ? _GEN7391 : _GEN7388;
wire  _GEN7393 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7394 = io_x[27] ? _GEN7278 : _GEN7393;
wire  _GEN7395 = io_x[19] ? _GEN7394 : _GEN7280;
wire  _GEN7396 = io_x[23] ? _GEN7395 : _GEN7305;
wire  _GEN7397 = io_x[18] ? _GEN7396 : _GEN7392;
wire  _GEN7398 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7399 = io_x[27] ? _GEN7278 : _GEN7398;
wire  _GEN7400 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7401 = io_x[27] ? _GEN7400 : _GEN7278;
wire  _GEN7402 = io_x[19] ? _GEN7401 : _GEN7399;
wire  _GEN7403 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7404 = io_x[19] ? _GEN7403 : _GEN7280;
wire  _GEN7405 = io_x[23] ? _GEN7404 : _GEN7402;
wire  _GEN7406 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7407 = io_x[27] ? _GEN7406 : _GEN7278;
wire  _GEN7408 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7409 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7410 = io_x[27] ? _GEN7409 : _GEN7408;
wire  _GEN7411 = io_x[19] ? _GEN7410 : _GEN7407;
wire  _GEN7412 = io_x[23] ? _GEN7411 : _GEN7267;
wire  _GEN7413 = io_x[18] ? _GEN7412 : _GEN7405;
wire  _GEN7414 = io_x[33] ? _GEN7413 : _GEN7397;
wire  _GEN7415 = io_x[31] ? _GEN7414 : _GEN7386;
wire  _GEN7416 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7417 = io_x[27] ? _GEN7278 : _GEN7416;
wire  _GEN7418 = io_x[19] ? _GEN7417 : _GEN7280;
wire  _GEN7419 = io_x[23] ? _GEN7418 : _GEN7267;
wire  _GEN7420 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN7421 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7422 = io_x[27] ? _GEN7421 : _GEN7271;
wire  _GEN7423 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7424 = io_x[27] ? _GEN7423 : _GEN7278;
wire  _GEN7425 = io_x[19] ? _GEN7424 : _GEN7422;
wire  _GEN7426 = io_x[23] ? _GEN7425 : _GEN7420;
wire  _GEN7427 = io_x[18] ? _GEN7426 : _GEN7419;
wire  _GEN7428 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN7429 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7430 = io_x[27] ? _GEN7271 : _GEN7429;
wire  _GEN7431 = io_x[19] ? _GEN7430 : _GEN7280;
wire  _GEN7432 = io_x[23] ? _GEN7431 : _GEN7428;
wire  _GEN7433 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7434 = io_x[27] ? _GEN7271 : _GEN7433;
wire  _GEN7435 = io_x[19] ? _GEN7434 : _GEN7273;
wire  _GEN7436 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7437 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7438 = io_x[19] ? _GEN7437 : _GEN7436;
wire  _GEN7439 = io_x[23] ? _GEN7438 : _GEN7435;
wire  _GEN7440 = io_x[18] ? _GEN7439 : _GEN7432;
wire  _GEN7441 = io_x[33] ? _GEN7440 : _GEN7427;
wire  _GEN7442 = io_x[23] ? _GEN7267 : _GEN7305;
wire  _GEN7443 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7444 = io_x[27] ? _GEN7443 : _GEN7271;
wire  _GEN7445 = io_x[19] ? _GEN7444 : _GEN7280;
wire  _GEN7446 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7447 = io_x[27] ? _GEN7446 : _GEN7278;
wire  _GEN7448 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7449 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7450 = io_x[27] ? _GEN7449 : _GEN7448;
wire  _GEN7451 = io_x[19] ? _GEN7450 : _GEN7447;
wire  _GEN7452 = io_x[23] ? _GEN7451 : _GEN7445;
wire  _GEN7453 = io_x[18] ? _GEN7452 : _GEN7442;
wire  _GEN7454 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7455 = io_x[19] ? _GEN7454 : _GEN7280;
wire  _GEN7456 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7457 = io_x[27] ? _GEN7456 : _GEN7278;
wire  _GEN7458 = io_x[19] ? _GEN7457 : _GEN7280;
wire  _GEN7459 = io_x[23] ? _GEN7458 : _GEN7455;
wire  _GEN7460 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7461 = io_x[27] ? _GEN7460 : _GEN7278;
wire  _GEN7462 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7463 = io_x[27] ? _GEN7271 : _GEN7462;
wire  _GEN7464 = io_x[19] ? _GEN7463 : _GEN7461;
wire  _GEN7465 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7466 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7467 = io_x[27] ? _GEN7466 : _GEN7465;
wire  _GEN7468 = io_x[19] ? _GEN7467 : _GEN7273;
wire  _GEN7469 = io_x[23] ? _GEN7468 : _GEN7464;
wire  _GEN7470 = io_x[18] ? _GEN7469 : _GEN7459;
wire  _GEN7471 = io_x[33] ? _GEN7470 : _GEN7453;
wire  _GEN7472 = io_x[31] ? _GEN7471 : _GEN7441;
wire  _GEN7473 = io_x[28] ? _GEN7472 : _GEN7415;
wire  _GEN7474 = io_x[26] ? _GEN7473 : _GEN7367;
wire  _GEN7475 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7476 = io_x[27] ? _GEN7475 : _GEN7278;
wire  _GEN7477 = io_x[19] ? _GEN7280 : _GEN7476;
wire  _GEN7478 = io_x[23] ? _GEN7477 : _GEN7267;
wire  _GEN7479 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7480 = io_x[27] ? _GEN7479 : _GEN7278;
wire  _GEN7481 = io_x[19] ? _GEN7273 : _GEN7480;
wire  _GEN7482 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7483 = io_x[27] ? _GEN7482 : _GEN7278;
wire  _GEN7484 = io_x[19] ? _GEN7273 : _GEN7483;
wire  _GEN7485 = io_x[23] ? _GEN7484 : _GEN7481;
wire  _GEN7486 = io_x[18] ? _GEN7485 : _GEN7478;
wire  _GEN7487 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7488 = io_x[27] ? _GEN7487 : _GEN7278;
wire  _GEN7489 = io_x[19] ? _GEN7280 : _GEN7488;
wire  _GEN7490 = io_x[23] ? _GEN7489 : _GEN7267;
wire  _GEN7491 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7492 = io_x[19] ? _GEN7273 : _GEN7491;
wire  _GEN7493 = io_x[23] ? _GEN7492 : _GEN7305;
wire  _GEN7494 = io_x[18] ? _GEN7493 : _GEN7490;
wire  _GEN7495 = io_x[33] ? _GEN7494 : _GEN7486;
wire  _GEN7496 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7497 = io_x[19] ? _GEN7280 : _GEN7496;
wire  _GEN7498 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7499 = io_x[27] ? _GEN7498 : _GEN7278;
wire  _GEN7500 = io_x[19] ? _GEN7280 : _GEN7499;
wire  _GEN7501 = io_x[23] ? _GEN7500 : _GEN7497;
wire  _GEN7502 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7503 = io_x[27] ? _GEN7502 : _GEN7271;
wire  _GEN7504 = io_x[19] ? _GEN7280 : _GEN7503;
wire  _GEN7505 = io_x[23] ? _GEN7504 : _GEN7305;
wire  _GEN7506 = io_x[18] ? _GEN7505 : _GEN7501;
wire  _GEN7507 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7508 = io_x[27] ? _GEN7507 : _GEN7271;
wire  _GEN7509 = io_x[19] ? _GEN7280 : _GEN7508;
wire  _GEN7510 = io_x[23] ? _GEN7509 : _GEN7267;
wire  _GEN7511 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7512 = io_x[27] ? _GEN7511 : _GEN7271;
wire  _GEN7513 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7514 = io_x[27] ? _GEN7271 : _GEN7513;
wire  _GEN7515 = io_x[19] ? _GEN7514 : _GEN7512;
wire  _GEN7516 = io_x[23] ? _GEN7267 : _GEN7515;
wire  _GEN7517 = io_x[18] ? _GEN7516 : _GEN7510;
wire  _GEN7518 = io_x[33] ? _GEN7517 : _GEN7506;
wire  _GEN7519 = io_x[31] ? _GEN7518 : _GEN7495;
wire  _GEN7520 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7521 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7522 = io_x[27] ? _GEN7521 : _GEN7278;
wire  _GEN7523 = io_x[19] ? _GEN7522 : _GEN7520;
wire  _GEN7524 = io_x[23] ? _GEN7523 : _GEN7267;
wire  _GEN7525 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7526 = io_x[27] ? _GEN7525 : _GEN7271;
wire  _GEN7527 = io_x[19] ? _GEN7280 : _GEN7526;
wire  _GEN7528 = io_x[23] ? _GEN7267 : _GEN7527;
wire  _GEN7529 = io_x[18] ? _GEN7528 : _GEN7524;
wire  _GEN7530 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7531 = io_x[27] ? _GEN7530 : _GEN7278;
wire  _GEN7532 = io_x[19] ? _GEN7531 : _GEN7280;
wire  _GEN7533 = io_x[23] ? _GEN7532 : _GEN7305;
wire  _GEN7534 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7535 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7536 = io_x[27] ? _GEN7535 : _GEN7534;
wire  _GEN7537 = io_x[19] ? _GEN7280 : _GEN7536;
wire  _GEN7538 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7539 = io_x[27] ? _GEN7538 : _GEN7278;
wire  _GEN7540 = io_x[19] ? _GEN7539 : _GEN7280;
wire  _GEN7541 = io_x[23] ? _GEN7540 : _GEN7537;
wire  _GEN7542 = io_x[18] ? _GEN7541 : _GEN7533;
wire  _GEN7543 = io_x[33] ? _GEN7542 : _GEN7529;
wire  _GEN7544 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7545 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7546 = io_x[19] ? _GEN7545 : _GEN7544;
wire  _GEN7547 = io_x[23] ? _GEN7546 : _GEN7267;
wire  _GEN7548 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7549 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7550 = io_x[27] ? _GEN7549 : _GEN7548;
wire  _GEN7551 = io_x[19] ? _GEN7550 : _GEN7273;
wire  _GEN7552 = io_x[23] ? _GEN7551 : _GEN7267;
wire  _GEN7553 = io_x[18] ? _GEN7552 : _GEN7547;
wire  _GEN7554 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN7555 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7556 = io_x[27] ? _GEN7555 : _GEN7271;
wire  _GEN7557 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7558 = io_x[27] ? _GEN7557 : _GEN7271;
wire  _GEN7559 = io_x[19] ? _GEN7558 : _GEN7556;
wire  _GEN7560 = io_x[23] ? _GEN7559 : _GEN7554;
wire  _GEN7561 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7562 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7563 = io_x[27] ? _GEN7562 : _GEN7561;
wire  _GEN7564 = io_x[19] ? _GEN7563 : _GEN7273;
wire  _GEN7565 = io_x[23] ? _GEN7564 : _GEN7305;
wire  _GEN7566 = io_x[18] ? _GEN7565 : _GEN7560;
wire  _GEN7567 = io_x[33] ? _GEN7566 : _GEN7553;
wire  _GEN7568 = io_x[31] ? _GEN7567 : _GEN7543;
wire  _GEN7569 = io_x[28] ? _GEN7568 : _GEN7519;
wire  _GEN7570 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7571 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7572 = io_x[27] ? _GEN7571 : _GEN7278;
wire  _GEN7573 = io_x[19] ? _GEN7572 : _GEN7570;
wire  _GEN7574 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7575 = io_x[19] ? _GEN7280 : _GEN7574;
wire  _GEN7576 = io_x[23] ? _GEN7575 : _GEN7573;
wire  _GEN7577 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7578 = io_x[19] ? _GEN7280 : _GEN7577;
wire  _GEN7579 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7580 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7581 = io_x[27] ? _GEN7580 : _GEN7579;
wire  _GEN7582 = io_x[19] ? _GEN7280 : _GEN7581;
wire  _GEN7583 = io_x[23] ? _GEN7582 : _GEN7578;
wire  _GEN7584 = io_x[18] ? _GEN7583 : _GEN7576;
wire  _GEN7585 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7586 = io_x[27] ? _GEN7278 : _GEN7585;
wire  _GEN7587 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7588 = io_x[19] ? _GEN7587 : _GEN7586;
wire  _GEN7589 = io_x[23] ? _GEN7588 : _GEN7305;
wire  _GEN7590 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN7591 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7592 = io_x[27] ? _GEN7591 : _GEN7278;
wire  _GEN7593 = io_x[19] ? _GEN7592 : _GEN7273;
wire  _GEN7594 = io_x[23] ? _GEN7593 : _GEN7590;
wire  _GEN7595 = io_x[18] ? _GEN7594 : _GEN7589;
wire  _GEN7596 = io_x[33] ? _GEN7595 : _GEN7584;
wire  _GEN7597 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN7598 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7599 = io_x[27] ? _GEN7278 : _GEN7598;
wire  _GEN7600 = io_x[19] ? _GEN7599 : _GEN7280;
wire  _GEN7601 = io_x[23] ? _GEN7600 : _GEN7597;
wire  _GEN7602 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7603 = io_x[27] ? _GEN7271 : _GEN7602;
wire  _GEN7604 = io_x[19] ? _GEN7603 : _GEN7280;
wire  _GEN7605 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7606 = io_x[27] ? _GEN7271 : _GEN7605;
wire  _GEN7607 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7608 = io_x[19] ? _GEN7607 : _GEN7606;
wire  _GEN7609 = io_x[23] ? _GEN7608 : _GEN7604;
wire  _GEN7610 = io_x[18] ? _GEN7609 : _GEN7601;
wire  _GEN7611 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7612 = io_x[27] ? _GEN7611 : _GEN7271;
wire  _GEN7613 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7614 = io_x[27] ? _GEN7613 : _GEN7271;
wire  _GEN7615 = io_x[19] ? _GEN7614 : _GEN7612;
wire  _GEN7616 = io_x[23] ? _GEN7615 : _GEN7267;
wire  _GEN7617 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7618 = io_x[27] ? _GEN7278 : _GEN7617;
wire  _GEN7619 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7620 = io_x[27] ? _GEN7278 : _GEN7619;
wire  _GEN7621 = io_x[19] ? _GEN7620 : _GEN7618;
wire  _GEN7622 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7623 = io_x[27] ? _GEN7622 : _GEN7271;
wire  _GEN7624 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7625 = io_x[27] ? _GEN7624 : _GEN7278;
wire  _GEN7626 = io_x[19] ? _GEN7625 : _GEN7623;
wire  _GEN7627 = io_x[23] ? _GEN7626 : _GEN7621;
wire  _GEN7628 = io_x[18] ? _GEN7627 : _GEN7616;
wire  _GEN7629 = io_x[33] ? _GEN7628 : _GEN7610;
wire  _GEN7630 = io_x[31] ? _GEN7629 : _GEN7596;
wire  _GEN7631 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN7632 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7633 = io_x[19] ? _GEN7280 : _GEN7632;
wire  _GEN7634 = io_x[23] ? _GEN7633 : _GEN7631;
wire  _GEN7635 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7636 = io_x[27] ? _GEN7635 : _GEN7271;
wire  _GEN7637 = io_x[19] ? _GEN7636 : _GEN7273;
wire  _GEN7638 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN7639 = io_x[23] ? _GEN7638 : _GEN7637;
wire  _GEN7640 = io_x[18] ? _GEN7639 : _GEN7634;
wire  _GEN7641 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7642 = io_x[27] ? _GEN7641 : _GEN7271;
wire  _GEN7643 = io_x[19] ? _GEN7280 : _GEN7642;
wire  _GEN7644 = io_x[23] ? _GEN7643 : _GEN7305;
wire  _GEN7645 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7646 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7647 = io_x[27] ? _GEN7278 : _GEN7646;
wire  _GEN7648 = io_x[19] ? _GEN7647 : _GEN7645;
wire  _GEN7649 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN7650 = io_x[23] ? _GEN7649 : _GEN7648;
wire  _GEN7651 = io_x[18] ? _GEN7650 : _GEN7644;
wire  _GEN7652 = io_x[33] ? _GEN7651 : _GEN7640;
wire  _GEN7653 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7654 = io_x[27] ? _GEN7278 : _GEN7653;
wire  _GEN7655 = io_x[19] ? _GEN7654 : _GEN7273;
wire  _GEN7656 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7657 = io_x[27] ? _GEN7656 : _GEN7278;
wire  _GEN7658 = io_x[19] ? _GEN7273 : _GEN7657;
wire  _GEN7659 = io_x[23] ? _GEN7658 : _GEN7655;
wire  _GEN7660 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7661 = io_x[19] ? _GEN7273 : _GEN7660;
wire  _GEN7662 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7663 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7664 = io_x[27] ? _GEN7663 : _GEN7662;
wire  _GEN7665 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7666 = io_x[19] ? _GEN7665 : _GEN7664;
wire  _GEN7667 = io_x[23] ? _GEN7666 : _GEN7661;
wire  _GEN7668 = io_x[18] ? _GEN7667 : _GEN7659;
wire  _GEN7669 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7670 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7671 = io_x[27] ? _GEN7670 : _GEN7278;
wire  _GEN7672 = io_x[19] ? _GEN7671 : _GEN7669;
wire  _GEN7673 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7674 = io_x[27] ? _GEN7673 : _GEN7278;
wire  _GEN7675 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7676 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7677 = io_x[27] ? _GEN7676 : _GEN7675;
wire  _GEN7678 = io_x[19] ? _GEN7677 : _GEN7674;
wire  _GEN7679 = io_x[23] ? _GEN7678 : _GEN7672;
wire  _GEN7680 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7681 = io_x[27] ? _GEN7278 : _GEN7680;
wire  _GEN7682 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7683 = io_x[27] ? _GEN7682 : _GEN7278;
wire  _GEN7684 = io_x[19] ? _GEN7683 : _GEN7681;
wire  _GEN7685 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7686 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7687 = io_x[27] ? _GEN7686 : _GEN7685;
wire  _GEN7688 = io_x[19] ? _GEN7687 : _GEN7280;
wire  _GEN7689 = io_x[23] ? _GEN7688 : _GEN7684;
wire  _GEN7690 = io_x[18] ? _GEN7689 : _GEN7679;
wire  _GEN7691 = io_x[33] ? _GEN7690 : _GEN7668;
wire  _GEN7692 = io_x[31] ? _GEN7691 : _GEN7652;
wire  _GEN7693 = io_x[28] ? _GEN7692 : _GEN7630;
wire  _GEN7694 = io_x[26] ? _GEN7693 : _GEN7569;
wire  _GEN7695 = io_x[20] ? _GEN7694 : _GEN7474;
wire  _GEN7696 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7697 = io_x[19] ? _GEN7696 : _GEN7280;
wire  _GEN7698 = io_x[23] ? _GEN7697 : _GEN7267;
wire  _GEN7699 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7700 = io_x[19] ? _GEN7699 : _GEN7280;
wire  _GEN7701 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7702 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7703 = io_x[19] ? _GEN7702 : _GEN7701;
wire  _GEN7704 = io_x[23] ? _GEN7703 : _GEN7700;
wire  _GEN7705 = io_x[18] ? _GEN7704 : _GEN7698;
wire  _GEN7706 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7707 = io_x[27] ? _GEN7706 : _GEN7278;
wire  _GEN7708 = io_x[19] ? _GEN7280 : _GEN7707;
wire  _GEN7709 = io_x[23] ? _GEN7305 : _GEN7708;
wire  _GEN7710 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7711 = io_x[27] ? _GEN7710 : _GEN7271;
wire  _GEN7712 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7713 = io_x[19] ? _GEN7712 : _GEN7711;
wire  _GEN7714 = io_x[23] ? _GEN7713 : _GEN7305;
wire  _GEN7715 = io_x[18] ? _GEN7714 : _GEN7709;
wire  _GEN7716 = io_x[33] ? _GEN7715 : _GEN7705;
wire  _GEN7717 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN7718 = io_x[23] ? _GEN7267 : _GEN7717;
wire  _GEN7719 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN7720 = io_x[23] ? _GEN7719 : _GEN7267;
wire  _GEN7721 = io_x[18] ? _GEN7720 : _GEN7718;
wire  _GEN7722 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7723 = io_x[27] ? _GEN7722 : _GEN7278;
wire  _GEN7724 = io_x[19] ? _GEN7723 : _GEN7280;
wire  _GEN7725 = io_x[23] ? _GEN7724 : _GEN7267;
wire  _GEN7726 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7727 = io_x[27] ? _GEN7726 : _GEN7278;
wire  _GEN7728 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7729 = io_x[27] ? _GEN7728 : _GEN7278;
wire  _GEN7730 = io_x[19] ? _GEN7729 : _GEN7727;
wire  _GEN7731 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7732 = io_x[27] ? _GEN7731 : _GEN7278;
wire  _GEN7733 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7734 = io_x[19] ? _GEN7733 : _GEN7732;
wire  _GEN7735 = io_x[23] ? _GEN7734 : _GEN7730;
wire  _GEN7736 = io_x[18] ? _GEN7735 : _GEN7725;
wire  _GEN7737 = io_x[33] ? _GEN7736 : _GEN7721;
wire  _GEN7738 = io_x[31] ? _GEN7737 : _GEN7716;
wire  _GEN7739 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7740 = io_x[27] ? _GEN7739 : _GEN7278;
wire  _GEN7741 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7742 = io_x[27] ? _GEN7741 : _GEN7271;
wire  _GEN7743 = io_x[19] ? _GEN7742 : _GEN7740;
wire  _GEN7744 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7745 = io_x[27] ? _GEN7744 : _GEN7278;
wire  _GEN7746 = io_x[19] ? _GEN7273 : _GEN7745;
wire  _GEN7747 = io_x[23] ? _GEN7746 : _GEN7743;
wire  _GEN7748 = io_x[18] ? _GEN7747 : _GEN7266;
wire  _GEN7749 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN7750 = io_x[23] ? _GEN7267 : _GEN7749;
wire  _GEN7751 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7752 = io_x[27] ? _GEN7751 : _GEN7271;
wire  _GEN7753 = io_x[19] ? _GEN7752 : _GEN7280;
wire  _GEN7754 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7755 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7756 = io_x[27] ? _GEN7755 : _GEN7278;
wire  _GEN7757 = io_x[19] ? _GEN7756 : _GEN7754;
wire  _GEN7758 = io_x[23] ? _GEN7757 : _GEN7753;
wire  _GEN7759 = io_x[18] ? _GEN7758 : _GEN7750;
wire  _GEN7760 = io_x[33] ? _GEN7759 : _GEN7748;
wire  _GEN7761 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7762 = io_x[27] ? _GEN7278 : _GEN7761;
wire  _GEN7763 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7764 = io_x[19] ? _GEN7763 : _GEN7762;
wire  _GEN7765 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN7766 = io_x[23] ? _GEN7765 : _GEN7764;
wire  _GEN7767 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7768 = io_x[27] ? _GEN7271 : _GEN7767;
wire  _GEN7769 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7770 = io_x[27] ? _GEN7278 : _GEN7769;
wire  _GEN7771 = io_x[19] ? _GEN7770 : _GEN7768;
wire  _GEN7772 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7773 = io_x[27] ? _GEN7772 : _GEN7278;
wire  _GEN7774 = io_x[19] ? _GEN7273 : _GEN7773;
wire  _GEN7775 = io_x[23] ? _GEN7774 : _GEN7771;
wire  _GEN7776 = io_x[18] ? _GEN7775 : _GEN7766;
wire  _GEN7777 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7778 = io_x[27] ? _GEN7278 : _GEN7777;
wire  _GEN7779 = io_x[19] ? _GEN7778 : _GEN7280;
wire  _GEN7780 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7781 = io_x[27] ? _GEN7278 : _GEN7780;
wire  _GEN7782 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7783 = io_x[19] ? _GEN7782 : _GEN7781;
wire  _GEN7784 = io_x[23] ? _GEN7783 : _GEN7779;
wire  _GEN7785 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7786 = io_x[27] ? _GEN7278 : _GEN7785;
wire  _GEN7787 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7788 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7789 = io_x[27] ? _GEN7788 : _GEN7787;
wire  _GEN7790 = io_x[19] ? _GEN7789 : _GEN7786;
wire  _GEN7791 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7792 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7793 = io_x[27] ? _GEN7792 : _GEN7791;
wire  _GEN7794 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7795 = io_x[27] ? _GEN7794 : _GEN7278;
wire  _GEN7796 = io_x[19] ? _GEN7795 : _GEN7793;
wire  _GEN7797 = io_x[23] ? _GEN7796 : _GEN7790;
wire  _GEN7798 = io_x[18] ? _GEN7797 : _GEN7784;
wire  _GEN7799 = io_x[33] ? _GEN7798 : _GEN7776;
wire  _GEN7800 = io_x[31] ? _GEN7799 : _GEN7760;
wire  _GEN7801 = io_x[28] ? _GEN7800 : _GEN7738;
wire  _GEN7802 = io_x[23] ? _GEN7267 : _GEN7305;
wire  _GEN7803 = io_x[18] ? _GEN7297 : _GEN7802;
wire  _GEN7804 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7805 = io_x[19] ? _GEN7273 : _GEN7804;
wire  _GEN7806 = io_x[23] ? _GEN7267 : _GEN7805;
wire  _GEN7807 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7808 = io_x[27] ? _GEN7271 : _GEN7807;
wire  _GEN7809 = io_x[19] ? _GEN7273 : _GEN7808;
wire  _GEN7810 = io_x[23] ? _GEN7267 : _GEN7809;
wire  _GEN7811 = io_x[18] ? _GEN7810 : _GEN7806;
wire  _GEN7812 = io_x[33] ? _GEN7811 : _GEN7803;
wire  _GEN7813 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7814 = io_x[27] ? _GEN7271 : _GEN7813;
wire  _GEN7815 = io_x[19] ? _GEN7814 : _GEN7280;
wire  _GEN7816 = io_x[23] ? _GEN7305 : _GEN7815;
wire  _GEN7817 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7818 = io_x[27] ? _GEN7817 : _GEN7278;
wire  _GEN7819 = io_x[19] ? _GEN7280 : _GEN7818;
wire  _GEN7820 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7821 = io_x[27] ? _GEN7820 : _GEN7271;
wire  _GEN7822 = io_x[19] ? _GEN7821 : _GEN7280;
wire  _GEN7823 = io_x[23] ? _GEN7822 : _GEN7819;
wire  _GEN7824 = io_x[18] ? _GEN7823 : _GEN7816;
wire  _GEN7825 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7826 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7827 = io_x[27] ? _GEN7826 : _GEN7825;
wire  _GEN7828 = io_x[19] ? _GEN7827 : _GEN7273;
wire  _GEN7829 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7830 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7831 = io_x[27] ? _GEN7830 : _GEN7829;
wire  _GEN7832 = io_x[19] ? _GEN7831 : _GEN7273;
wire  _GEN7833 = io_x[23] ? _GEN7832 : _GEN7828;
wire  _GEN7834 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7835 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7836 = io_x[27] ? _GEN7835 : _GEN7834;
wire  _GEN7837 = io_x[19] ? _GEN7836 : _GEN7280;
wire  _GEN7838 = io_x[23] ? _GEN7837 : _GEN7305;
wire  _GEN7839 = io_x[18] ? _GEN7838 : _GEN7833;
wire  _GEN7840 = io_x[33] ? _GEN7839 : _GEN7824;
wire  _GEN7841 = io_x[31] ? _GEN7840 : _GEN7812;
wire  _GEN7842 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7843 = io_x[27] ? _GEN7278 : _GEN7842;
wire  _GEN7844 = io_x[19] ? _GEN7843 : _GEN7280;
wire  _GEN7845 = io_x[23] ? _GEN7305 : _GEN7844;
wire  _GEN7846 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7847 = io_x[27] ? _GEN7846 : _GEN7278;
wire  _GEN7848 = io_x[19] ? _GEN7273 : _GEN7847;
wire  _GEN7849 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7850 = io_x[27] ? _GEN7849 : _GEN7278;
wire  _GEN7851 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7852 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7853 = io_x[27] ? _GEN7852 : _GEN7851;
wire  _GEN7854 = io_x[19] ? _GEN7853 : _GEN7850;
wire  _GEN7855 = io_x[23] ? _GEN7854 : _GEN7848;
wire  _GEN7856 = io_x[18] ? _GEN7855 : _GEN7845;
wire  _GEN7857 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7858 = io_x[27] ? _GEN7278 : _GEN7857;
wire  _GEN7859 = io_x[19] ? _GEN7858 : _GEN7280;
wire  _GEN7860 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7861 = io_x[27] ? _GEN7860 : _GEN7278;
wire  _GEN7862 = io_x[19] ? _GEN7861 : _GEN7280;
wire  _GEN7863 = io_x[23] ? _GEN7862 : _GEN7859;
wire  _GEN7864 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7865 = io_x[19] ? _GEN7273 : _GEN7864;
wire  _GEN7866 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7867 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7868 = io_x[27] ? _GEN7867 : _GEN7866;
wire  _GEN7869 = io_x[19] ? _GEN7868 : _GEN7273;
wire  _GEN7870 = io_x[23] ? _GEN7869 : _GEN7865;
wire  _GEN7871 = io_x[18] ? _GEN7870 : _GEN7863;
wire  _GEN7872 = io_x[33] ? _GEN7871 : _GEN7856;
wire  _GEN7873 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7874 = io_x[27] ? _GEN7873 : _GEN7278;
wire  _GEN7875 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7876 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7877 = io_x[27] ? _GEN7876 : _GEN7875;
wire  _GEN7878 = io_x[19] ? _GEN7877 : _GEN7874;
wire  _GEN7879 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7880 = io_x[27] ? _GEN7879 : _GEN7278;
wire  _GEN7881 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7882 = io_x[19] ? _GEN7881 : _GEN7880;
wire  _GEN7883 = io_x[23] ? _GEN7882 : _GEN7878;
wire  _GEN7884 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7885 = io_x[19] ? _GEN7280 : _GEN7884;
wire  _GEN7886 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7887 = io_x[27] ? _GEN7886 : _GEN7271;
wire  _GEN7888 = io_x[19] ? _GEN7887 : _GEN7280;
wire  _GEN7889 = io_x[23] ? _GEN7888 : _GEN7885;
wire  _GEN7890 = io_x[18] ? _GEN7889 : _GEN7883;
wire  _GEN7891 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7892 = io_x[27] ? _GEN7891 : _GEN7875;
wire  _GEN7893 = io_x[19] ? _GEN7892 : _GEN7273;
wire  _GEN7894 = io_x[27] ? _GEN7879 : _GEN7278;
wire  _GEN7895 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7896 = io_x[27] ? _GEN7895 : _GEN7271;
wire  _GEN7897 = io_x[19] ? _GEN7896 : _GEN7894;
wire  _GEN7898 = io_x[23] ? _GEN7897 : _GEN7893;
wire  _GEN7899 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7900 = io_x[27] ? _GEN7271 : _GEN7899;
wire  _GEN7901 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7902 = io_x[27] ? _GEN7901 : _GEN7278;
wire  _GEN7903 = io_x[19] ? _GEN7902 : _GEN7900;
wire  _GEN7904 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7905 = io_x[27] ? _GEN7904 : _GEN7278;
wire  _GEN7906 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7907 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7908 = io_x[27] ? _GEN7907 : _GEN7906;
wire  _GEN7909 = io_x[19] ? _GEN7908 : _GEN7905;
wire  _GEN7910 = io_x[23] ? _GEN7909 : _GEN7903;
wire  _GEN7911 = io_x[18] ? _GEN7910 : _GEN7898;
wire  _GEN7912 = io_x[33] ? _GEN7911 : _GEN7890;
wire  _GEN7913 = io_x[31] ? _GEN7912 : _GEN7872;
wire  _GEN7914 = io_x[28] ? _GEN7913 : _GEN7841;
wire  _GEN7915 = io_x[26] ? _GEN7914 : _GEN7801;
wire  _GEN7916 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7917 = io_x[27] ? _GEN7916 : _GEN7278;
wire  _GEN7918 = io_x[19] ? _GEN7917 : _GEN7280;
wire  _GEN7919 = io_x[23] ? _GEN7918 : _GEN7305;
wire  _GEN7920 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7921 = io_x[27] ? _GEN7920 : _GEN7278;
wire  _GEN7922 = io_x[19] ? _GEN7280 : _GEN7921;
wire  _GEN7923 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7924 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7925 = io_x[27] ? _GEN7924 : _GEN7278;
wire  _GEN7926 = io_x[19] ? _GEN7925 : _GEN7923;
wire  _GEN7927 = io_x[23] ? _GEN7926 : _GEN7922;
wire  _GEN7928 = io_x[18] ? _GEN7927 : _GEN7919;
wire  _GEN7929 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7930 = io_x[27] ? _GEN7929 : _GEN7271;
wire  _GEN7931 = io_x[19] ? _GEN7280 : _GEN7930;
wire  _GEN7932 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7933 = io_x[27] ? _GEN7932 : _GEN7278;
wire  _GEN7934 = io_x[19] ? _GEN7933 : _GEN7280;
wire  _GEN7935 = io_x[23] ? _GEN7934 : _GEN7931;
wire  _GEN7936 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN7937 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7938 = io_x[27] ? _GEN7937 : _GEN7278;
wire  _GEN7939 = io_x[19] ? _GEN7938 : _GEN7273;
wire  _GEN7940 = io_x[23] ? _GEN7939 : _GEN7936;
wire  _GEN7941 = io_x[18] ? _GEN7940 : _GEN7935;
wire  _GEN7942 = io_x[33] ? _GEN7941 : _GEN7928;
wire  _GEN7943 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7944 = io_x[19] ? _GEN7273 : _GEN7943;
wire  _GEN7945 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN7946 = io_x[19] ? _GEN7280 : _GEN7945;
wire  _GEN7947 = io_x[23] ? _GEN7946 : _GEN7944;
wire  _GEN7948 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7949 = io_x[27] ? _GEN7948 : _GEN7278;
wire  _GEN7950 = io_x[19] ? _GEN7280 : _GEN7949;
wire  _GEN7951 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN7952 = io_x[23] ? _GEN7951 : _GEN7950;
wire  _GEN7953 = io_x[18] ? _GEN7952 : _GEN7947;
wire  _GEN7954 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7955 = io_x[27] ? _GEN7954 : _GEN7278;
wire  _GEN7956 = io_x[19] ? _GEN7273 : _GEN7955;
wire  _GEN7957 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7958 = io_x[27] ? _GEN7957 : _GEN7278;
wire  _GEN7959 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7960 = io_x[27] ? _GEN7959 : _GEN7278;
wire  _GEN7961 = io_x[19] ? _GEN7960 : _GEN7958;
wire  _GEN7962 = io_x[23] ? _GEN7961 : _GEN7956;
wire  _GEN7963 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7964 = io_x[27] ? _GEN7963 : _GEN7278;
wire  _GEN7965 = io_x[19] ? _GEN7280 : _GEN7964;
wire  _GEN7966 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7967 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7968 = io_x[27] ? _GEN7967 : _GEN7966;
wire  _GEN7969 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7970 = io_x[27] ? _GEN7969 : _GEN7278;
wire  _GEN7971 = io_x[19] ? _GEN7970 : _GEN7968;
wire  _GEN7972 = io_x[23] ? _GEN7971 : _GEN7965;
wire  _GEN7973 = io_x[18] ? _GEN7972 : _GEN7962;
wire  _GEN7974 = io_x[33] ? _GEN7973 : _GEN7953;
wire  _GEN7975 = io_x[31] ? _GEN7974 : _GEN7942;
wire  _GEN7976 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7977 = io_x[19] ? _GEN7976 : _GEN7280;
wire  _GEN7978 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7979 = io_x[27] ? _GEN7978 : _GEN7278;
wire  _GEN7980 = io_x[19] ? _GEN7280 : _GEN7979;
wire  _GEN7981 = io_x[23] ? _GEN7980 : _GEN7977;
wire  _GEN7982 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7983 = io_x[27] ? _GEN7982 : _GEN7278;
wire  _GEN7984 = io_x[19] ? _GEN7983 : _GEN7280;
wire  _GEN7985 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7986 = io_x[19] ? _GEN7985 : _GEN7273;
wire  _GEN7987 = io_x[23] ? _GEN7986 : _GEN7984;
wire  _GEN7988 = io_x[18] ? _GEN7987 : _GEN7981;
wire  _GEN7989 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN7990 = io_x[19] ? _GEN7989 : _GEN7280;
wire  _GEN7991 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN7992 = io_x[27] ? _GEN7991 : _GEN7278;
wire  _GEN7993 = io_x[19] ? _GEN7992 : _GEN7273;
wire  _GEN7994 = io_x[23] ? _GEN7993 : _GEN7990;
wire  _GEN7995 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7996 = io_x[27] ? _GEN7995 : _GEN7271;
wire  _GEN7997 = io_x[19] ? _GEN7996 : _GEN7280;
wire  _GEN7998 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN7999 = io_x[27] ? _GEN7998 : _GEN7278;
wire  _GEN8000 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8001 = io_x[27] ? _GEN8000 : _GEN7271;
wire  _GEN8002 = io_x[19] ? _GEN8001 : _GEN7999;
wire  _GEN8003 = io_x[23] ? _GEN8002 : _GEN7997;
wire  _GEN8004 = io_x[18] ? _GEN8003 : _GEN7994;
wire  _GEN8005 = io_x[33] ? _GEN8004 : _GEN7988;
wire  _GEN8006 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8007 = io_x[27] ? _GEN7278 : _GEN8006;
wire  _GEN8008 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8009 = io_x[19] ? _GEN8008 : _GEN8007;
wire  _GEN8010 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8011 = io_x[27] ? _GEN8010 : _GEN7278;
wire  _GEN8012 = io_x[19] ? _GEN7273 : _GEN8011;
wire  _GEN8013 = io_x[23] ? _GEN8012 : _GEN8009;
wire  _GEN8014 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8015 = io_x[27] ? _GEN7271 : _GEN8014;
wire  _GEN8016 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8017 = io_x[27] ? _GEN8016 : _GEN7278;
wire  _GEN8018 = io_x[19] ? _GEN8017 : _GEN8015;
wire  _GEN8019 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8020 = io_x[27] ? _GEN7271 : _GEN8019;
wire  _GEN8021 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8022 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8023 = io_x[27] ? _GEN8022 : _GEN8021;
wire  _GEN8024 = io_x[19] ? _GEN8023 : _GEN8020;
wire  _GEN8025 = io_x[23] ? _GEN8024 : _GEN8018;
wire  _GEN8026 = io_x[18] ? _GEN8025 : _GEN8013;
wire  _GEN8027 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8028 = io_x[27] ? _GEN7278 : _GEN8027;
wire  _GEN8029 = io_x[19] ? _GEN8028 : _GEN7280;
wire  _GEN8030 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8031 = io_x[27] ? _GEN8030 : _GEN7278;
wire  _GEN8032 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8033 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8034 = io_x[27] ? _GEN8033 : _GEN8032;
wire  _GEN8035 = io_x[19] ? _GEN8034 : _GEN8031;
wire  _GEN8036 = io_x[23] ? _GEN8035 : _GEN8029;
wire  _GEN8037 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8038 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8039 = io_x[27] ? _GEN8038 : _GEN8037;
wire  _GEN8040 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8041 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8042 = io_x[27] ? _GEN8041 : _GEN8040;
wire  _GEN8043 = io_x[19] ? _GEN8042 : _GEN8039;
wire  _GEN8044 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8045 = io_x[27] ? _GEN8044 : _GEN7278;
wire  _GEN8046 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8047 = io_x[27] ? _GEN8046 : _GEN7278;
wire  _GEN8048 = io_x[19] ? _GEN8047 : _GEN8045;
wire  _GEN8049 = io_x[23] ? _GEN8048 : _GEN8043;
wire  _GEN8050 = io_x[18] ? _GEN8049 : _GEN8036;
wire  _GEN8051 = io_x[33] ? _GEN8050 : _GEN8026;
wire  _GEN8052 = io_x[31] ? _GEN8051 : _GEN8005;
wire  _GEN8053 = io_x[28] ? _GEN8052 : _GEN7975;
wire  _GEN8054 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8055 = io_x[27] ? _GEN8054 : _GEN7278;
wire  _GEN8056 = io_x[19] ? _GEN8055 : _GEN7280;
wire  _GEN8057 = io_x[23] ? _GEN8056 : _GEN7267;
wire  _GEN8058 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8059 = io_x[27] ? _GEN8058 : _GEN7278;
wire  _GEN8060 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8061 = io_x[27] ? _GEN8060 : _GEN7278;
wire  _GEN8062 = io_x[19] ? _GEN8061 : _GEN8059;
wire  _GEN8063 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8064 = io_x[27] ? _GEN7271 : _GEN8063;
wire  _GEN8065 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8066 = io_x[19] ? _GEN8065 : _GEN8064;
wire  _GEN8067 = io_x[23] ? _GEN8066 : _GEN8062;
wire  _GEN8068 = io_x[18] ? _GEN8067 : _GEN8057;
wire  _GEN8069 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8070 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8071 = io_x[27] ? _GEN8070 : _GEN8069;
wire  _GEN8072 = io_x[19] ? _GEN8071 : _GEN7273;
wire  _GEN8073 = io_x[23] ? _GEN7305 : _GEN8072;
wire  _GEN8074 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8075 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8076 = io_x[27] ? _GEN8075 : _GEN8074;
wire  _GEN8077 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8078 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8079 = io_x[27] ? _GEN8078 : _GEN8077;
wire  _GEN8080 = io_x[19] ? _GEN8079 : _GEN8076;
wire  _GEN8081 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8082 = io_x[27] ? _GEN7271 : _GEN8081;
wire  _GEN8083 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8084 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8085 = io_x[27] ? _GEN8084 : _GEN8083;
wire  _GEN8086 = io_x[19] ? _GEN8085 : _GEN8082;
wire  _GEN8087 = io_x[23] ? _GEN8086 : _GEN8080;
wire  _GEN8088 = io_x[18] ? _GEN8087 : _GEN8073;
wire  _GEN8089 = io_x[33] ? _GEN8088 : _GEN8068;
wire  _GEN8090 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8091 = io_x[27] ? _GEN7271 : _GEN8090;
wire  _GEN8092 = io_x[19] ? _GEN8091 : _GEN7280;
wire  _GEN8093 = io_x[23] ? _GEN7267 : _GEN8092;
wire  _GEN8094 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8095 = io_x[27] ? _GEN8094 : _GEN7278;
wire  _GEN8096 = io_x[19] ? _GEN8095 : _GEN7280;
wire  _GEN8097 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8098 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8099 = io_x[27] ? _GEN8098 : _GEN7271;
wire  _GEN8100 = io_x[19] ? _GEN8099 : _GEN8097;
wire  _GEN8101 = io_x[23] ? _GEN8100 : _GEN8096;
wire  _GEN8102 = io_x[18] ? _GEN8101 : _GEN8093;
wire  _GEN8103 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8104 = io_x[27] ? _GEN8103 : _GEN7278;
wire  _GEN8105 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8106 = io_x[27] ? _GEN7271 : _GEN8105;
wire  _GEN8107 = io_x[19] ? _GEN8106 : _GEN8104;
wire  _GEN8108 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8109 = io_x[27] ? _GEN8108 : _GEN7278;
wire  _GEN8110 = io_x[19] ? _GEN8109 : _GEN7273;
wire  _GEN8111 = io_x[23] ? _GEN8110 : _GEN8107;
wire  _GEN8112 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8113 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8114 = io_x[27] ? _GEN8113 : _GEN8112;
wire  _GEN8115 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8116 = io_x[27] ? _GEN8115 : _GEN7278;
wire  _GEN8117 = io_x[19] ? _GEN8116 : _GEN8114;
wire  _GEN8118 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8119 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8120 = io_x[27] ? _GEN8119 : _GEN8118;
wire  _GEN8121 = io_x[19] ? _GEN8120 : _GEN7280;
wire  _GEN8122 = io_x[23] ? _GEN8121 : _GEN8117;
wire  _GEN8123 = io_x[18] ? _GEN8122 : _GEN8111;
wire  _GEN8124 = io_x[33] ? _GEN8123 : _GEN8102;
wire  _GEN8125 = io_x[31] ? _GEN8124 : _GEN8089;
wire  _GEN8126 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8127 = io_x[27] ? _GEN8126 : _GEN7271;
wire  _GEN8128 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8129 = io_x[27] ? _GEN7278 : _GEN8128;
wire  _GEN8130 = io_x[19] ? _GEN8129 : _GEN8127;
wire  _GEN8131 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8132 = io_x[27] ? _GEN8131 : _GEN7278;
wire  _GEN8133 = io_x[19] ? _GEN7280 : _GEN8132;
wire  _GEN8134 = io_x[23] ? _GEN8133 : _GEN8130;
wire  _GEN8135 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8136 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8137 = io_x[27] ? _GEN8136 : _GEN8135;
wire  _GEN8138 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8139 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8140 = io_x[27] ? _GEN8139 : _GEN8138;
wire  _GEN8141 = io_x[19] ? _GEN8140 : _GEN8137;
wire  _GEN8142 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8143 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8144 = io_x[27] ? _GEN8143 : _GEN8142;
wire  _GEN8145 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8146 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8147 = io_x[27] ? _GEN8146 : _GEN8145;
wire  _GEN8148 = io_x[19] ? _GEN8147 : _GEN8144;
wire  _GEN8149 = io_x[23] ? _GEN8148 : _GEN8141;
wire  _GEN8150 = io_x[18] ? _GEN8149 : _GEN8134;
wire  _GEN8151 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8152 = io_x[27] ? _GEN8151 : _GEN7271;
wire  _GEN8153 = io_x[19] ? _GEN8152 : _GEN7273;
wire  _GEN8154 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8155 = io_x[19] ? _GEN8154 : _GEN7280;
wire  _GEN8156 = io_x[23] ? _GEN8155 : _GEN8153;
wire  _GEN8157 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8158 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8159 = io_x[27] ? _GEN8158 : _GEN8157;
wire  _GEN8160 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8161 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8162 = io_x[27] ? _GEN8161 : _GEN8160;
wire  _GEN8163 = io_x[19] ? _GEN8162 : _GEN8159;
wire  _GEN8164 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8165 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8166 = io_x[27] ? _GEN8165 : _GEN8164;
wire  _GEN8167 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8168 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8169 = io_x[27] ? _GEN8168 : _GEN8167;
wire  _GEN8170 = io_x[19] ? _GEN8169 : _GEN8166;
wire  _GEN8171 = io_x[23] ? _GEN8170 : _GEN8163;
wire  _GEN8172 = io_x[18] ? _GEN8171 : _GEN8156;
wire  _GEN8173 = io_x[33] ? _GEN8172 : _GEN8150;
wire  _GEN8174 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8175 = io_x[27] ? _GEN8174 : _GEN7278;
wire  _GEN8176 = io_x[19] ? _GEN8175 : _GEN7280;
wire  _GEN8177 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8178 = io_x[27] ? _GEN8177 : _GEN7278;
wire  _GEN8179 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8180 = io_x[27] ? _GEN8179 : _GEN7278;
wire  _GEN8181 = io_x[19] ? _GEN8180 : _GEN8178;
wire  _GEN8182 = io_x[23] ? _GEN8181 : _GEN8176;
wire  _GEN8183 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8184 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8185 = io_x[27] ? _GEN8184 : _GEN8183;
wire  _GEN8186 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8187 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8188 = io_x[27] ? _GEN8187 : _GEN8186;
wire  _GEN8189 = io_x[19] ? _GEN8188 : _GEN8185;
wire  _GEN8190 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8191 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8192 = io_x[27] ? _GEN8191 : _GEN8190;
wire  _GEN8193 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8194 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8195 = io_x[27] ? _GEN8194 : _GEN8193;
wire  _GEN8196 = io_x[19] ? _GEN8195 : _GEN8192;
wire  _GEN8197 = io_x[23] ? _GEN8196 : _GEN8189;
wire  _GEN8198 = io_x[18] ? _GEN8197 : _GEN8182;
wire  _GEN8199 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8200 = io_x[27] ? _GEN8199 : _GEN7278;
wire  _GEN8201 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8202 = io_x[19] ? _GEN8201 : _GEN8200;
wire  _GEN8203 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8204 = io_x[27] ? _GEN8203 : _GEN7271;
wire  _GEN8205 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8206 = io_x[27] ? _GEN8205 : _GEN7278;
wire  _GEN8207 = io_x[19] ? _GEN8206 : _GEN8204;
wire  _GEN8208 = io_x[23] ? _GEN8207 : _GEN8202;
wire  _GEN8209 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8210 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8211 = io_x[27] ? _GEN8210 : _GEN8209;
wire  _GEN8212 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8213 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8214 = io_x[27] ? _GEN8213 : _GEN8212;
wire  _GEN8215 = io_x[19] ? _GEN8214 : _GEN8211;
wire  _GEN8216 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8217 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8218 = io_x[27] ? _GEN8217 : _GEN8216;
wire  _GEN8219 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8220 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8221 = io_x[27] ? _GEN8220 : _GEN8219;
wire  _GEN8222 = io_x[19] ? _GEN8221 : _GEN8218;
wire  _GEN8223 = io_x[23] ? _GEN8222 : _GEN8215;
wire  _GEN8224 = io_x[18] ? _GEN8223 : _GEN8208;
wire  _GEN8225 = io_x[33] ? _GEN8224 : _GEN8198;
wire  _GEN8226 = io_x[31] ? _GEN8225 : _GEN8173;
wire  _GEN8227 = io_x[28] ? _GEN8226 : _GEN8125;
wire  _GEN8228 = io_x[26] ? _GEN8227 : _GEN8053;
wire  _GEN8229 = io_x[20] ? _GEN8228 : _GEN7915;
wire  _GEN8230 = io_x[24] ? _GEN8229 : _GEN7695;
wire  _GEN8231 = io_x[18] ? _GEN7297 : _GEN7266;
wire  _GEN8232 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8233 = io_x[27] ? _GEN8232 : _GEN7278;
wire  _GEN8234 = io_x[19] ? _GEN8233 : _GEN7280;
wire  _GEN8235 = io_x[23] ? _GEN8234 : _GEN7305;
wire  _GEN8236 = io_x[18] ? _GEN7297 : _GEN8235;
wire  _GEN8237 = io_x[33] ? _GEN8236 : _GEN8231;
wire  _GEN8238 = io_x[23] ? _GEN7267 : _GEN7305;
wire  _GEN8239 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8240 = io_x[27] ? _GEN8239 : _GEN7278;
wire  _GEN8241 = io_x[19] ? _GEN8240 : _GEN7273;
wire  _GEN8242 = io_x[23] ? _GEN8241 : _GEN7267;
wire  _GEN8243 = io_x[18] ? _GEN8242 : _GEN8238;
wire  _GEN8244 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8245 = io_x[19] ? _GEN8244 : _GEN7280;
wire  _GEN8246 = io_x[23] ? _GEN7267 : _GEN8245;
wire  _GEN8247 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8248 = io_x[27] ? _GEN8247 : _GEN7278;
wire  _GEN8249 = io_x[19] ? _GEN8248 : _GEN7280;
wire  _GEN8250 = io_x[23] ? _GEN8249 : _GEN7267;
wire  _GEN8251 = io_x[18] ? _GEN8250 : _GEN8246;
wire  _GEN8252 = io_x[33] ? _GEN8251 : _GEN8243;
wire  _GEN8253 = io_x[31] ? _GEN8252 : _GEN8237;
wire  _GEN8254 = io_x[23] ? _GEN7267 : _GEN7305;
wire  _GEN8255 = io_x[18] ? _GEN8254 : _GEN7266;
wire  _GEN8256 = io_x[23] ? _GEN7267 : _GEN7305;
wire  _GEN8257 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8258 = io_x[19] ? _GEN8257 : _GEN7280;
wire  _GEN8259 = io_x[23] ? _GEN8258 : _GEN7267;
wire  _GEN8260 = io_x[18] ? _GEN8259 : _GEN8256;
wire  _GEN8261 = io_x[33] ? _GEN8260 : _GEN8255;
wire  _GEN8262 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8263 = io_x[19] ? _GEN8262 : _GEN7280;
wire  _GEN8264 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8265 = io_x[19] ? _GEN8264 : _GEN7280;
wire  _GEN8266 = io_x[23] ? _GEN8265 : _GEN8263;
wire  _GEN8267 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8268 = io_x[23] ? _GEN7305 : _GEN8267;
wire  _GEN8269 = io_x[18] ? _GEN8268 : _GEN8266;
wire  _GEN8270 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8271 = io_x[19] ? _GEN8270 : _GEN7280;
wire  _GEN8272 = io_x[23] ? _GEN7267 : _GEN8271;
wire  _GEN8273 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8274 = io_x[23] ? _GEN7305 : _GEN8273;
wire  _GEN8275 = io_x[18] ? _GEN8274 : _GEN8272;
wire  _GEN8276 = io_x[33] ? _GEN8275 : _GEN8269;
wire  _GEN8277 = io_x[31] ? _GEN8276 : _GEN8261;
wire  _GEN8278 = io_x[28] ? _GEN8277 : _GEN8253;
wire  _GEN8279 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8280 = io_x[19] ? _GEN8279 : _GEN7280;
wire  _GEN8281 = io_x[23] ? _GEN8280 : _GEN7305;
wire  _GEN8282 = io_x[18] ? _GEN8281 : _GEN7297;
wire  _GEN8283 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8284 = io_x[19] ? _GEN8283 : _GEN7280;
wire  _GEN8285 = io_x[23] ? _GEN8284 : _GEN7267;
wire  _GEN8286 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8287 = io_x[27] ? _GEN8286 : _GEN7271;
wire  _GEN8288 = io_x[19] ? _GEN8287 : _GEN7280;
wire  _GEN8289 = io_x[23] ? _GEN8288 : _GEN7305;
wire  _GEN8290 = io_x[18] ? _GEN8289 : _GEN8285;
wire  _GEN8291 = io_x[33] ? _GEN8290 : _GEN8282;
wire  _GEN8292 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8293 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8294 = io_x[27] ? _GEN8293 : _GEN8292;
wire  _GEN8295 = io_x[19] ? _GEN8294 : _GEN7280;
wire  _GEN8296 = io_x[23] ? _GEN8295 : _GEN7267;
wire  _GEN8297 = io_x[18] ? _GEN8296 : _GEN7266;
wire  _GEN8298 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN8299 = io_x[23] ? _GEN8298 : _GEN7267;
wire  _GEN8300 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8301 = io_x[19] ? _GEN7280 : _GEN8300;
wire  _GEN8302 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8303 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8304 = io_x[27] ? _GEN8303 : _GEN7278;
wire  _GEN8305 = io_x[19] ? _GEN8304 : _GEN8302;
wire  _GEN8306 = io_x[23] ? _GEN8305 : _GEN8301;
wire  _GEN8307 = io_x[18] ? _GEN8306 : _GEN8299;
wire  _GEN8308 = io_x[33] ? _GEN8307 : _GEN8297;
wire  _GEN8309 = io_x[31] ? _GEN8308 : _GEN8291;
wire  _GEN8310 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8311 = io_x[19] ? _GEN8310 : _GEN7280;
wire  _GEN8312 = io_x[23] ? _GEN7267 : _GEN8311;
wire  _GEN8313 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8314 = io_x[27] ? _GEN7278 : _GEN8313;
wire  _GEN8315 = io_x[19] ? _GEN8314 : _GEN7280;
wire  _GEN8316 = io_x[23] ? _GEN8315 : _GEN7267;
wire  _GEN8317 = io_x[18] ? _GEN8316 : _GEN8312;
wire  _GEN8318 = io_x[18] ? _GEN7266 : _GEN7297;
wire  _GEN8319 = io_x[33] ? _GEN8318 : _GEN8317;
wire  _GEN8320 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8321 = io_x[23] ? _GEN8320 : _GEN7267;
wire  _GEN8322 = io_x[18] ? _GEN8321 : _GEN7297;
wire  _GEN8323 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8324 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8325 = io_x[27] ? _GEN7278 : _GEN8324;
wire  _GEN8326 = io_x[19] ? _GEN8325 : _GEN7280;
wire  _GEN8327 = io_x[23] ? _GEN8326 : _GEN8323;
wire  _GEN8328 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8329 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8330 = io_x[27] ? _GEN8329 : _GEN8328;
wire  _GEN8331 = io_x[19] ? _GEN8330 : _GEN7280;
wire  _GEN8332 = io_x[23] ? _GEN8331 : _GEN7267;
wire  _GEN8333 = io_x[18] ? _GEN8332 : _GEN8327;
wire  _GEN8334 = io_x[33] ? _GEN8333 : _GEN8322;
wire  _GEN8335 = io_x[31] ? _GEN8334 : _GEN8319;
wire  _GEN8336 = io_x[28] ? _GEN8335 : _GEN8309;
wire  _GEN8337 = io_x[26] ? _GEN8336 : _GEN8278;
wire  _GEN8338 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8339 = io_x[19] ? _GEN8338 : _GEN7280;
wire  _GEN8340 = io_x[23] ? _GEN8339 : _GEN7267;
wire  _GEN8341 = io_x[18] ? _GEN7266 : _GEN8340;
wire  _GEN8342 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8343 = io_x[23] ? _GEN8342 : _GEN7267;
wire  _GEN8344 = io_x[18] ? _GEN8343 : _GEN7297;
wire  _GEN8345 = io_x[33] ? _GEN8344 : _GEN8341;
wire  _GEN8346 = 1'b0;
wire  _GEN8347 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8348 = io_x[27] ? _GEN8347 : _GEN7278;
wire  _GEN8349 = io_x[19] ? _GEN8348 : _GEN7273;
wire  _GEN8350 = io_x[23] ? _GEN8349 : _GEN7305;
wire  _GEN8351 = io_x[18] ? _GEN8350 : _GEN7297;
wire  _GEN8352 = io_x[33] ? _GEN8351 : _GEN8346;
wire  _GEN8353 = io_x[31] ? _GEN8352 : _GEN8345;
wire  _GEN8354 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8355 = io_x[19] ? _GEN7280 : _GEN8354;
wire  _GEN8356 = io_x[23] ? _GEN8355 : _GEN7267;
wire  _GEN8357 = io_x[18] ? _GEN7297 : _GEN8356;
wire  _GEN8358 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8359 = io_x[19] ? _GEN7273 : _GEN8358;
wire  _GEN8360 = io_x[23] ? _GEN8359 : _GEN7267;
wire  _GEN8361 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN8362 = io_x[18] ? _GEN8361 : _GEN8360;
wire  _GEN8363 = io_x[33] ? _GEN8362 : _GEN8357;
wire  _GEN8364 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8365 = io_x[27] ? _GEN8364 : _GEN7271;
wire  _GEN8366 = io_x[19] ? _GEN7280 : _GEN8365;
wire  _GEN8367 = io_x[23] ? _GEN8366 : _GEN7267;
wire  _GEN8368 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8369 = io_x[19] ? _GEN8368 : _GEN7280;
wire  _GEN8370 = io_x[23] ? _GEN8369 : _GEN7305;
wire  _GEN8371 = io_x[18] ? _GEN8370 : _GEN8367;
wire  _GEN8372 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8373 = io_x[19] ? _GEN7280 : _GEN8372;
wire  _GEN8374 = io_x[23] ? _GEN8373 : _GEN7267;
wire  _GEN8375 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8376 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8377 = io_x[27] ? _GEN8376 : _GEN8375;
wire  _GEN8378 = io_x[19] ? _GEN8377 : _GEN7280;
wire  _GEN8379 = io_x[23] ? _GEN8378 : _GEN7305;
wire  _GEN8380 = io_x[18] ? _GEN8379 : _GEN8374;
wire  _GEN8381 = io_x[33] ? _GEN8380 : _GEN8371;
wire  _GEN8382 = io_x[31] ? _GEN8381 : _GEN8363;
wire  _GEN8383 = io_x[28] ? _GEN8382 : _GEN8353;
wire  _GEN8384 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8385 = io_x[27] ? _GEN7271 : _GEN8384;
wire  _GEN8386 = io_x[19] ? _GEN7280 : _GEN8385;
wire  _GEN8387 = io_x[23] ? _GEN8386 : _GEN7267;
wire  _GEN8388 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8389 = io_x[27] ? _GEN8388 : _GEN7271;
wire  _GEN8390 = io_x[19] ? _GEN8389 : _GEN7280;
wire  _GEN8391 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8392 = io_x[27] ? _GEN8391 : _GEN7278;
wire  _GEN8393 = io_x[19] ? _GEN8392 : _GEN7280;
wire  _GEN8394 = io_x[23] ? _GEN8393 : _GEN8390;
wire  _GEN8395 = io_x[18] ? _GEN8394 : _GEN8387;
wire  _GEN8396 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8397 = io_x[27] ? _GEN7278 : _GEN8396;
wire  _GEN8398 = io_x[19] ? _GEN8397 : _GEN7280;
wire  _GEN8399 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8400 = io_x[27] ? _GEN7271 : _GEN8399;
wire  _GEN8401 = io_x[19] ? _GEN7280 : _GEN8400;
wire  _GEN8402 = io_x[23] ? _GEN8401 : _GEN8398;
wire  _GEN8403 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8404 = io_x[27] ? _GEN8403 : _GEN7278;
wire  _GEN8405 = io_x[19] ? _GEN8404 : _GEN7280;
wire  _GEN8406 = io_x[23] ? _GEN7267 : _GEN8405;
wire  _GEN8407 = io_x[18] ? _GEN8406 : _GEN8402;
wire  _GEN8408 = io_x[33] ? _GEN8407 : _GEN8395;
wire  _GEN8409 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN8410 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8411 = io_x[27] ? _GEN8410 : _GEN7278;
wire  _GEN8412 = io_x[19] ? _GEN8411 : _GEN7280;
wire  _GEN8413 = io_x[23] ? _GEN8412 : _GEN7267;
wire  _GEN8414 = io_x[18] ? _GEN8413 : _GEN8409;
wire  _GEN8415 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8416 = io_x[19] ? _GEN7273 : _GEN8415;
wire  _GEN8417 = io_x[23] ? _GEN8416 : _GEN7267;
wire  _GEN8418 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8419 = io_x[27] ? _GEN8418 : _GEN7278;
wire  _GEN8420 = io_x[19] ? _GEN8419 : _GEN7280;
wire  _GEN8421 = io_x[23] ? _GEN8420 : _GEN7267;
wire  _GEN8422 = io_x[18] ? _GEN8421 : _GEN8417;
wire  _GEN8423 = io_x[33] ? _GEN8422 : _GEN8414;
wire  _GEN8424 = io_x[31] ? _GEN8423 : _GEN8408;
wire  _GEN8425 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8426 = io_x[23] ? _GEN8425 : _GEN7267;
wire  _GEN8427 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN8428 = io_x[18] ? _GEN8427 : _GEN8426;
wire  _GEN8429 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8430 = io_x[23] ? _GEN8429 : _GEN7267;
wire  _GEN8431 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8432 = io_x[27] ? _GEN7271 : _GEN8431;
wire  _GEN8433 = io_x[19] ? _GEN8432 : _GEN7280;
wire  _GEN8434 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8435 = io_x[19] ? _GEN8434 : _GEN7280;
wire  _GEN8436 = io_x[23] ? _GEN8435 : _GEN8433;
wire  _GEN8437 = io_x[18] ? _GEN8436 : _GEN8430;
wire  _GEN8438 = io_x[33] ? _GEN8437 : _GEN8428;
wire  _GEN8439 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN8440 = io_x[23] ? _GEN8439 : _GEN7267;
wire  _GEN8441 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8442 = io_x[27] ? _GEN8441 : _GEN7271;
wire  _GEN8443 = io_x[19] ? _GEN7273 : _GEN8442;
wire  _GEN8444 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8445 = io_x[27] ? _GEN8444 : _GEN7278;
wire  _GEN8446 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8447 = io_x[27] ? _GEN8446 : _GEN7278;
wire  _GEN8448 = io_x[19] ? _GEN8447 : _GEN8445;
wire  _GEN8449 = io_x[23] ? _GEN8448 : _GEN8443;
wire  _GEN8450 = io_x[18] ? _GEN8449 : _GEN8440;
wire  _GEN8451 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN8452 = io_x[23] ? _GEN8451 : _GEN7267;
wire  _GEN8453 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8454 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8455 = io_x[27] ? _GEN8454 : _GEN8453;
wire  _GEN8456 = io_x[19] ? _GEN8455 : _GEN7280;
wire  _GEN8457 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8458 = io_x[27] ? _GEN8457 : _GEN7278;
wire  _GEN8459 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8460 = io_x[27] ? _GEN8459 : _GEN7278;
wire  _GEN8461 = io_x[19] ? _GEN8460 : _GEN8458;
wire  _GEN8462 = io_x[23] ? _GEN8461 : _GEN8456;
wire  _GEN8463 = io_x[18] ? _GEN8462 : _GEN8452;
wire  _GEN8464 = io_x[33] ? _GEN8463 : _GEN8450;
wire  _GEN8465 = io_x[31] ? _GEN8464 : _GEN8438;
wire  _GEN8466 = io_x[28] ? _GEN8465 : _GEN8424;
wire  _GEN8467 = io_x[26] ? _GEN8466 : _GEN8383;
wire  _GEN8468 = io_x[20] ? _GEN8467 : _GEN8337;
wire  _GEN8469 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8470 = io_x[27] ? _GEN8469 : _GEN7278;
wire  _GEN8471 = io_x[19] ? _GEN8470 : _GEN7273;
wire  _GEN8472 = io_x[23] ? _GEN7267 : _GEN8471;
wire  _GEN8473 = io_x[18] ? _GEN8472 : _GEN7297;
wire  _GEN8474 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8475 = io_x[19] ? _GEN7273 : _GEN8474;
wire  _GEN8476 = io_x[23] ? _GEN7267 : _GEN8475;
wire  _GEN8477 = io_x[18] ? _GEN8476 : _GEN7266;
wire  _GEN8478 = io_x[33] ? _GEN8477 : _GEN8473;
wire  _GEN8479 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN8480 = io_x[18] ? _GEN8479 : _GEN7266;
wire  _GEN8481 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8482 = io_x[27] ? _GEN8481 : _GEN7278;
wire  _GEN8483 = io_x[19] ? _GEN8482 : _GEN7280;
wire  _GEN8484 = io_x[23] ? _GEN8483 : _GEN7305;
wire  _GEN8485 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8486 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8487 = io_x[27] ? _GEN8486 : _GEN7278;
wire  _GEN8488 = io_x[19] ? _GEN8487 : _GEN8485;
wire  _GEN8489 = io_x[23] ? _GEN7305 : _GEN8488;
wire  _GEN8490 = io_x[18] ? _GEN8489 : _GEN8484;
wire  _GEN8491 = io_x[33] ? _GEN8490 : _GEN8480;
wire  _GEN8492 = io_x[31] ? _GEN8491 : _GEN8478;
wire  _GEN8493 = io_x[18] ? _GEN7266 : _GEN7297;
wire  _GEN8494 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8495 = io_x[27] ? _GEN8494 : _GEN7278;
wire  _GEN8496 = io_x[19] ? _GEN8495 : _GEN7273;
wire  _GEN8497 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8498 = io_x[19] ? _GEN8497 : _GEN7280;
wire  _GEN8499 = io_x[23] ? _GEN8498 : _GEN8496;
wire  _GEN8500 = io_x[18] ? _GEN8499 : _GEN7297;
wire  _GEN8501 = io_x[33] ? _GEN8500 : _GEN8493;
wire  _GEN8502 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8503 = io_x[23] ? _GEN7267 : _GEN8502;
wire  _GEN8504 = io_x[18] ? _GEN8503 : _GEN7266;
wire  _GEN8505 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8506 = io_x[27] ? _GEN8505 : _GEN7278;
wire  _GEN8507 = io_x[19] ? _GEN8506 : _GEN7280;
wire  _GEN8508 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8509 = io_x[19] ? _GEN8508 : _GEN7280;
wire  _GEN8510 = io_x[23] ? _GEN8509 : _GEN8507;
wire  _GEN8511 = io_x[18] ? _GEN8510 : _GEN7297;
wire  _GEN8512 = io_x[33] ? _GEN8511 : _GEN8504;
wire  _GEN8513 = io_x[31] ? _GEN8512 : _GEN8501;
wire  _GEN8514 = io_x[28] ? _GEN8513 : _GEN8492;
wire  _GEN8515 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN8516 = io_x[23] ? _GEN7305 : _GEN8515;
wire  _GEN8517 = io_x[18] ? _GEN8516 : _GEN7266;
wire  _GEN8518 = io_x[33] ? _GEN8346 : _GEN8517;
wire  _GEN8519 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8520 = io_x[19] ? _GEN8519 : _GEN7280;
wire  _GEN8521 = io_x[23] ? _GEN8520 : _GEN7267;
wire  _GEN8522 = io_x[18] ? _GEN8521 : _GEN7297;
wire  _GEN8523 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8524 = io_x[19] ? _GEN8523 : _GEN7280;
wire  _GEN8525 = io_x[23] ? _GEN8524 : _GEN7267;
wire  _GEN8526 = io_x[18] ? _GEN8525 : _GEN7266;
wire  _GEN8527 = io_x[33] ? _GEN8526 : _GEN8522;
wire  _GEN8528 = io_x[31] ? _GEN8527 : _GEN8518;
wire  _GEN8529 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8530 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8531 = io_x[27] ? _GEN8530 : _GEN7278;
wire  _GEN8532 = io_x[19] ? _GEN8531 : _GEN7280;
wire  _GEN8533 = io_x[23] ? _GEN8532 : _GEN8529;
wire  _GEN8534 = io_x[18] ? _GEN8533 : _GEN7297;
wire  _GEN8535 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8536 = io_x[19] ? _GEN7280 : _GEN8535;
wire  _GEN8537 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8538 = io_x[27] ? _GEN8537 : _GEN7278;
wire  _GEN8539 = io_x[19] ? _GEN8538 : _GEN7280;
wire  _GEN8540 = io_x[23] ? _GEN8539 : _GEN8536;
wire  _GEN8541 = io_x[18] ? _GEN8540 : _GEN7297;
wire  _GEN8542 = io_x[33] ? _GEN8541 : _GEN8534;
wire  _GEN8543 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8544 = io_x[27] ? _GEN8543 : _GEN7278;
wire  _GEN8545 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8546 = io_x[27] ? _GEN8545 : _GEN7278;
wire  _GEN8547 = io_x[19] ? _GEN8546 : _GEN8544;
wire  _GEN8548 = io_x[23] ? _GEN8547 : _GEN7305;
wire  _GEN8549 = io_x[18] ? _GEN7266 : _GEN8548;
wire  _GEN8550 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8551 = io_x[27] ? _GEN8550 : _GEN7278;
wire  _GEN8552 = io_x[19] ? _GEN7280 : _GEN8551;
wire  _GEN8553 = io_x[23] ? _GEN8552 : _GEN7305;
wire  _GEN8554 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8555 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8556 = io_x[27] ? _GEN8555 : _GEN8554;
wire  _GEN8557 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8558 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8559 = io_x[27] ? _GEN8558 : _GEN8557;
wire  _GEN8560 = io_x[19] ? _GEN8559 : _GEN8556;
wire  _GEN8561 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8562 = io_x[27] ? _GEN8561 : _GEN7278;
wire  _GEN8563 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8564 = io_x[27] ? _GEN8563 : _GEN7278;
wire  _GEN8565 = io_x[19] ? _GEN8564 : _GEN8562;
wire  _GEN8566 = io_x[23] ? _GEN8565 : _GEN8560;
wire  _GEN8567 = io_x[18] ? _GEN8566 : _GEN8553;
wire  _GEN8568 = io_x[33] ? _GEN8567 : _GEN8549;
wire  _GEN8569 = io_x[31] ? _GEN8568 : _GEN8542;
wire  _GEN8570 = io_x[28] ? _GEN8569 : _GEN8528;
wire  _GEN8571 = io_x[26] ? _GEN8570 : _GEN8514;
wire  _GEN8572 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8573 = io_x[19] ? _GEN7280 : _GEN8572;
wire  _GEN8574 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8575 = io_x[23] ? _GEN8574 : _GEN8573;
wire  _GEN8576 = io_x[18] ? _GEN7297 : _GEN8575;
wire  _GEN8577 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8578 = io_x[19] ? _GEN7280 : _GEN8577;
wire  _GEN8579 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8580 = io_x[23] ? _GEN8579 : _GEN8578;
wire  _GEN8581 = io_x[18] ? _GEN7266 : _GEN8580;
wire  _GEN8582 = io_x[33] ? _GEN8581 : _GEN8576;
wire  _GEN8583 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8584 = io_x[23] ? _GEN7267 : _GEN8583;
wire  _GEN8585 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8586 = io_x[27] ? _GEN8585 : _GEN7278;
wire  _GEN8587 = io_x[19] ? _GEN8586 : _GEN7280;
wire  _GEN8588 = io_x[23] ? _GEN8587 : _GEN7267;
wire  _GEN8589 = io_x[18] ? _GEN8588 : _GEN8584;
wire  _GEN8590 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8591 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8592 = io_x[27] ? _GEN8591 : _GEN7278;
wire  _GEN8593 = io_x[19] ? _GEN8592 : _GEN7280;
wire  _GEN8594 = io_x[23] ? _GEN8593 : _GEN8590;
wire  _GEN8595 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8596 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8597 = io_x[27] ? _GEN8596 : _GEN8595;
wire  _GEN8598 = io_x[19] ? _GEN8597 : _GEN7273;
wire  _GEN8599 = io_x[23] ? _GEN8598 : _GEN7267;
wire  _GEN8600 = io_x[18] ? _GEN8599 : _GEN8594;
wire  _GEN8601 = io_x[33] ? _GEN8600 : _GEN8589;
wire  _GEN8602 = io_x[31] ? _GEN8601 : _GEN8582;
wire  _GEN8603 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8604 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8605 = io_x[27] ? _GEN7271 : _GEN8604;
wire  _GEN8606 = io_x[19] ? _GEN8605 : _GEN8603;
wire  _GEN8607 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8608 = io_x[23] ? _GEN8607 : _GEN8606;
wire  _GEN8609 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8610 = io_x[19] ? _GEN8609 : _GEN7273;
wire  _GEN8611 = io_x[23] ? _GEN8610 : _GEN7305;
wire  _GEN8612 = io_x[18] ? _GEN8611 : _GEN8608;
wire  _GEN8613 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8614 = io_x[27] ? _GEN7278 : _GEN8613;
wire  _GEN8615 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8616 = io_x[19] ? _GEN8615 : _GEN8614;
wire  _GEN8617 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8618 = io_x[27] ? _GEN8617 : _GEN7271;
wire  _GEN8619 = io_x[19] ? _GEN8618 : _GEN7273;
wire  _GEN8620 = io_x[23] ? _GEN8619 : _GEN8616;
wire  _GEN8621 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8622 = io_x[27] ? _GEN8621 : _GEN7278;
wire  _GEN8623 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8624 = io_x[27] ? _GEN8623 : _GEN7278;
wire  _GEN8625 = io_x[19] ? _GEN8624 : _GEN8622;
wire  _GEN8626 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8627 = io_x[23] ? _GEN8626 : _GEN8625;
wire  _GEN8628 = io_x[18] ? _GEN8627 : _GEN8620;
wire  _GEN8629 = io_x[33] ? _GEN8628 : _GEN8612;
wire  _GEN8630 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8631 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8632 = io_x[27] ? _GEN8631 : _GEN7278;
wire  _GEN8633 = io_x[19] ? _GEN8632 : _GEN7280;
wire  _GEN8634 = io_x[23] ? _GEN8633 : _GEN8630;
wire  _GEN8635 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8636 = io_x[27] ? _GEN7278 : _GEN8635;
wire  _GEN8637 = io_x[19] ? _GEN8636 : _GEN7273;
wire  _GEN8638 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8639 = io_x[27] ? _GEN8638 : _GEN7278;
wire  _GEN8640 = io_x[19] ? _GEN8639 : _GEN7280;
wire  _GEN8641 = io_x[23] ? _GEN8640 : _GEN8637;
wire  _GEN8642 = io_x[18] ? _GEN8641 : _GEN8634;
wire  _GEN8643 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8644 = io_x[19] ? _GEN8643 : _GEN7273;
wire  _GEN8645 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8646 = io_x[27] ? _GEN8645 : _GEN7278;
wire  _GEN8647 = io_x[19] ? _GEN8646 : _GEN7280;
wire  _GEN8648 = io_x[23] ? _GEN8647 : _GEN8644;
wire  _GEN8649 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8650 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8651 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8652 = io_x[27] ? _GEN8651 : _GEN8650;
wire  _GEN8653 = io_x[19] ? _GEN8652 : _GEN7280;
wire  _GEN8654 = io_x[23] ? _GEN8653 : _GEN8649;
wire  _GEN8655 = io_x[18] ? _GEN8654 : _GEN8648;
wire  _GEN8656 = io_x[33] ? _GEN8655 : _GEN8642;
wire  _GEN8657 = io_x[31] ? _GEN8656 : _GEN8629;
wire  _GEN8658 = io_x[28] ? _GEN8657 : _GEN8602;
wire  _GEN8659 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8660 = io_x[27] ? _GEN8659 : _GEN7278;
wire  _GEN8661 = io_x[19] ? _GEN8660 : _GEN7280;
wire  _GEN8662 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8663 = io_x[19] ? _GEN8662 : _GEN7280;
wire  _GEN8664 = io_x[23] ? _GEN8663 : _GEN8661;
wire  _GEN8665 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8666 = io_x[27] ? _GEN7278 : _GEN8665;
wire  _GEN8667 = io_x[19] ? _GEN8666 : _GEN7280;
wire  _GEN8668 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8669 = io_x[27] ? _GEN8668 : _GEN7278;
wire  _GEN8670 = io_x[19] ? _GEN8669 : _GEN7280;
wire  _GEN8671 = io_x[23] ? _GEN8670 : _GEN8667;
wire  _GEN8672 = io_x[18] ? _GEN8671 : _GEN8664;
wire  _GEN8673 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8674 = io_x[19] ? _GEN7273 : _GEN8673;
wire  _GEN8675 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8676 = io_x[27] ? _GEN8675 : _GEN7278;
wire  _GEN8677 = io_x[19] ? _GEN8676 : _GEN7280;
wire  _GEN8678 = io_x[23] ? _GEN8677 : _GEN8674;
wire  _GEN8679 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8680 = io_x[27] ? _GEN7271 : _GEN8679;
wire  _GEN8681 = io_x[19] ? _GEN8680 : _GEN7280;
wire  _GEN8682 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8683 = io_x[27] ? _GEN8682 : _GEN7278;
wire  _GEN8684 = io_x[19] ? _GEN8683 : _GEN7280;
wire  _GEN8685 = io_x[23] ? _GEN8684 : _GEN8681;
wire  _GEN8686 = io_x[18] ? _GEN8685 : _GEN8678;
wire  _GEN8687 = io_x[33] ? _GEN8686 : _GEN8672;
wire  _GEN8688 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8689 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8690 = io_x[27] ? _GEN8689 : _GEN7278;
wire  _GEN8691 = io_x[19] ? _GEN8690 : _GEN8688;
wire  _GEN8692 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8693 = io_x[27] ? _GEN8692 : _GEN7278;
wire  _GEN8694 = io_x[19] ? _GEN8693 : _GEN7280;
wire  _GEN8695 = io_x[23] ? _GEN8694 : _GEN8691;
wire  _GEN8696 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8697 = io_x[27] ? _GEN8696 : _GEN7278;
wire  _GEN8698 = io_x[19] ? _GEN7273 : _GEN8697;
wire  _GEN8699 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8700 = io_x[27] ? _GEN8699 : _GEN7278;
wire  _GEN8701 = io_x[19] ? _GEN8700 : _GEN7273;
wire  _GEN8702 = io_x[23] ? _GEN8701 : _GEN8698;
wire  _GEN8703 = io_x[18] ? _GEN8702 : _GEN8695;
wire  _GEN8704 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8705 = io_x[27] ? _GEN8704 : _GEN7278;
wire  _GEN8706 = io_x[19] ? _GEN8705 : _GEN7273;
wire  _GEN8707 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8708 = io_x[27] ? _GEN8707 : _GEN7278;
wire  _GEN8709 = io_x[19] ? _GEN8708 : _GEN7280;
wire  _GEN8710 = io_x[23] ? _GEN8709 : _GEN8706;
wire  _GEN8711 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN8712 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8713 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8714 = io_x[27] ? _GEN8713 : _GEN8712;
wire  _GEN8715 = io_x[19] ? _GEN8714 : _GEN7280;
wire  _GEN8716 = io_x[23] ? _GEN8715 : _GEN8711;
wire  _GEN8717 = io_x[18] ? _GEN8716 : _GEN8710;
wire  _GEN8718 = io_x[33] ? _GEN8717 : _GEN8703;
wire  _GEN8719 = io_x[31] ? _GEN8718 : _GEN8687;
wire  _GEN8720 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8721 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8722 = io_x[27] ? _GEN7271 : _GEN8721;
wire  _GEN8723 = io_x[19] ? _GEN8722 : _GEN8720;
wire  _GEN8724 = io_x[23] ? _GEN8723 : _GEN7305;
wire  _GEN8725 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8726 = io_x[27] ? _GEN7278 : _GEN8725;
wire  _GEN8727 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8728 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8729 = io_x[27] ? _GEN8728 : _GEN8727;
wire  _GEN8730 = io_x[19] ? _GEN8729 : _GEN8726;
wire  _GEN8731 = io_x[23] ? _GEN8730 : _GEN7267;
wire  _GEN8732 = io_x[18] ? _GEN8731 : _GEN8724;
wire  _GEN8733 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8734 = io_x[19] ? _GEN7273 : _GEN8733;
wire  _GEN8735 = io_x[23] ? _GEN7305 : _GEN8734;
wire  _GEN8736 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8737 = io_x[27] ? _GEN7278 : _GEN8736;
wire  _GEN8738 = io_x[19] ? _GEN8737 : _GEN7280;
wire  _GEN8739 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8740 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8741 = io_x[27] ? _GEN8740 : _GEN8739;
wire  _GEN8742 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8743 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8744 = io_x[27] ? _GEN8743 : _GEN8742;
wire  _GEN8745 = io_x[19] ? _GEN8744 : _GEN8741;
wire  _GEN8746 = io_x[23] ? _GEN8745 : _GEN8738;
wire  _GEN8747 = io_x[18] ? _GEN8746 : _GEN8735;
wire  _GEN8748 = io_x[33] ? _GEN8747 : _GEN8732;
wire  _GEN8749 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8750 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8751 = io_x[19] ? _GEN8750 : _GEN8749;
wire  _GEN8752 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8753 = io_x[27] ? _GEN8752 : _GEN7271;
wire  _GEN8754 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8755 = io_x[27] ? _GEN8754 : _GEN7278;
wire  _GEN8756 = io_x[19] ? _GEN8755 : _GEN8753;
wire  _GEN8757 = io_x[23] ? _GEN8756 : _GEN8751;
wire  _GEN8758 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8759 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8760 = io_x[27] ? _GEN8759 : _GEN8758;
wire  _GEN8761 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8762 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8763 = io_x[27] ? _GEN8762 : _GEN8761;
wire  _GEN8764 = io_x[19] ? _GEN8763 : _GEN8760;
wire  _GEN8765 = io_x[23] ? _GEN8764 : _GEN7305;
wire  _GEN8766 = io_x[18] ? _GEN8765 : _GEN8757;
wire  _GEN8767 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8768 = io_x[27] ? _GEN8767 : _GEN7278;
wire  _GEN8769 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8770 = io_x[19] ? _GEN8769 : _GEN8768;
wire  _GEN8771 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8772 = io_x[27] ? _GEN8771 : _GEN7271;
wire  _GEN8773 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8774 = io_x[27] ? _GEN8773 : _GEN7278;
wire  _GEN8775 = io_x[19] ? _GEN8774 : _GEN8772;
wire  _GEN8776 = io_x[23] ? _GEN8775 : _GEN8770;
wire  _GEN8777 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8778 = io_x[27] ? _GEN8777 : _GEN7271;
wire  _GEN8779 = io_x[19] ? _GEN8778 : _GEN7273;
wire  _GEN8780 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8781 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8782 = io_x[27] ? _GEN8781 : _GEN8780;
wire  _GEN8783 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8784 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8785 = io_x[27] ? _GEN8784 : _GEN8783;
wire  _GEN8786 = io_x[19] ? _GEN8785 : _GEN8782;
wire  _GEN8787 = io_x[23] ? _GEN8786 : _GEN8779;
wire  _GEN8788 = io_x[18] ? _GEN8787 : _GEN8776;
wire  _GEN8789 = io_x[33] ? _GEN8788 : _GEN8766;
wire  _GEN8790 = io_x[31] ? _GEN8789 : _GEN8748;
wire  _GEN8791 = io_x[28] ? _GEN8790 : _GEN8719;
wire  _GEN8792 = io_x[26] ? _GEN8791 : _GEN8658;
wire  _GEN8793 = io_x[20] ? _GEN8792 : _GEN8571;
wire  _GEN8794 = io_x[24] ? _GEN8793 : _GEN8468;
wire  _GEN8795 = io_x[78] ? _GEN8794 : _GEN8230;
wire  _GEN8796 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8797 = io_x[23] ? _GEN8796 : _GEN7305;
wire  _GEN8798 = io_x[18] ? _GEN7297 : _GEN8797;
wire  _GEN8799 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8800 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8801 = io_x[27] ? _GEN8800 : _GEN8799;
wire  _GEN8802 = io_x[19] ? _GEN8801 : _GEN7273;
wire  _GEN8803 = io_x[23] ? _GEN8802 : _GEN7267;
wire  _GEN8804 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8805 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8806 = io_x[27] ? _GEN8805 : _GEN8804;
wire  _GEN8807 = io_x[19] ? _GEN8806 : _GEN7273;
wire  _GEN8808 = io_x[23] ? _GEN8807 : _GEN7267;
wire  _GEN8809 = io_x[18] ? _GEN8808 : _GEN8803;
wire  _GEN8810 = io_x[33] ? _GEN8809 : _GEN8798;
wire  _GEN8811 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8812 = io_x[27] ? _GEN8811 : _GEN7278;
wire  _GEN8813 = io_x[19] ? _GEN8812 : _GEN7280;
wire  _GEN8814 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8815 = io_x[19] ? _GEN8814 : _GEN7280;
wire  _GEN8816 = io_x[23] ? _GEN8815 : _GEN8813;
wire  _GEN8817 = io_x[18] ? _GEN7297 : _GEN8816;
wire  _GEN8818 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN8819 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8820 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8821 = io_x[27] ? _GEN8820 : _GEN8819;
wire  _GEN8822 = io_x[19] ? _GEN8821 : _GEN7280;
wire  _GEN8823 = io_x[23] ? _GEN8822 : _GEN8818;
wire  _GEN8824 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8825 = io_x[27] ? _GEN8824 : _GEN7278;
wire  _GEN8826 = io_x[19] ? _GEN8825 : _GEN7280;
wire  _GEN8827 = io_x[23] ? _GEN8826 : _GEN7305;
wire  _GEN8828 = io_x[18] ? _GEN8827 : _GEN8823;
wire  _GEN8829 = io_x[33] ? _GEN8828 : _GEN8817;
wire  _GEN8830 = io_x[31] ? _GEN8829 : _GEN8810;
wire  _GEN8831 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN8832 = io_x[18] ? _GEN7297 : _GEN8831;
wire  _GEN8833 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8834 = io_x[19] ? _GEN8833 : _GEN7280;
wire  _GEN8835 = io_x[23] ? _GEN7305 : _GEN8834;
wire  _GEN8836 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8837 = io_x[27] ? _GEN8836 : _GEN7278;
wire  _GEN8838 = io_x[19] ? _GEN8837 : _GEN7273;
wire  _GEN8839 = io_x[23] ? _GEN7305 : _GEN8838;
wire  _GEN8840 = io_x[18] ? _GEN8839 : _GEN8835;
wire  _GEN8841 = io_x[33] ? _GEN8840 : _GEN8832;
wire  _GEN8842 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8843 = io_x[19] ? _GEN8842 : _GEN7280;
wire  _GEN8844 = io_x[23] ? _GEN7267 : _GEN8843;
wire  _GEN8845 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8846 = io_x[19] ? _GEN8845 : _GEN7280;
wire  _GEN8847 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8848 = io_x[27] ? _GEN8847 : _GEN7278;
wire  _GEN8849 = io_x[19] ? _GEN8848 : _GEN7273;
wire  _GEN8850 = io_x[23] ? _GEN8849 : _GEN8846;
wire  _GEN8851 = io_x[18] ? _GEN8850 : _GEN8844;
wire  _GEN8852 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8853 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8854 = io_x[27] ? _GEN8853 : _GEN8852;
wire  _GEN8855 = io_x[19] ? _GEN8854 : _GEN7273;
wire  _GEN8856 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8857 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8858 = io_x[27] ? _GEN8857 : _GEN8856;
wire  _GEN8859 = io_x[19] ? _GEN8858 : _GEN7280;
wire  _GEN8860 = io_x[23] ? _GEN8859 : _GEN8855;
wire  _GEN8861 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8862 = io_x[27] ? _GEN8861 : _GEN7271;
wire  _GEN8863 = io_x[19] ? _GEN8862 : _GEN7280;
wire  _GEN8864 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8865 = io_x[27] ? _GEN8864 : _GEN7278;
wire  _GEN8866 = io_x[19] ? _GEN8865 : _GEN7280;
wire  _GEN8867 = io_x[23] ? _GEN8866 : _GEN8863;
wire  _GEN8868 = io_x[18] ? _GEN8867 : _GEN8860;
wire  _GEN8869 = io_x[33] ? _GEN8868 : _GEN8851;
wire  _GEN8870 = io_x[31] ? _GEN8869 : _GEN8841;
wire  _GEN8871 = io_x[28] ? _GEN8870 : _GEN8830;
wire  _GEN8872 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8873 = io_x[27] ? _GEN8872 : _GEN7278;
wire  _GEN8874 = io_x[19] ? _GEN8873 : _GEN7280;
wire  _GEN8875 = io_x[23] ? _GEN8874 : _GEN7267;
wire  _GEN8876 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN8877 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN8878 = io_x[23] ? _GEN8877 : _GEN8876;
wire  _GEN8879 = io_x[18] ? _GEN8878 : _GEN8875;
wire  _GEN8880 = io_x[33] ? _GEN8879 : _GEN8346;
wire  _GEN8881 = io_x[18] ? _GEN7266 : _GEN7297;
wire  _GEN8882 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8883 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8884 = io_x[27] ? _GEN8883 : _GEN7271;
wire  _GEN8885 = io_x[19] ? _GEN8884 : _GEN8882;
wire  _GEN8886 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8887 = io_x[27] ? _GEN8886 : _GEN7278;
wire  _GEN8888 = io_x[19] ? _GEN8887 : _GEN7280;
wire  _GEN8889 = io_x[23] ? _GEN8888 : _GEN8885;
wire  _GEN8890 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8891 = io_x[27] ? _GEN8890 : _GEN7271;
wire  _GEN8892 = io_x[19] ? _GEN8891 : _GEN7280;
wire  _GEN8893 = io_x[23] ? _GEN8892 : _GEN7305;
wire  _GEN8894 = io_x[18] ? _GEN8893 : _GEN8889;
wire  _GEN8895 = io_x[33] ? _GEN8894 : _GEN8881;
wire  _GEN8896 = io_x[31] ? _GEN8895 : _GEN8880;
wire  _GEN8897 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8898 = io_x[27] ? _GEN7278 : _GEN8897;
wire  _GEN8899 = io_x[19] ? _GEN8898 : _GEN7273;
wire  _GEN8900 = io_x[23] ? _GEN7267 : _GEN8899;
wire  _GEN8901 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8902 = io_x[19] ? _GEN8901 : _GEN7280;
wire  _GEN8903 = io_x[23] ? _GEN8902 : _GEN7305;
wire  _GEN8904 = io_x[18] ? _GEN8903 : _GEN8900;
wire  _GEN8905 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN8906 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8907 = io_x[27] ? _GEN7278 : _GEN8906;
wire  _GEN8908 = io_x[19] ? _GEN8907 : _GEN7280;
wire  _GEN8909 = io_x[23] ? _GEN8908 : _GEN8905;
wire  _GEN8910 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8911 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8912 = io_x[27] ? _GEN8911 : _GEN8910;
wire  _GEN8913 = io_x[19] ? _GEN8912 : _GEN7273;
wire  _GEN8914 = io_x[23] ? _GEN8913 : _GEN7267;
wire  _GEN8915 = io_x[18] ? _GEN8914 : _GEN8909;
wire  _GEN8916 = io_x[33] ? _GEN8915 : _GEN8904;
wire  _GEN8917 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN8918 = io_x[18] ? _GEN7266 : _GEN8917;
wire  _GEN8919 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8920 = io_x[27] ? _GEN7271 : _GEN8919;
wire  _GEN8921 = io_x[19] ? _GEN8920 : _GEN7280;
wire  _GEN8922 = io_x[23] ? _GEN8921 : _GEN7267;
wire  _GEN8923 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN8924 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8925 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8926 = io_x[27] ? _GEN8925 : _GEN7271;
wire  _GEN8927 = io_x[19] ? _GEN8926 : _GEN8924;
wire  _GEN8928 = io_x[23] ? _GEN8927 : _GEN8923;
wire  _GEN8929 = io_x[18] ? _GEN8928 : _GEN8922;
wire  _GEN8930 = io_x[33] ? _GEN8929 : _GEN8918;
wire  _GEN8931 = io_x[31] ? _GEN8930 : _GEN8916;
wire  _GEN8932 = io_x[28] ? _GEN8931 : _GEN8896;
wire  _GEN8933 = io_x[26] ? _GEN8932 : _GEN8871;
wire  _GEN8934 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8935 = io_x[27] ? _GEN8934 : _GEN7278;
wire  _GEN8936 = io_x[19] ? _GEN8935 : _GEN7273;
wire  _GEN8937 = io_x[23] ? _GEN8936 : _GEN7305;
wire  _GEN8938 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN8939 = io_x[23] ? _GEN8938 : _GEN7267;
wire  _GEN8940 = io_x[18] ? _GEN8939 : _GEN8937;
wire  _GEN8941 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8942 = io_x[27] ? _GEN8941 : _GEN7278;
wire  _GEN8943 = io_x[19] ? _GEN8942 : _GEN7280;
wire  _GEN8944 = io_x[23] ? _GEN8943 : _GEN7305;
wire  _GEN8945 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8946 = io_x[27] ? _GEN8945 : _GEN7271;
wire  _GEN8947 = io_x[19] ? _GEN8946 : _GEN7273;
wire  _GEN8948 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8949 = io_x[27] ? _GEN7278 : _GEN8948;
wire  _GEN8950 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8951 = io_x[27] ? _GEN8950 : _GEN7278;
wire  _GEN8952 = io_x[19] ? _GEN8951 : _GEN8949;
wire  _GEN8953 = io_x[23] ? _GEN8952 : _GEN8947;
wire  _GEN8954 = io_x[18] ? _GEN8953 : _GEN8944;
wire  _GEN8955 = io_x[33] ? _GEN8954 : _GEN8940;
wire  _GEN8956 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8957 = io_x[27] ? _GEN8956 : _GEN7278;
wire  _GEN8958 = io_x[19] ? _GEN8957 : _GEN7273;
wire  _GEN8959 = io_x[23] ? _GEN8958 : _GEN7267;
wire  _GEN8960 = io_x[18] ? _GEN7266 : _GEN8959;
wire  _GEN8961 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN8962 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8963 = io_x[27] ? _GEN8962 : _GEN7278;
wire  _GEN8964 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8965 = io_x[27] ? _GEN8964 : _GEN7278;
wire  _GEN8966 = io_x[19] ? _GEN8965 : _GEN8963;
wire  _GEN8967 = io_x[23] ? _GEN8966 : _GEN8961;
wire  _GEN8968 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8969 = io_x[27] ? _GEN7278 : _GEN8968;
wire  _GEN8970 = io_x[19] ? _GEN8969 : _GEN7273;
wire  _GEN8971 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8972 = io_x[27] ? _GEN8971 : _GEN7278;
wire  _GEN8973 = io_x[19] ? _GEN8972 : _GEN7273;
wire  _GEN8974 = io_x[23] ? _GEN8973 : _GEN8970;
wire  _GEN8975 = io_x[18] ? _GEN8974 : _GEN8967;
wire  _GEN8976 = io_x[33] ? _GEN8975 : _GEN8960;
wire  _GEN8977 = io_x[31] ? _GEN8976 : _GEN8955;
wire  _GEN8978 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN8979 = io_x[18] ? _GEN8978 : _GEN7266;
wire  _GEN8980 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN8981 = io_x[19] ? _GEN8980 : _GEN7280;
wire  _GEN8982 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN8983 = io_x[23] ? _GEN8982 : _GEN8981;
wire  _GEN8984 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8985 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8986 = io_x[27] ? _GEN8985 : _GEN8984;
wire  _GEN8987 = io_x[19] ? _GEN8986 : _GEN7280;
wire  _GEN8988 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN8989 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8990 = io_x[27] ? _GEN8989 : _GEN8988;
wire  _GEN8991 = io_x[19] ? _GEN8990 : _GEN7280;
wire  _GEN8992 = io_x[23] ? _GEN8991 : _GEN8987;
wire  _GEN8993 = io_x[18] ? _GEN8992 : _GEN8983;
wire  _GEN8994 = io_x[33] ? _GEN8993 : _GEN8979;
wire  _GEN8995 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN8996 = io_x[19] ? _GEN7273 : _GEN8995;
wire  _GEN8997 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN8998 = io_x[27] ? _GEN8997 : _GEN7278;
wire  _GEN8999 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9000 = io_x[19] ? _GEN8999 : _GEN8998;
wire  _GEN9001 = io_x[23] ? _GEN9000 : _GEN8996;
wire  _GEN9002 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9003 = io_x[27] ? _GEN9002 : _GEN7278;
wire  _GEN9004 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9005 = io_x[27] ? _GEN7278 : _GEN9004;
wire  _GEN9006 = io_x[19] ? _GEN9005 : _GEN9003;
wire  _GEN9007 = io_x[23] ? _GEN9006 : _GEN7305;
wire  _GEN9008 = io_x[18] ? _GEN9007 : _GEN9001;
wire  _GEN9009 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9010 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9011 = io_x[27] ? _GEN7278 : _GEN9010;
wire  _GEN9012 = io_x[19] ? _GEN9011 : _GEN9009;
wire  _GEN9013 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9014 = io_x[27] ? _GEN9013 : _GEN7278;
wire  _GEN9015 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9016 = io_x[27] ? _GEN9015 : _GEN7278;
wire  _GEN9017 = io_x[19] ? _GEN9016 : _GEN9014;
wire  _GEN9018 = io_x[23] ? _GEN9017 : _GEN9012;
wire  _GEN9019 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9020 = io_x[19] ? _GEN9019 : _GEN7273;
wire  _GEN9021 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9022 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9023 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9024 = io_x[27] ? _GEN9023 : _GEN9022;
wire  _GEN9025 = io_x[19] ? _GEN9024 : _GEN9021;
wire  _GEN9026 = io_x[23] ? _GEN9025 : _GEN9020;
wire  _GEN9027 = io_x[18] ? _GEN9026 : _GEN9018;
wire  _GEN9028 = io_x[33] ? _GEN9027 : _GEN9008;
wire  _GEN9029 = io_x[31] ? _GEN9028 : _GEN8994;
wire  _GEN9030 = io_x[28] ? _GEN9029 : _GEN8977;
wire  _GEN9031 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9032 = io_x[27] ? _GEN9031 : _GEN7271;
wire  _GEN9033 = io_x[19] ? _GEN7280 : _GEN9032;
wire  _GEN9034 = io_x[23] ? _GEN9033 : _GEN7305;
wire  _GEN9035 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9036 = io_x[27] ? _GEN7271 : _GEN9035;
wire  _GEN9037 = io_x[19] ? _GEN9036 : _GEN7273;
wire  _GEN9038 = io_x[23] ? _GEN9037 : _GEN7267;
wire  _GEN9039 = io_x[18] ? _GEN9038 : _GEN9034;
wire  _GEN9040 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9041 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9042 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9043 = io_x[27] ? _GEN9042 : _GEN9041;
wire  _GEN9044 = io_x[19] ? _GEN9043 : _GEN9040;
wire  _GEN9045 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9046 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9047 = io_x[27] ? _GEN9046 : _GEN9045;
wire  _GEN9048 = io_x[19] ? _GEN7280 : _GEN9047;
wire  _GEN9049 = io_x[23] ? _GEN9048 : _GEN9044;
wire  _GEN9050 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9051 = io_x[19] ? _GEN9050 : _GEN7280;
wire  _GEN9052 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9053 = io_x[19] ? _GEN9052 : _GEN7273;
wire  _GEN9054 = io_x[23] ? _GEN9053 : _GEN9051;
wire  _GEN9055 = io_x[18] ? _GEN9054 : _GEN9049;
wire  _GEN9056 = io_x[33] ? _GEN9055 : _GEN9039;
wire  _GEN9057 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9058 = io_x[19] ? _GEN7280 : _GEN9057;
wire  _GEN9059 = io_x[23] ? _GEN7267 : _GEN9058;
wire  _GEN9060 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9061 = io_x[27] ? _GEN9060 : _GEN7278;
wire  _GEN9062 = io_x[19] ? _GEN7280 : _GEN9061;
wire  _GEN9063 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9064 = io_x[27] ? _GEN9063 : _GEN7278;
wire  _GEN9065 = io_x[19] ? _GEN9064 : _GEN7280;
wire  _GEN9066 = io_x[23] ? _GEN9065 : _GEN9062;
wire  _GEN9067 = io_x[18] ? _GEN9066 : _GEN9059;
wire  _GEN9068 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9069 = io_x[19] ? _GEN7280 : _GEN9068;
wire  _GEN9070 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9071 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9072 = io_x[27] ? _GEN9071 : _GEN9070;
wire  _GEN9073 = io_x[19] ? _GEN9072 : _GEN7280;
wire  _GEN9074 = io_x[23] ? _GEN9073 : _GEN9069;
wire  _GEN9075 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9076 = io_x[27] ? _GEN9075 : _GEN7278;
wire  _GEN9077 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9078 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9079 = io_x[27] ? _GEN9078 : _GEN9077;
wire  _GEN9080 = io_x[19] ? _GEN9079 : _GEN9076;
wire  _GEN9081 = io_x[23] ? _GEN9080 : _GEN7267;
wire  _GEN9082 = io_x[18] ? _GEN9081 : _GEN9074;
wire  _GEN9083 = io_x[33] ? _GEN9082 : _GEN9067;
wire  _GEN9084 = io_x[31] ? _GEN9083 : _GEN9056;
wire  _GEN9085 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9086 = io_x[27] ? _GEN7278 : _GEN9085;
wire  _GEN9087 = io_x[19] ? _GEN9086 : _GEN7273;
wire  _GEN9088 = io_x[23] ? _GEN9087 : _GEN7267;
wire  _GEN9089 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9090 = io_x[27] ? _GEN7278 : _GEN9089;
wire  _GEN9091 = io_x[19] ? _GEN7280 : _GEN9090;
wire  _GEN9092 = io_x[23] ? _GEN7305 : _GEN9091;
wire  _GEN9093 = io_x[18] ? _GEN9092 : _GEN9088;
wire  _GEN9094 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9095 = io_x[19] ? _GEN9094 : _GEN7280;
wire  _GEN9096 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9097 = io_x[27] ? _GEN9096 : _GEN7271;
wire  _GEN9098 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9099 = io_x[27] ? _GEN7278 : _GEN9098;
wire  _GEN9100 = io_x[19] ? _GEN9099 : _GEN9097;
wire  _GEN9101 = io_x[23] ? _GEN9100 : _GEN9095;
wire  _GEN9102 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9103 = io_x[27] ? _GEN7278 : _GEN9102;
wire  _GEN9104 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9105 = io_x[27] ? _GEN7278 : _GEN9104;
wire  _GEN9106 = io_x[19] ? _GEN9105 : _GEN9103;
wire  _GEN9107 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9108 = io_x[27] ? _GEN9107 : _GEN7271;
wire  _GEN9109 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9110 = io_x[27] ? _GEN7278 : _GEN9109;
wire  _GEN9111 = io_x[19] ? _GEN9110 : _GEN9108;
wire  _GEN9112 = io_x[23] ? _GEN9111 : _GEN9106;
wire  _GEN9113 = io_x[18] ? _GEN9112 : _GEN9101;
wire  _GEN9114 = io_x[33] ? _GEN9113 : _GEN9093;
wire  _GEN9115 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9116 = io_x[27] ? _GEN9115 : _GEN7278;
wire  _GEN9117 = io_x[19] ? _GEN9116 : _GEN7273;
wire  _GEN9118 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9119 = io_x[23] ? _GEN9118 : _GEN9117;
wire  _GEN9120 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9121 = io_x[27] ? _GEN9120 : _GEN7278;
wire  _GEN9122 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9123 = io_x[27] ? _GEN9122 : _GEN7278;
wire  _GEN9124 = io_x[19] ? _GEN9123 : _GEN9121;
wire  _GEN9125 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9126 = io_x[27] ? _GEN9125 : _GEN7278;
wire  _GEN9127 = io_x[19] ? _GEN9126 : _GEN7280;
wire  _GEN9128 = io_x[23] ? _GEN9127 : _GEN9124;
wire  _GEN9129 = io_x[18] ? _GEN9128 : _GEN9119;
wire  _GEN9130 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9131 = io_x[27] ? _GEN9130 : _GEN7278;
wire  _GEN9132 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9133 = io_x[27] ? _GEN7271 : _GEN9132;
wire  _GEN9134 = io_x[19] ? _GEN9133 : _GEN9131;
wire  _GEN9135 = io_x[23] ? _GEN9134 : _GEN7305;
wire  _GEN9136 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9137 = io_x[27] ? _GEN9136 : _GEN7278;
wire  _GEN9138 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9139 = io_x[27] ? _GEN9138 : _GEN7271;
wire  _GEN9140 = io_x[19] ? _GEN9139 : _GEN9137;
wire  _GEN9141 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9142 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9143 = io_x[27] ? _GEN9142 : _GEN9141;
wire  _GEN9144 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9145 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9146 = io_x[27] ? _GEN9145 : _GEN9144;
wire  _GEN9147 = io_x[19] ? _GEN9146 : _GEN9143;
wire  _GEN9148 = io_x[23] ? _GEN9147 : _GEN9140;
wire  _GEN9149 = io_x[18] ? _GEN9148 : _GEN9135;
wire  _GEN9150 = io_x[33] ? _GEN9149 : _GEN9129;
wire  _GEN9151 = io_x[31] ? _GEN9150 : _GEN9114;
wire  _GEN9152 = io_x[28] ? _GEN9151 : _GEN9084;
wire  _GEN9153 = io_x[26] ? _GEN9152 : _GEN9030;
wire  _GEN9154 = io_x[20] ? _GEN9153 : _GEN8933;
wire  _GEN9155 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN9156 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9157 = io_x[27] ? _GEN9156 : _GEN7278;
wire  _GEN9158 = io_x[19] ? _GEN9157 : _GEN7280;
wire  _GEN9159 = io_x[23] ? _GEN9158 : _GEN7305;
wire  _GEN9160 = io_x[18] ? _GEN9159 : _GEN9155;
wire  _GEN9161 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9162 = io_x[27] ? _GEN9161 : _GEN7278;
wire  _GEN9163 = io_x[19] ? _GEN9162 : _GEN7280;
wire  _GEN9164 = io_x[23] ? _GEN9163 : _GEN7267;
wire  _GEN9165 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9166 = io_x[19] ? _GEN9165 : _GEN7273;
wire  _GEN9167 = io_x[23] ? _GEN7267 : _GEN9166;
wire  _GEN9168 = io_x[18] ? _GEN9167 : _GEN9164;
wire  _GEN9169 = io_x[33] ? _GEN9168 : _GEN9160;
wire  _GEN9170 = io_x[23] ? _GEN7267 : _GEN7305;
wire  _GEN9171 = io_x[23] ? _GEN7267 : _GEN7305;
wire  _GEN9172 = io_x[18] ? _GEN9171 : _GEN9170;
wire  _GEN9173 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9174 = io_x[27] ? _GEN9173 : _GEN7278;
wire  _GEN9175 = io_x[19] ? _GEN9174 : _GEN7273;
wire  _GEN9176 = io_x[23] ? _GEN9175 : _GEN7305;
wire  _GEN9177 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9178 = io_x[27] ? _GEN9177 : _GEN7278;
wire  _GEN9179 = io_x[19] ? _GEN7280 : _GEN9178;
wire  _GEN9180 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9181 = io_x[27] ? _GEN9180 : _GEN7278;
wire  _GEN9182 = io_x[19] ? _GEN9181 : _GEN7273;
wire  _GEN9183 = io_x[23] ? _GEN9182 : _GEN9179;
wire  _GEN9184 = io_x[18] ? _GEN9183 : _GEN9176;
wire  _GEN9185 = io_x[33] ? _GEN9184 : _GEN9172;
wire  _GEN9186 = io_x[31] ? _GEN9185 : _GEN9169;
wire  _GEN9187 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9188 = io_x[19] ? _GEN7280 : _GEN9187;
wire  _GEN9189 = io_x[23] ? _GEN7305 : _GEN9188;
wire  _GEN9190 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9191 = io_x[19] ? _GEN9190 : _GEN7280;
wire  _GEN9192 = io_x[23] ? _GEN9191 : _GEN7267;
wire  _GEN9193 = io_x[18] ? _GEN9192 : _GEN9189;
wire  _GEN9194 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9195 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9196 = io_x[27] ? _GEN9195 : _GEN7278;
wire  _GEN9197 = io_x[19] ? _GEN9196 : _GEN9194;
wire  _GEN9198 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9199 = io_x[27] ? _GEN9198 : _GEN7278;
wire  _GEN9200 = io_x[19] ? _GEN9199 : _GEN7280;
wire  _GEN9201 = io_x[23] ? _GEN9200 : _GEN9197;
wire  _GEN9202 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9203 = io_x[27] ? _GEN9202 : _GEN7278;
wire  _GEN9204 = io_x[19] ? _GEN9203 : _GEN7273;
wire  _GEN9205 = io_x[23] ? _GEN9204 : _GEN7267;
wire  _GEN9206 = io_x[18] ? _GEN9205 : _GEN9201;
wire  _GEN9207 = io_x[33] ? _GEN9206 : _GEN9193;
wire  _GEN9208 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN9209 = io_x[18] ? _GEN9208 : _GEN7266;
wire  _GEN9210 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9211 = io_x[27] ? _GEN7278 : _GEN9210;
wire  _GEN9212 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9213 = io_x[27] ? _GEN9212 : _GEN7278;
wire  _GEN9214 = io_x[19] ? _GEN9213 : _GEN9211;
wire  _GEN9215 = io_x[23] ? _GEN9214 : _GEN7267;
wire  _GEN9216 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9217 = io_x[27] ? _GEN7271 : _GEN9216;
wire  _GEN9218 = io_x[19] ? _GEN7280 : _GEN9217;
wire  _GEN9219 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9220 = io_x[27] ? _GEN7271 : _GEN9219;
wire  _GEN9221 = io_x[19] ? _GEN9220 : _GEN7273;
wire  _GEN9222 = io_x[23] ? _GEN9221 : _GEN9218;
wire  _GEN9223 = io_x[18] ? _GEN9222 : _GEN9215;
wire  _GEN9224 = io_x[33] ? _GEN9223 : _GEN9209;
wire  _GEN9225 = io_x[31] ? _GEN9224 : _GEN9207;
wire  _GEN9226 = io_x[28] ? _GEN9225 : _GEN9186;
wire  _GEN9227 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9228 = io_x[19] ? _GEN7280 : _GEN9227;
wire  _GEN9229 = io_x[23] ? _GEN7267 : _GEN9228;
wire  _GEN9230 = io_x[18] ? _GEN9229 : _GEN7297;
wire  _GEN9231 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9232 = io_x[27] ? _GEN9231 : _GEN7278;
wire  _GEN9233 = io_x[19] ? _GEN9232 : _GEN7280;
wire  _GEN9234 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9235 = io_x[27] ? _GEN7278 : _GEN9234;
wire  _GEN9236 = io_x[19] ? _GEN9235 : _GEN7280;
wire  _GEN9237 = io_x[23] ? _GEN9236 : _GEN9233;
wire  _GEN9238 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9239 = io_x[27] ? _GEN7278 : _GEN9238;
wire  _GEN9240 = io_x[19] ? _GEN9239 : _GEN7273;
wire  _GEN9241 = io_x[23] ? _GEN7267 : _GEN9240;
wire  _GEN9242 = io_x[18] ? _GEN9241 : _GEN9237;
wire  _GEN9243 = io_x[33] ? _GEN9242 : _GEN9230;
wire  _GEN9244 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9245 = io_x[27] ? _GEN9244 : _GEN7278;
wire  _GEN9246 = io_x[19] ? _GEN9245 : _GEN7273;
wire  _GEN9247 = io_x[23] ? _GEN7305 : _GEN9246;
wire  _GEN9248 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9249 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9250 = io_x[27] ? _GEN9249 : _GEN9248;
wire  _GEN9251 = io_x[19] ? _GEN9250 : _GEN7280;
wire  _GEN9252 = io_x[23] ? _GEN9251 : _GEN7267;
wire  _GEN9253 = io_x[18] ? _GEN9252 : _GEN9247;
wire  _GEN9254 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9255 = io_x[27] ? _GEN9254 : _GEN7278;
wire  _GEN9256 = io_x[19] ? _GEN9255 : _GEN7280;
wire  _GEN9257 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9258 = io_x[27] ? _GEN7271 : _GEN9257;
wire  _GEN9259 = io_x[19] ? _GEN9258 : _GEN7273;
wire  _GEN9260 = io_x[23] ? _GEN9259 : _GEN9256;
wire  _GEN9261 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9262 = io_x[27] ? _GEN7271 : _GEN9261;
wire  _GEN9263 = io_x[19] ? _GEN7273 : _GEN9262;
wire  _GEN9264 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9265 = io_x[27] ? _GEN9264 : _GEN7271;
wire  _GEN9266 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9267 = io_x[27] ? _GEN9266 : _GEN7278;
wire  _GEN9268 = io_x[19] ? _GEN9267 : _GEN9265;
wire  _GEN9269 = io_x[23] ? _GEN9268 : _GEN9263;
wire  _GEN9270 = io_x[18] ? _GEN9269 : _GEN9260;
wire  _GEN9271 = io_x[33] ? _GEN9270 : _GEN9253;
wire  _GEN9272 = io_x[31] ? _GEN9271 : _GEN9243;
wire  _GEN9273 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9274 = io_x[27] ? _GEN9273 : _GEN7278;
wire  _GEN9275 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9276 = io_x[27] ? _GEN7278 : _GEN9275;
wire  _GEN9277 = io_x[19] ? _GEN9276 : _GEN9274;
wire  _GEN9278 = io_x[23] ? _GEN9277 : _GEN7305;
wire  _GEN9279 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9280 = io_x[19] ? _GEN9279 : _GEN7280;
wire  _GEN9281 = io_x[23] ? _GEN7267 : _GEN9280;
wire  _GEN9282 = io_x[18] ? _GEN9281 : _GEN9278;
wire  _GEN9283 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9284 = io_x[27] ? _GEN7278 : _GEN9283;
wire  _GEN9285 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9286 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9287 = io_x[27] ? _GEN9286 : _GEN9285;
wire  _GEN9288 = io_x[19] ? _GEN9287 : _GEN9284;
wire  _GEN9289 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9290 = io_x[27] ? _GEN9289 : _GEN7278;
wire  _GEN9291 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9292 = io_x[27] ? _GEN7278 : _GEN9291;
wire  _GEN9293 = io_x[19] ? _GEN9292 : _GEN9290;
wire  _GEN9294 = io_x[23] ? _GEN9293 : _GEN9288;
wire  _GEN9295 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9296 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9297 = io_x[19] ? _GEN9296 : _GEN9295;
wire  _GEN9298 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9299 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9300 = io_x[27] ? _GEN9299 : _GEN7271;
wire  _GEN9301 = io_x[19] ? _GEN9300 : _GEN9298;
wire  _GEN9302 = io_x[23] ? _GEN9301 : _GEN9297;
wire  _GEN9303 = io_x[18] ? _GEN9302 : _GEN9294;
wire  _GEN9304 = io_x[33] ? _GEN9303 : _GEN9282;
wire  _GEN9305 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9306 = io_x[23] ? _GEN9305 : _GEN7267;
wire  _GEN9307 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9308 = io_x[27] ? _GEN9307 : _GEN7271;
wire  _GEN9309 = io_x[19] ? _GEN9308 : _GEN7280;
wire  _GEN9310 = io_x[23] ? _GEN9309 : _GEN7267;
wire  _GEN9311 = io_x[18] ? _GEN9310 : _GEN9306;
wire  _GEN9312 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9313 = io_x[27] ? _GEN7278 : _GEN9312;
wire  _GEN9314 = io_x[19] ? _GEN9313 : _GEN7273;
wire  _GEN9315 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9316 = io_x[27] ? _GEN9315 : _GEN7278;
wire  _GEN9317 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9318 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9319 = io_x[27] ? _GEN9318 : _GEN9317;
wire  _GEN9320 = io_x[19] ? _GEN9319 : _GEN9316;
wire  _GEN9321 = io_x[23] ? _GEN9320 : _GEN9314;
wire  _GEN9322 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9323 = io_x[27] ? _GEN7271 : _GEN9322;
wire  _GEN9324 = io_x[19] ? _GEN7280 : _GEN9323;
wire  _GEN9325 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9326 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9327 = io_x[27] ? _GEN9326 : _GEN9325;
wire  _GEN9328 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9329 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9330 = io_x[27] ? _GEN9329 : _GEN9328;
wire  _GEN9331 = io_x[19] ? _GEN9330 : _GEN9327;
wire  _GEN9332 = io_x[23] ? _GEN9331 : _GEN9324;
wire  _GEN9333 = io_x[18] ? _GEN9332 : _GEN9321;
wire  _GEN9334 = io_x[33] ? _GEN9333 : _GEN9311;
wire  _GEN9335 = io_x[31] ? _GEN9334 : _GEN9304;
wire  _GEN9336 = io_x[28] ? _GEN9335 : _GEN9272;
wire  _GEN9337 = io_x[26] ? _GEN9336 : _GEN9226;
wire  _GEN9338 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9339 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9340 = io_x[27] ? _GEN9339 : _GEN7278;
wire  _GEN9341 = io_x[19] ? _GEN9340 : _GEN9338;
wire  _GEN9342 = io_x[23] ? _GEN7267 : _GEN9341;
wire  _GEN9343 = io_x[18] ? _GEN9342 : _GEN7266;
wire  _GEN9344 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9345 = io_x[27] ? _GEN9344 : _GEN7271;
wire  _GEN9346 = io_x[19] ? _GEN9345 : _GEN7273;
wire  _GEN9347 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9348 = io_x[27] ? _GEN9347 : _GEN7271;
wire  _GEN9349 = io_x[19] ? _GEN9348 : _GEN7273;
wire  _GEN9350 = io_x[23] ? _GEN9349 : _GEN9346;
wire  _GEN9351 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9352 = io_x[27] ? _GEN9351 : _GEN7278;
wire  _GEN9353 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9354 = io_x[27] ? _GEN9353 : _GEN7271;
wire  _GEN9355 = io_x[19] ? _GEN9354 : _GEN9352;
wire  _GEN9356 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9357 = io_x[27] ? _GEN9356 : _GEN7278;
wire  _GEN9358 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9359 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9360 = io_x[27] ? _GEN9359 : _GEN9358;
wire  _GEN9361 = io_x[19] ? _GEN9360 : _GEN9357;
wire  _GEN9362 = io_x[23] ? _GEN9361 : _GEN9355;
wire  _GEN9363 = io_x[18] ? _GEN9362 : _GEN9350;
wire  _GEN9364 = io_x[33] ? _GEN9363 : _GEN9343;
wire  _GEN9365 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9366 = io_x[19] ? _GEN7280 : _GEN9365;
wire  _GEN9367 = io_x[23] ? _GEN9366 : _GEN7267;
wire  _GEN9368 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9369 = io_x[19] ? _GEN7273 : _GEN9368;
wire  _GEN9370 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9371 = io_x[27] ? _GEN9370 : _GEN7278;
wire  _GEN9372 = io_x[19] ? _GEN9371 : _GEN7273;
wire  _GEN9373 = io_x[23] ? _GEN9372 : _GEN9369;
wire  _GEN9374 = io_x[18] ? _GEN9373 : _GEN9367;
wire  _GEN9375 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9376 = io_x[27] ? _GEN9375 : _GEN7278;
wire  _GEN9377 = io_x[19] ? _GEN9376 : _GEN7280;
wire  _GEN9378 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9379 = io_x[27] ? _GEN9378 : _GEN7271;
wire  _GEN9380 = io_x[19] ? _GEN9379 : _GEN7280;
wire  _GEN9381 = io_x[23] ? _GEN9380 : _GEN9377;
wire  _GEN9382 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9383 = io_x[27] ? _GEN9382 : _GEN7278;
wire  _GEN9384 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9385 = io_x[27] ? _GEN9384 : _GEN7278;
wire  _GEN9386 = io_x[19] ? _GEN9385 : _GEN9383;
wire  _GEN9387 = io_x[23] ? _GEN7305 : _GEN9386;
wire  _GEN9388 = io_x[18] ? _GEN9387 : _GEN9381;
wire  _GEN9389 = io_x[33] ? _GEN9388 : _GEN9374;
wire  _GEN9390 = io_x[31] ? _GEN9389 : _GEN9364;
wire  _GEN9391 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9392 = io_x[19] ? _GEN9391 : _GEN7273;
wire  _GEN9393 = io_x[23] ? _GEN9392 : _GEN7267;
wire  _GEN9394 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9395 = io_x[27] ? _GEN9394 : _GEN7278;
wire  _GEN9396 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9397 = io_x[27] ? _GEN9396 : _GEN7271;
wire  _GEN9398 = io_x[19] ? _GEN9397 : _GEN9395;
wire  _GEN9399 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9400 = io_x[27] ? _GEN9399 : _GEN7278;
wire  _GEN9401 = io_x[19] ? _GEN9400 : _GEN7280;
wire  _GEN9402 = io_x[23] ? _GEN9401 : _GEN9398;
wire  _GEN9403 = io_x[18] ? _GEN9402 : _GEN9393;
wire  _GEN9404 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9405 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9406 = io_x[27] ? _GEN9405 : _GEN9404;
wire  _GEN9407 = io_x[19] ? _GEN9406 : _GEN7273;
wire  _GEN9408 = io_x[23] ? _GEN9407 : _GEN7267;
wire  _GEN9409 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9410 = io_x[27] ? _GEN9409 : _GEN7278;
wire  _GEN9411 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9412 = io_x[27] ? _GEN9411 : _GEN7278;
wire  _GEN9413 = io_x[19] ? _GEN9412 : _GEN9410;
wire  _GEN9414 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9415 = io_x[27] ? _GEN7278 : _GEN9414;
wire  _GEN9416 = io_x[19] ? _GEN9415 : _GEN7273;
wire  _GEN9417 = io_x[23] ? _GEN9416 : _GEN9413;
wire  _GEN9418 = io_x[18] ? _GEN9417 : _GEN9408;
wire  _GEN9419 = io_x[33] ? _GEN9418 : _GEN9403;
wire  _GEN9420 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9421 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9422 = io_x[19] ? _GEN9421 : _GEN9420;
wire  _GEN9423 = io_x[23] ? _GEN9422 : _GEN7267;
wire  _GEN9424 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9425 = io_x[27] ? _GEN7271 : _GEN9424;
wire  _GEN9426 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9427 = io_x[27] ? _GEN9426 : _GEN7278;
wire  _GEN9428 = io_x[19] ? _GEN9427 : _GEN9425;
wire  _GEN9429 = io_x[23] ? _GEN9428 : _GEN7305;
wire  _GEN9430 = io_x[18] ? _GEN9429 : _GEN9423;
wire  _GEN9431 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9432 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9433 = io_x[27] ? _GEN9432 : _GEN9431;
wire  _GEN9434 = io_x[19] ? _GEN9433 : _GEN7273;
wire  _GEN9435 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9436 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9437 = io_x[27] ? _GEN9436 : _GEN9435;
wire  _GEN9438 = io_x[19] ? _GEN9437 : _GEN7280;
wire  _GEN9439 = io_x[23] ? _GEN9438 : _GEN9434;
wire  _GEN9440 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9441 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9442 = io_x[27] ? _GEN9441 : _GEN9440;
wire  _GEN9443 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9444 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9445 = io_x[27] ? _GEN9444 : _GEN9443;
wire  _GEN9446 = io_x[19] ? _GEN9445 : _GEN9442;
wire  _GEN9447 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9448 = io_x[27] ? _GEN9447 : _GEN7278;
wire  _GEN9449 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9450 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9451 = io_x[27] ? _GEN9450 : _GEN9449;
wire  _GEN9452 = io_x[19] ? _GEN9451 : _GEN9448;
wire  _GEN9453 = io_x[23] ? _GEN9452 : _GEN9446;
wire  _GEN9454 = io_x[18] ? _GEN9453 : _GEN9439;
wire  _GEN9455 = io_x[33] ? _GEN9454 : _GEN9430;
wire  _GEN9456 = io_x[31] ? _GEN9455 : _GEN9419;
wire  _GEN9457 = io_x[28] ? _GEN9456 : _GEN9390;
wire  _GEN9458 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9459 = io_x[19] ? _GEN9458 : _GEN7280;
wire  _GEN9460 = io_x[23] ? _GEN9459 : _GEN7305;
wire  _GEN9461 = io_x[18] ? _GEN9460 : _GEN7297;
wire  _GEN9462 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9463 = io_x[19] ? _GEN9462 : _GEN7280;
wire  _GEN9464 = io_x[23] ? _GEN9463 : _GEN7267;
wire  _GEN9465 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9466 = io_x[27] ? _GEN9465 : _GEN7271;
wire  _GEN9467 = io_x[19] ? _GEN9466 : _GEN7280;
wire  _GEN9468 = io_x[23] ? _GEN9467 : _GEN7305;
wire  _GEN9469 = io_x[18] ? _GEN9468 : _GEN9464;
wire  _GEN9470 = io_x[33] ? _GEN9469 : _GEN9461;
wire  _GEN9471 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9472 = io_x[27] ? _GEN9471 : _GEN7278;
wire  _GEN9473 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9474 = io_x[19] ? _GEN9473 : _GEN9472;
wire  _GEN9475 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9476 = io_x[27] ? _GEN9475 : _GEN7278;
wire  _GEN9477 = io_x[19] ? _GEN9476 : _GEN7280;
wire  _GEN9478 = io_x[23] ? _GEN9477 : _GEN9474;
wire  _GEN9479 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9480 = io_x[27] ? _GEN9479 : _GEN7278;
wire  _GEN9481 = io_x[19] ? _GEN9480 : _GEN7280;
wire  _GEN9482 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9483 = io_x[27] ? _GEN9482 : _GEN7278;
wire  _GEN9484 = io_x[19] ? _GEN9483 : _GEN7273;
wire  _GEN9485 = io_x[23] ? _GEN9484 : _GEN9481;
wire  _GEN9486 = io_x[18] ? _GEN9485 : _GEN9478;
wire  _GEN9487 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9488 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9489 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9490 = io_x[27] ? _GEN9489 : _GEN9488;
wire  _GEN9491 = io_x[19] ? _GEN9490 : _GEN9487;
wire  _GEN9492 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9493 = io_x[27] ? _GEN7278 : _GEN9492;
wire  _GEN9494 = io_x[19] ? _GEN7273 : _GEN9493;
wire  _GEN9495 = io_x[23] ? _GEN9494 : _GEN9491;
wire  _GEN9496 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9497 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9498 = io_x[27] ? _GEN9497 : _GEN9496;
wire  _GEN9499 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9500 = io_x[27] ? _GEN9499 : _GEN7278;
wire  _GEN9501 = io_x[19] ? _GEN9500 : _GEN9498;
wire  _GEN9502 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9503 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9504 = io_x[27] ? _GEN9503 : _GEN9502;
wire  _GEN9505 = io_x[19] ? _GEN9504 : _GEN7280;
wire  _GEN9506 = io_x[23] ? _GEN9505 : _GEN9501;
wire  _GEN9507 = io_x[18] ? _GEN9506 : _GEN9495;
wire  _GEN9508 = io_x[33] ? _GEN9507 : _GEN9486;
wire  _GEN9509 = io_x[31] ? _GEN9508 : _GEN9470;
wire  _GEN9510 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9511 = io_x[19] ? _GEN9510 : _GEN7273;
wire  _GEN9512 = io_x[23] ? _GEN7267 : _GEN9511;
wire  _GEN9513 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9514 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9515 = io_x[27] ? _GEN9514 : _GEN9513;
wire  _GEN9516 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9517 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9518 = io_x[27] ? _GEN9517 : _GEN9516;
wire  _GEN9519 = io_x[19] ? _GEN9518 : _GEN9515;
wire  _GEN9520 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9521 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9522 = io_x[27] ? _GEN9521 : _GEN7278;
wire  _GEN9523 = io_x[19] ? _GEN9522 : _GEN9520;
wire  _GEN9524 = io_x[23] ? _GEN9523 : _GEN9519;
wire  _GEN9525 = io_x[18] ? _GEN9524 : _GEN9512;
wire  _GEN9526 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9527 = io_x[27] ? _GEN7278 : _GEN9526;
wire  _GEN9528 = io_x[19] ? _GEN9527 : _GEN7273;
wire  _GEN9529 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9530 = io_x[27] ? _GEN7271 : _GEN9529;
wire  _GEN9531 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9532 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9533 = io_x[27] ? _GEN9532 : _GEN9531;
wire  _GEN9534 = io_x[19] ? _GEN9533 : _GEN9530;
wire  _GEN9535 = io_x[23] ? _GEN9534 : _GEN9528;
wire  _GEN9536 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9537 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9538 = io_x[27] ? _GEN9537 : _GEN9536;
wire  _GEN9539 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9540 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9541 = io_x[27] ? _GEN9540 : _GEN9539;
wire  _GEN9542 = io_x[19] ? _GEN9541 : _GEN9538;
wire  _GEN9543 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9544 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9545 = io_x[27] ? _GEN9544 : _GEN9543;
wire  _GEN9546 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9547 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9548 = io_x[27] ? _GEN9547 : _GEN9546;
wire  _GEN9549 = io_x[19] ? _GEN9548 : _GEN9545;
wire  _GEN9550 = io_x[23] ? _GEN9549 : _GEN9542;
wire  _GEN9551 = io_x[18] ? _GEN9550 : _GEN9535;
wire  _GEN9552 = io_x[33] ? _GEN9551 : _GEN9525;
wire  _GEN9553 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9554 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9555 = io_x[27] ? _GEN9554 : _GEN7278;
wire  _GEN9556 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9557 = io_x[27] ? _GEN9556 : _GEN7271;
wire  _GEN9558 = io_x[19] ? _GEN9557 : _GEN9555;
wire  _GEN9559 = io_x[23] ? _GEN9558 : _GEN9553;
wire  _GEN9560 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9561 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9562 = io_x[27] ? _GEN9561 : _GEN7278;
wire  _GEN9563 = io_x[19] ? _GEN9562 : _GEN9560;
wire  _GEN9564 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9565 = io_x[27] ? _GEN9564 : _GEN7278;
wire  _GEN9566 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9567 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9568 = io_x[27] ? _GEN9567 : _GEN9566;
wire  _GEN9569 = io_x[19] ? _GEN9568 : _GEN9565;
wire  _GEN9570 = io_x[23] ? _GEN9569 : _GEN9563;
wire  _GEN9571 = io_x[18] ? _GEN9570 : _GEN9559;
wire  _GEN9572 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9573 = io_x[27] ? _GEN9572 : _GEN7278;
wire  _GEN9574 = io_x[19] ? _GEN9573 : _GEN7280;
wire  _GEN9575 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9576 = io_x[27] ? _GEN9575 : _GEN7271;
wire  _GEN9577 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9578 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9579 = io_x[27] ? _GEN9578 : _GEN9577;
wire  _GEN9580 = io_x[19] ? _GEN9579 : _GEN9576;
wire  _GEN9581 = io_x[23] ? _GEN9580 : _GEN9574;
wire  _GEN9582 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9583 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9584 = io_x[27] ? _GEN9583 : _GEN9582;
wire  _GEN9585 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9586 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9587 = io_x[27] ? _GEN9586 : _GEN9585;
wire  _GEN9588 = io_x[19] ? _GEN9587 : _GEN9584;
wire  _GEN9589 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9590 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9591 = io_x[27] ? _GEN9590 : _GEN9589;
wire  _GEN9592 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9593 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9594 = io_x[27] ? _GEN9593 : _GEN9592;
wire  _GEN9595 = io_x[19] ? _GEN9594 : _GEN9591;
wire  _GEN9596 = io_x[23] ? _GEN9595 : _GEN9588;
wire  _GEN9597 = io_x[18] ? _GEN9596 : _GEN9581;
wire  _GEN9598 = io_x[33] ? _GEN9597 : _GEN9571;
wire  _GEN9599 = io_x[31] ? _GEN9598 : _GEN9552;
wire  _GEN9600 = io_x[28] ? _GEN9599 : _GEN9509;
wire  _GEN9601 = io_x[26] ? _GEN9600 : _GEN9457;
wire  _GEN9602 = io_x[20] ? _GEN9601 : _GEN9337;
wire  _GEN9603 = io_x[24] ? _GEN9602 : _GEN9154;
wire  _GEN9604 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN9605 = io_x[18] ? _GEN7297 : _GEN9604;
wire  _GEN9606 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9607 = io_x[27] ? _GEN9606 : _GEN7278;
wire  _GEN9608 = io_x[19] ? _GEN9607 : _GEN7273;
wire  _GEN9609 = io_x[23] ? _GEN9608 : _GEN7267;
wire  _GEN9610 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9611 = io_x[19] ? _GEN7273 : _GEN9610;
wire  _GEN9612 = io_x[23] ? _GEN9611 : _GEN7267;
wire  _GEN9613 = io_x[18] ? _GEN9612 : _GEN9609;
wire  _GEN9614 = io_x[33] ? _GEN9613 : _GEN9605;
wire  _GEN9615 = io_x[23] ? _GEN7267 : _GEN7305;
wire  _GEN9616 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9617 = io_x[27] ? _GEN9616 : _GEN7278;
wire  _GEN9618 = io_x[19] ? _GEN9617 : _GEN7280;
wire  _GEN9619 = io_x[23] ? _GEN9618 : _GEN7267;
wire  _GEN9620 = io_x[18] ? _GEN9619 : _GEN9615;
wire  _GEN9621 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9622 = io_x[27] ? _GEN9621 : _GEN7278;
wire  _GEN9623 = io_x[19] ? _GEN9622 : _GEN7280;
wire  _GEN9624 = io_x[23] ? _GEN9623 : _GEN7267;
wire  _GEN9625 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9626 = io_x[27] ? _GEN9625 : _GEN7278;
wire  _GEN9627 = io_x[19] ? _GEN9626 : _GEN7280;
wire  _GEN9628 = io_x[23] ? _GEN9627 : _GEN7267;
wire  _GEN9629 = io_x[18] ? _GEN9628 : _GEN9624;
wire  _GEN9630 = io_x[33] ? _GEN9629 : _GEN9620;
wire  _GEN9631 = io_x[31] ? _GEN9630 : _GEN9614;
wire  _GEN9632 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9633 = io_x[27] ? _GEN7278 : _GEN9632;
wire  _GEN9634 = io_x[19] ? _GEN9633 : _GEN7280;
wire  _GEN9635 = io_x[23] ? _GEN7267 : _GEN9634;
wire  _GEN9636 = io_x[18] ? _GEN7297 : _GEN9635;
wire  _GEN9637 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN9638 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9639 = io_x[27] ? _GEN9638 : _GEN7278;
wire  _GEN9640 = io_x[19] ? _GEN9639 : _GEN7273;
wire  _GEN9641 = io_x[23] ? _GEN9640 : _GEN9637;
wire  _GEN9642 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9643 = io_x[27] ? _GEN9642 : _GEN7278;
wire  _GEN9644 = io_x[19] ? _GEN9643 : _GEN7273;
wire  _GEN9645 = io_x[23] ? _GEN9644 : _GEN7267;
wire  _GEN9646 = io_x[18] ? _GEN9645 : _GEN9641;
wire  _GEN9647 = io_x[33] ? _GEN9646 : _GEN9636;
wire  _GEN9648 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN9649 = io_x[18] ? _GEN9648 : _GEN7266;
wire  _GEN9650 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9651 = io_x[19] ? _GEN7273 : _GEN9650;
wire  _GEN9652 = io_x[23] ? _GEN9651 : _GEN7305;
wire  _GEN9653 = io_x[18] ? _GEN9652 : _GEN7266;
wire  _GEN9654 = io_x[33] ? _GEN9653 : _GEN9649;
wire  _GEN9655 = io_x[31] ? _GEN9654 : _GEN9647;
wire  _GEN9656 = io_x[28] ? _GEN9655 : _GEN9631;
wire  _GEN9657 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9658 = io_x[27] ? _GEN9657 : _GEN7278;
wire  _GEN9659 = io_x[19] ? _GEN9658 : _GEN7280;
wire  _GEN9660 = io_x[23] ? _GEN7267 : _GEN9659;
wire  _GEN9661 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9662 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN9663 = io_x[23] ? _GEN9662 : _GEN9661;
wire  _GEN9664 = io_x[18] ? _GEN9663 : _GEN9660;
wire  _GEN9665 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9666 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9667 = io_x[19] ? _GEN9666 : _GEN7280;
wire  _GEN9668 = io_x[23] ? _GEN9667 : _GEN9665;
wire  _GEN9669 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9670 = io_x[19] ? _GEN7273 : _GEN9669;
wire  _GEN9671 = io_x[23] ? _GEN7305 : _GEN9670;
wire  _GEN9672 = io_x[18] ? _GEN9671 : _GEN9668;
wire  _GEN9673 = io_x[33] ? _GEN9672 : _GEN9664;
wire  _GEN9674 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN9675 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9676 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9677 = io_x[27] ? _GEN9676 : _GEN7271;
wire  _GEN9678 = io_x[19] ? _GEN9677 : _GEN9675;
wire  _GEN9679 = io_x[23] ? _GEN9678 : _GEN9674;
wire  _GEN9680 = io_x[18] ? _GEN9679 : _GEN7297;
wire  _GEN9681 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9682 = io_x[19] ? _GEN7280 : _GEN9681;
wire  _GEN9683 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9684 = io_x[19] ? _GEN9683 : _GEN7273;
wire  _GEN9685 = io_x[23] ? _GEN9684 : _GEN9682;
wire  _GEN9686 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9687 = io_x[19] ? _GEN9686 : _GEN7280;
wire  _GEN9688 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9689 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9690 = io_x[19] ? _GEN9689 : _GEN9688;
wire  _GEN9691 = io_x[23] ? _GEN9690 : _GEN9687;
wire  _GEN9692 = io_x[18] ? _GEN9691 : _GEN9685;
wire  _GEN9693 = io_x[33] ? _GEN9692 : _GEN9680;
wire  _GEN9694 = io_x[31] ? _GEN9693 : _GEN9673;
wire  _GEN9695 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9696 = io_x[27] ? _GEN7278 : _GEN9695;
wire  _GEN9697 = io_x[19] ? _GEN9696 : _GEN7280;
wire  _GEN9698 = io_x[23] ? _GEN9697 : _GEN7305;
wire  _GEN9699 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9700 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9701 = io_x[27] ? _GEN7278 : _GEN9700;
wire  _GEN9702 = io_x[19] ? _GEN9701 : _GEN9699;
wire  _GEN9703 = io_x[23] ? _GEN9702 : _GEN7305;
wire  _GEN9704 = io_x[18] ? _GEN9703 : _GEN9698;
wire  _GEN9705 = io_x[33] ? _GEN9704 : _GEN8346;
wire  _GEN9706 = io_x[23] ? _GEN7267 : _GEN7305;
wire  _GEN9707 = io_x[18] ? _GEN9706 : _GEN7297;
wire  _GEN9708 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN9709 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9710 = io_x[19] ? _GEN9709 : _GEN7280;
wire  _GEN9711 = io_x[23] ? _GEN9710 : _GEN9708;
wire  _GEN9712 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9713 = io_x[19] ? _GEN7280 : _GEN9712;
wire  _GEN9714 = io_x[23] ? _GEN9713 : _GEN7305;
wire  _GEN9715 = io_x[18] ? _GEN9714 : _GEN9711;
wire  _GEN9716 = io_x[33] ? _GEN9715 : _GEN9707;
wire  _GEN9717 = io_x[31] ? _GEN9716 : _GEN9705;
wire  _GEN9718 = io_x[28] ? _GEN9717 : _GEN9694;
wire  _GEN9719 = io_x[26] ? _GEN9718 : _GEN9656;
wire  _GEN9720 = 1'b1;
wire  _GEN9721 = io_x[23] ? _GEN7267 : _GEN7305;
wire  _GEN9722 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9723 = io_x[27] ? _GEN9722 : _GEN7278;
wire  _GEN9724 = io_x[19] ? _GEN9723 : _GEN7280;
wire  _GEN9725 = io_x[23] ? _GEN9724 : _GEN7267;
wire  _GEN9726 = io_x[18] ? _GEN9725 : _GEN9721;
wire  _GEN9727 = io_x[33] ? _GEN9726 : _GEN9720;
wire  _GEN9728 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN9729 = io_x[23] ? _GEN9728 : _GEN7305;
wire  _GEN9730 = io_x[18] ? _GEN9729 : _GEN7266;
wire  _GEN9731 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9732 = io_x[27] ? _GEN9731 : _GEN7278;
wire  _GEN9733 = io_x[19] ? _GEN9732 : _GEN7280;
wire  _GEN9734 = io_x[23] ? _GEN9733 : _GEN7267;
wire  _GEN9735 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9736 = io_x[27] ? _GEN9735 : _GEN7278;
wire  _GEN9737 = io_x[19] ? _GEN9736 : _GEN7273;
wire  _GEN9738 = io_x[23] ? _GEN9737 : _GEN7267;
wire  _GEN9739 = io_x[18] ? _GEN9738 : _GEN9734;
wire  _GEN9740 = io_x[33] ? _GEN9739 : _GEN9730;
wire  _GEN9741 = io_x[31] ? _GEN9740 : _GEN9727;
wire  _GEN9742 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9743 = io_x[23] ? _GEN9742 : _GEN7305;
wire  _GEN9744 = io_x[18] ? _GEN9743 : _GEN7297;
wire  _GEN9745 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN9746 = io_x[23] ? _GEN7267 : _GEN9745;
wire  _GEN9747 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9748 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9749 = io_x[19] ? _GEN9748 : _GEN9747;
wire  _GEN9750 = io_x[23] ? _GEN9749 : _GEN7305;
wire  _GEN9751 = io_x[18] ? _GEN9750 : _GEN9746;
wire  _GEN9752 = io_x[33] ? _GEN9751 : _GEN9744;
wire  _GEN9753 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9754 = io_x[23] ? _GEN9753 : _GEN7267;
wire  _GEN9755 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9756 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9757 = io_x[27] ? _GEN9756 : _GEN9755;
wire  _GEN9758 = io_x[19] ? _GEN9757 : _GEN7273;
wire  _GEN9759 = io_x[23] ? _GEN9758 : _GEN7267;
wire  _GEN9760 = io_x[18] ? _GEN9759 : _GEN9754;
wire  _GEN9761 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9762 = io_x[27] ? _GEN9761 : _GEN7271;
wire  _GEN9763 = io_x[19] ? _GEN9762 : _GEN7273;
wire  _GEN9764 = io_x[23] ? _GEN9763 : _GEN7305;
wire  _GEN9765 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9766 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9767 = io_x[27] ? _GEN9766 : _GEN9765;
wire  _GEN9768 = io_x[19] ? _GEN9767 : _GEN7273;
wire  _GEN9769 = io_x[23] ? _GEN9768 : _GEN7267;
wire  _GEN9770 = io_x[18] ? _GEN9769 : _GEN9764;
wire  _GEN9771 = io_x[33] ? _GEN9770 : _GEN9760;
wire  _GEN9772 = io_x[31] ? _GEN9771 : _GEN9752;
wire  _GEN9773 = io_x[28] ? _GEN9772 : _GEN9741;
wire  _GEN9774 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9775 = io_x[19] ? _GEN7280 : _GEN9774;
wire  _GEN9776 = io_x[23] ? _GEN9775 : _GEN7267;
wire  _GEN9777 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9778 = io_x[19] ? _GEN7273 : _GEN9777;
wire  _GEN9779 = io_x[23] ? _GEN9778 : _GEN7267;
wire  _GEN9780 = io_x[18] ? _GEN9779 : _GEN9776;
wire  _GEN9781 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9782 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9783 = io_x[27] ? _GEN7278 : _GEN9782;
wire  _GEN9784 = io_x[19] ? _GEN7280 : _GEN9783;
wire  _GEN9785 = io_x[23] ? _GEN9784 : _GEN9781;
wire  _GEN9786 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9787 = io_x[19] ? _GEN9786 : _GEN7280;
wire  _GEN9788 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9789 = io_x[27] ? _GEN7271 : _GEN9788;
wire  _GEN9790 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9791 = io_x[19] ? _GEN9790 : _GEN9789;
wire  _GEN9792 = io_x[23] ? _GEN9791 : _GEN9787;
wire  _GEN9793 = io_x[18] ? _GEN9792 : _GEN9785;
wire  _GEN9794 = io_x[33] ? _GEN9793 : _GEN9780;
wire  _GEN9795 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9796 = io_x[23] ? _GEN9795 : _GEN7267;
wire  _GEN9797 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9798 = io_x[19] ? _GEN7280 : _GEN9797;
wire  _GEN9799 = io_x[23] ? _GEN9798 : _GEN7305;
wire  _GEN9800 = io_x[18] ? _GEN9799 : _GEN9796;
wire  _GEN9801 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9802 = io_x[27] ? _GEN7278 : _GEN9801;
wire  _GEN9803 = io_x[19] ? _GEN7273 : _GEN9802;
wire  _GEN9804 = io_x[23] ? _GEN9803 : _GEN7267;
wire  _GEN9805 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9806 = io_x[19] ? _GEN9805 : _GEN7273;
wire  _GEN9807 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9808 = io_x[27] ? _GEN9807 : _GEN7271;
wire  _GEN9809 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9810 = io_x[27] ? _GEN9809 : _GEN7278;
wire  _GEN9811 = io_x[19] ? _GEN9810 : _GEN9808;
wire  _GEN9812 = io_x[23] ? _GEN9811 : _GEN9806;
wire  _GEN9813 = io_x[18] ? _GEN9812 : _GEN9804;
wire  _GEN9814 = io_x[33] ? _GEN9813 : _GEN9800;
wire  _GEN9815 = io_x[31] ? _GEN9814 : _GEN9794;
wire  _GEN9816 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9817 = io_x[27] ? _GEN7278 : _GEN9816;
wire  _GEN9818 = io_x[19] ? _GEN7280 : _GEN9817;
wire  _GEN9819 = io_x[23] ? _GEN7305 : _GEN9818;
wire  _GEN9820 = io_x[18] ? _GEN9819 : _GEN7266;
wire  _GEN9821 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9822 = io_x[19] ? _GEN9821 : _GEN7280;
wire  _GEN9823 = io_x[23] ? _GEN7305 : _GEN9822;
wire  _GEN9824 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9825 = io_x[19] ? _GEN9824 : _GEN7280;
wire  _GEN9826 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9827 = io_x[27] ? _GEN9826 : _GEN7271;
wire  _GEN9828 = io_x[19] ? _GEN9827 : _GEN7273;
wire  _GEN9829 = io_x[23] ? _GEN9828 : _GEN9825;
wire  _GEN9830 = io_x[18] ? _GEN9829 : _GEN9823;
wire  _GEN9831 = io_x[33] ? _GEN9830 : _GEN9820;
wire  _GEN9832 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN9833 = io_x[23] ? _GEN9832 : _GEN7267;
wire  _GEN9834 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9835 = io_x[19] ? _GEN9834 : _GEN7280;
wire  _GEN9836 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9837 = io_x[23] ? _GEN9836 : _GEN9835;
wire  _GEN9838 = io_x[18] ? _GEN9837 : _GEN9833;
wire  _GEN9839 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9840 = io_x[27] ? _GEN9839 : _GEN7278;
wire  _GEN9841 = io_x[19] ? _GEN7280 : _GEN9840;
wire  _GEN9842 = io_x[23] ? _GEN9841 : _GEN7267;
wire  _GEN9843 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9844 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9845 = io_x[27] ? _GEN9844 : _GEN9843;
wire  _GEN9846 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9847 = io_x[27] ? _GEN9846 : _GEN7271;
wire  _GEN9848 = io_x[19] ? _GEN9847 : _GEN9845;
wire  _GEN9849 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9850 = io_x[27] ? _GEN9849 : _GEN7278;
wire  _GEN9851 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9852 = io_x[27] ? _GEN9851 : _GEN7271;
wire  _GEN9853 = io_x[19] ? _GEN9852 : _GEN9850;
wire  _GEN9854 = io_x[23] ? _GEN9853 : _GEN9848;
wire  _GEN9855 = io_x[18] ? _GEN9854 : _GEN9842;
wire  _GEN9856 = io_x[33] ? _GEN9855 : _GEN9838;
wire  _GEN9857 = io_x[31] ? _GEN9856 : _GEN9831;
wire  _GEN9858 = io_x[28] ? _GEN9857 : _GEN9815;
wire  _GEN9859 = io_x[26] ? _GEN9858 : _GEN9773;
wire  _GEN9860 = io_x[20] ? _GEN9859 : _GEN9719;
wire  _GEN9861 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9862 = io_x[27] ? _GEN9861 : _GEN7278;
wire  _GEN9863 = io_x[19] ? _GEN7273 : _GEN9862;
wire  _GEN9864 = io_x[23] ? _GEN7305 : _GEN9863;
wire  _GEN9865 = io_x[18] ? _GEN9864 : _GEN7297;
wire  _GEN9866 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9867 = io_x[19] ? _GEN9866 : _GEN7273;
wire  _GEN9868 = io_x[23] ? _GEN9867 : _GEN7305;
wire  _GEN9869 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9870 = io_x[27] ? _GEN9869 : _GEN7278;
wire  _GEN9871 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9872 = io_x[27] ? _GEN9871 : _GEN7278;
wire  _GEN9873 = io_x[19] ? _GEN9872 : _GEN9870;
wire  _GEN9874 = io_x[23] ? _GEN7267 : _GEN9873;
wire  _GEN9875 = io_x[18] ? _GEN9874 : _GEN9868;
wire  _GEN9876 = io_x[33] ? _GEN9875 : _GEN9865;
wire  _GEN9877 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN9878 = io_x[23] ? _GEN7267 : _GEN9877;
wire  _GEN9879 = io_x[18] ? _GEN9878 : _GEN7266;
wire  _GEN9880 = io_x[23] ? _GEN7305 : _GEN7267;
wire  _GEN9881 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9882 = io_x[27] ? _GEN9881 : _GEN7271;
wire  _GEN9883 = io_x[19] ? _GEN9882 : _GEN7273;
wire  _GEN9884 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9885 = io_x[27] ? _GEN9884 : _GEN7278;
wire  _GEN9886 = io_x[19] ? _GEN9885 : _GEN7280;
wire  _GEN9887 = io_x[23] ? _GEN9886 : _GEN9883;
wire  _GEN9888 = io_x[18] ? _GEN9887 : _GEN9880;
wire  _GEN9889 = io_x[33] ? _GEN9888 : _GEN9879;
wire  _GEN9890 = io_x[31] ? _GEN9889 : _GEN9876;
wire  _GEN9891 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9892 = io_x[23] ? _GEN7267 : _GEN9891;
wire  _GEN9893 = io_x[18] ? _GEN9892 : _GEN7297;
wire  _GEN9894 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9895 = io_x[19] ? _GEN9894 : _GEN7280;
wire  _GEN9896 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9897 = io_x[19] ? _GEN9896 : _GEN7280;
wire  _GEN9898 = io_x[23] ? _GEN9897 : _GEN9895;
wire  _GEN9899 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9900 = io_x[19] ? _GEN9899 : _GEN7273;
wire  _GEN9901 = io_x[23] ? _GEN9900 : _GEN7267;
wire  _GEN9902 = io_x[18] ? _GEN9901 : _GEN9898;
wire  _GEN9903 = io_x[33] ? _GEN9902 : _GEN9893;
wire  _GEN9904 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN9905 = io_x[23] ? _GEN7267 : _GEN9904;
wire  _GEN9906 = io_x[18] ? _GEN9905 : _GEN7266;
wire  _GEN9907 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN9908 = io_x[23] ? _GEN9907 : _GEN7267;
wire  _GEN9909 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9910 = io_x[19] ? _GEN7280 : _GEN9909;
wire  _GEN9911 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9912 = io_x[19] ? _GEN9911 : _GEN7280;
wire  _GEN9913 = io_x[23] ? _GEN9912 : _GEN9910;
wire  _GEN9914 = io_x[18] ? _GEN9913 : _GEN9908;
wire  _GEN9915 = io_x[33] ? _GEN9914 : _GEN9906;
wire  _GEN9916 = io_x[31] ? _GEN9915 : _GEN9903;
wire  _GEN9917 = io_x[28] ? _GEN9916 : _GEN9890;
wire  _GEN9918 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9919 = io_x[19] ? _GEN7273 : _GEN9918;
wire  _GEN9920 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9921 = io_x[23] ? _GEN9920 : _GEN9919;
wire  _GEN9922 = io_x[18] ? _GEN9921 : _GEN7297;
wire  _GEN9923 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9924 = io_x[19] ? _GEN9923 : _GEN7280;
wire  _GEN9925 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9926 = io_x[19] ? _GEN9925 : _GEN7280;
wire  _GEN9927 = io_x[23] ? _GEN9926 : _GEN9924;
wire  _GEN9928 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9929 = io_x[27] ? _GEN7278 : _GEN9928;
wire  _GEN9930 = io_x[19] ? _GEN7273 : _GEN9929;
wire  _GEN9931 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN9932 = io_x[23] ? _GEN9931 : _GEN9930;
wire  _GEN9933 = io_x[18] ? _GEN9932 : _GEN9927;
wire  _GEN9934 = io_x[33] ? _GEN9933 : _GEN9922;
wire  _GEN9935 = io_x[18] ? _GEN7297 : _GEN7266;
wire  _GEN9936 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9937 = io_x[19] ? _GEN9936 : _GEN7280;
wire  _GEN9938 = io_x[23] ? _GEN9937 : _GEN7267;
wire  _GEN9939 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9940 = io_x[27] ? _GEN7278 : _GEN9939;
wire  _GEN9941 = io_x[19] ? _GEN9940 : _GEN7273;
wire  _GEN9942 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9943 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9944 = io_x[19] ? _GEN9943 : _GEN9942;
wire  _GEN9945 = io_x[23] ? _GEN9944 : _GEN9941;
wire  _GEN9946 = io_x[18] ? _GEN9945 : _GEN9938;
wire  _GEN9947 = io_x[33] ? _GEN9946 : _GEN9935;
wire  _GEN9948 = io_x[31] ? _GEN9947 : _GEN9934;
wire  _GEN9949 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9950 = io_x[27] ? _GEN7278 : _GEN9949;
wire  _GEN9951 = io_x[19] ? _GEN9950 : _GEN7280;
wire  _GEN9952 = io_x[23] ? _GEN9951 : _GEN7267;
wire  _GEN9953 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9954 = io_x[27] ? _GEN9953 : _GEN7278;
wire  _GEN9955 = io_x[19] ? _GEN9954 : _GEN7273;
wire  _GEN9956 = io_x[23] ? _GEN9955 : _GEN7267;
wire  _GEN9957 = io_x[18] ? _GEN9956 : _GEN9952;
wire  _GEN9958 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9959 = io_x[27] ? _GEN7278 : _GEN9958;
wire  _GEN9960 = io_x[19] ? _GEN9959 : _GEN7280;
wire  _GEN9961 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9962 = io_x[19] ? _GEN9961 : _GEN7280;
wire  _GEN9963 = io_x[23] ? _GEN9962 : _GEN9960;
wire  _GEN9964 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9965 = io_x[27] ? _GEN7278 : _GEN9964;
wire  _GEN9966 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9967 = io_x[27] ? _GEN7278 : _GEN9966;
wire  _GEN9968 = io_x[19] ? _GEN9967 : _GEN9965;
wire  _GEN9969 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9970 = io_x[19] ? _GEN7280 : _GEN9969;
wire  _GEN9971 = io_x[23] ? _GEN9970 : _GEN9968;
wire  _GEN9972 = io_x[18] ? _GEN9971 : _GEN9963;
wire  _GEN9973 = io_x[33] ? _GEN9972 : _GEN9957;
wire  _GEN9974 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9975 = io_x[27] ? _GEN9974 : _GEN7278;
wire  _GEN9976 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN9977 = io_x[19] ? _GEN9976 : _GEN9975;
wire  _GEN9978 = io_x[23] ? _GEN9977 : _GEN7267;
wire  _GEN9979 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN9980 = io_x[19] ? _GEN9979 : _GEN7280;
wire  _GEN9981 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9982 = io_x[27] ? _GEN9981 : _GEN7278;
wire  _GEN9983 = io_x[19] ? _GEN9982 : _GEN7280;
wire  _GEN9984 = io_x[23] ? _GEN9983 : _GEN9980;
wire  _GEN9985 = io_x[18] ? _GEN9984 : _GEN9978;
wire  _GEN9986 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9987 = io_x[27] ? _GEN9986 : _GEN7278;
wire  _GEN9988 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9989 = io_x[27] ? _GEN9988 : _GEN7278;
wire  _GEN9990 = io_x[19] ? _GEN9989 : _GEN9987;
wire  _GEN9991 = io_x[23] ? _GEN9990 : _GEN7305;
wire  _GEN9992 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9993 = io_x[27] ? _GEN7271 : _GEN9992;
wire  _GEN9994 = io_x[19] ? _GEN7273 : _GEN9993;
wire  _GEN9995 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN9996 = io_x[27] ? _GEN9995 : _GEN7278;
wire  _GEN9997 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN9998 = io_x[27] ? _GEN9997 : _GEN7278;
wire  _GEN9999 = io_x[19] ? _GEN9998 : _GEN9996;
wire  _GEN10000 = io_x[23] ? _GEN9999 : _GEN9994;
wire  _GEN10001 = io_x[18] ? _GEN10000 : _GEN9991;
wire  _GEN10002 = io_x[33] ? _GEN10001 : _GEN9985;
wire  _GEN10003 = io_x[31] ? _GEN10002 : _GEN9973;
wire  _GEN10004 = io_x[28] ? _GEN10003 : _GEN9948;
wire  _GEN10005 = io_x[26] ? _GEN10004 : _GEN9917;
wire  _GEN10006 = io_x[23] ? _GEN7267 : _GEN7305;
wire  _GEN10007 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10008 = io_x[27] ? _GEN10007 : _GEN7278;
wire  _GEN10009 = io_x[19] ? _GEN7280 : _GEN10008;
wire  _GEN10010 = io_x[23] ? _GEN7305 : _GEN10009;
wire  _GEN10011 = io_x[18] ? _GEN10010 : _GEN10006;
wire  _GEN10012 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN10013 = io_x[19] ? _GEN7273 : _GEN10012;
wire  _GEN10014 = io_x[23] ? _GEN7267 : _GEN10013;
wire  _GEN10015 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10016 = io_x[27] ? _GEN10015 : _GEN7278;
wire  _GEN10017 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN10018 = io_x[19] ? _GEN10017 : _GEN10016;
wire  _GEN10019 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN10020 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10021 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10022 = io_x[27] ? _GEN10021 : _GEN10020;
wire  _GEN10023 = io_x[19] ? _GEN10022 : _GEN10019;
wire  _GEN10024 = io_x[23] ? _GEN10023 : _GEN10018;
wire  _GEN10025 = io_x[18] ? _GEN10024 : _GEN10014;
wire  _GEN10026 = io_x[33] ? _GEN10025 : _GEN10011;
wire  _GEN10027 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10028 = io_x[27] ? _GEN10027 : _GEN7278;
wire  _GEN10029 = io_x[19] ? _GEN7280 : _GEN10028;
wire  _GEN10030 = io_x[23] ? _GEN7267 : _GEN10029;
wire  _GEN10031 = io_x[18] ? _GEN10030 : _GEN7297;
wire  _GEN10032 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10033 = io_x[27] ? _GEN10032 : _GEN7278;
wire  _GEN10034 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN10035 = io_x[19] ? _GEN10034 : _GEN10033;
wire  _GEN10036 = io_x[23] ? _GEN10035 : _GEN7267;
wire  _GEN10037 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN10038 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN10039 = io_x[19] ? _GEN10038 : _GEN10037;
wire  _GEN10040 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN10041 = io_x[19] ? _GEN10040 : _GEN7280;
wire  _GEN10042 = io_x[23] ? _GEN10041 : _GEN10039;
wire  _GEN10043 = io_x[18] ? _GEN10042 : _GEN10036;
wire  _GEN10044 = io_x[33] ? _GEN10043 : _GEN10031;
wire  _GEN10045 = io_x[31] ? _GEN10044 : _GEN10026;
wire  _GEN10046 = io_x[19] ? _GEN7273 : _GEN7280;
wire  _GEN10047 = io_x[23] ? _GEN7267 : _GEN10046;
wire  _GEN10048 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10049 = io_x[27] ? _GEN10048 : _GEN7278;
wire  _GEN10050 = io_x[19] ? _GEN7273 : _GEN10049;
wire  _GEN10051 = io_x[23] ? _GEN7305 : _GEN10050;
wire  _GEN10052 = io_x[18] ? _GEN10051 : _GEN10047;
wire  _GEN10053 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN10054 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN10055 = io_x[19] ? _GEN10054 : _GEN10053;
wire  _GEN10056 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN10057 = io_x[19] ? _GEN10056 : _GEN7273;
wire  _GEN10058 = io_x[23] ? _GEN10057 : _GEN10055;
wire  _GEN10059 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN10060 = io_x[19] ? _GEN10059 : _GEN7280;
wire  _GEN10061 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN10062 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10063 = io_x[27] ? _GEN7278 : _GEN10062;
wire  _GEN10064 = io_x[19] ? _GEN10063 : _GEN10061;
wire  _GEN10065 = io_x[23] ? _GEN10064 : _GEN10060;
wire  _GEN10066 = io_x[18] ? _GEN10065 : _GEN10058;
wire  _GEN10067 = io_x[33] ? _GEN10066 : _GEN10052;
wire  _GEN10068 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN10069 = io_x[23] ? _GEN10068 : _GEN7267;
wire  _GEN10070 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10071 = io_x[27] ? _GEN10070 : _GEN7271;
wire  _GEN10072 = io_x[19] ? _GEN7280 : _GEN10071;
wire  _GEN10073 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN10074 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10075 = io_x[27] ? _GEN10074 : _GEN7278;
wire  _GEN10076 = io_x[19] ? _GEN10075 : _GEN10073;
wire  _GEN10077 = io_x[23] ? _GEN10076 : _GEN10072;
wire  _GEN10078 = io_x[18] ? _GEN10077 : _GEN10069;
wire  _GEN10079 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN10080 = io_x[19] ? _GEN10079 : _GEN7280;
wire  _GEN10081 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10082 = io_x[27] ? _GEN10081 : _GEN7278;
wire  _GEN10083 = io_x[19] ? _GEN7273 : _GEN10082;
wire  _GEN10084 = io_x[23] ? _GEN10083 : _GEN10080;
wire  _GEN10085 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10086 = io_x[27] ? _GEN7278 : _GEN10085;
wire  _GEN10087 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10088 = io_x[27] ? _GEN7278 : _GEN10087;
wire  _GEN10089 = io_x[19] ? _GEN10088 : _GEN10086;
wire  _GEN10090 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10091 = io_x[27] ? _GEN10090 : _GEN7271;
wire  _GEN10092 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10093 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10094 = io_x[27] ? _GEN10093 : _GEN10092;
wire  _GEN10095 = io_x[19] ? _GEN10094 : _GEN10091;
wire  _GEN10096 = io_x[23] ? _GEN10095 : _GEN10089;
wire  _GEN10097 = io_x[18] ? _GEN10096 : _GEN10084;
wire  _GEN10098 = io_x[33] ? _GEN10097 : _GEN10078;
wire  _GEN10099 = io_x[31] ? _GEN10098 : _GEN10067;
wire  _GEN10100 = io_x[28] ? _GEN10099 : _GEN10045;
wire  _GEN10101 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN10102 = io_x[19] ? _GEN7280 : _GEN10101;
wire  _GEN10103 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN10104 = io_x[19] ? _GEN7280 : _GEN10103;
wire  _GEN10105 = io_x[23] ? _GEN10104 : _GEN10102;
wire  _GEN10106 = io_x[18] ? _GEN10105 : _GEN7266;
wire  _GEN10107 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN10108 = io_x[19] ? _GEN10107 : _GEN7273;
wire  _GEN10109 = io_x[23] ? _GEN10108 : _GEN7305;
wire  _GEN10110 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN10111 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN10112 = io_x[19] ? _GEN10111 : _GEN10110;
wire  _GEN10113 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10114 = io_x[27] ? _GEN10113 : _GEN7278;
wire  _GEN10115 = io_x[19] ? _GEN10114 : _GEN7280;
wire  _GEN10116 = io_x[23] ? _GEN10115 : _GEN10112;
wire  _GEN10117 = io_x[18] ? _GEN10116 : _GEN10109;
wire  _GEN10118 = io_x[33] ? _GEN10117 : _GEN10106;
wire  _GEN10119 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN10120 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN10121 = io_x[19] ? _GEN10120 : _GEN7273;
wire  _GEN10122 = io_x[23] ? _GEN10121 : _GEN10119;
wire  _GEN10123 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10124 = io_x[27] ? _GEN10123 : _GEN7278;
wire  _GEN10125 = io_x[19] ? _GEN7280 : _GEN10124;
wire  _GEN10126 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10127 = io_x[27] ? _GEN10126 : _GEN7278;
wire  _GEN10128 = io_x[19] ? _GEN10127 : _GEN7280;
wire  _GEN10129 = io_x[23] ? _GEN10128 : _GEN10125;
wire  _GEN10130 = io_x[18] ? _GEN10129 : _GEN10122;
wire  _GEN10131 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10132 = io_x[27] ? _GEN10131 : _GEN7278;
wire  _GEN10133 = io_x[19] ? _GEN10132 : _GEN7273;
wire  _GEN10134 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN10135 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10136 = io_x[27] ? _GEN10135 : _GEN7278;
wire  _GEN10137 = io_x[19] ? _GEN10136 : _GEN10134;
wire  _GEN10138 = io_x[23] ? _GEN10137 : _GEN10133;
wire  _GEN10139 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10140 = io_x[27] ? _GEN10139 : _GEN7278;
wire  _GEN10141 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10142 = io_x[27] ? _GEN10141 : _GEN7271;
wire  _GEN10143 = io_x[19] ? _GEN10142 : _GEN10140;
wire  _GEN10144 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10145 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10146 = io_x[27] ? _GEN10145 : _GEN10144;
wire  _GEN10147 = io_x[19] ? _GEN10146 : _GEN7273;
wire  _GEN10148 = io_x[23] ? _GEN10147 : _GEN10143;
wire  _GEN10149 = io_x[18] ? _GEN10148 : _GEN10138;
wire  _GEN10150 = io_x[33] ? _GEN10149 : _GEN10130;
wire  _GEN10151 = io_x[31] ? _GEN10150 : _GEN10118;
wire  _GEN10152 = io_x[19] ? _GEN7280 : _GEN7273;
wire  _GEN10153 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10154 = io_x[27] ? _GEN10153 : _GEN7278;
wire  _GEN10155 = io_x[19] ? _GEN10154 : _GEN7280;
wire  _GEN10156 = io_x[23] ? _GEN10155 : _GEN10152;
wire  _GEN10157 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10158 = io_x[27] ? _GEN7278 : _GEN10157;
wire  _GEN10159 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10160 = io_x[27] ? _GEN7271 : _GEN10159;
wire  _GEN10161 = io_x[19] ? _GEN10160 : _GEN10158;
wire  _GEN10162 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN10163 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10164 = io_x[27] ? _GEN10163 : _GEN7278;
wire  _GEN10165 = io_x[19] ? _GEN10164 : _GEN10162;
wire  _GEN10166 = io_x[23] ? _GEN10165 : _GEN10161;
wire  _GEN10167 = io_x[18] ? _GEN10166 : _GEN10156;
wire  _GEN10168 = io_x[27] ? _GEN7278 : _GEN7271;
wire  _GEN10169 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10170 = io_x[27] ? _GEN7278 : _GEN10169;
wire  _GEN10171 = io_x[19] ? _GEN10170 : _GEN10168;
wire  _GEN10172 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10173 = io_x[27] ? _GEN7271 : _GEN10172;
wire  _GEN10174 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10175 = io_x[27] ? _GEN10174 : _GEN7271;
wire  _GEN10176 = io_x[19] ? _GEN10175 : _GEN10173;
wire  _GEN10177 = io_x[23] ? _GEN10176 : _GEN10171;
wire  _GEN10178 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10179 = io_x[27] ? _GEN7278 : _GEN10178;
wire  _GEN10180 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10181 = io_x[27] ? _GEN7271 : _GEN10180;
wire  _GEN10182 = io_x[19] ? _GEN10181 : _GEN10179;
wire  _GEN10183 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10184 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10185 = io_x[27] ? _GEN10184 : _GEN10183;
wire  _GEN10186 = io_x[19] ? _GEN10185 : _GEN7280;
wire  _GEN10187 = io_x[23] ? _GEN10186 : _GEN10182;
wire  _GEN10188 = io_x[18] ? _GEN10187 : _GEN10177;
wire  _GEN10189 = io_x[33] ? _GEN10188 : _GEN10167;
wire  _GEN10190 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10191 = io_x[27] ? _GEN10190 : _GEN7271;
wire  _GEN10192 = io_x[19] ? _GEN10191 : _GEN7273;
wire  _GEN10193 = io_x[23] ? _GEN10192 : _GEN7305;
wire  _GEN10194 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10195 = io_x[27] ? _GEN7271 : _GEN10194;
wire  _GEN10196 = io_x[19] ? _GEN7280 : _GEN10195;
wire  _GEN10197 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10198 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10199 = io_x[27] ? _GEN10198 : _GEN10197;
wire  _GEN10200 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10201 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10202 = io_x[27] ? _GEN10201 : _GEN10200;
wire  _GEN10203 = io_x[19] ? _GEN10202 : _GEN10199;
wire  _GEN10204 = io_x[23] ? _GEN10203 : _GEN10196;
wire  _GEN10205 = io_x[18] ? _GEN10204 : _GEN10193;
wire  _GEN10206 = io_x[27] ? _GEN7271 : _GEN7278;
wire  _GEN10207 = io_x[19] ? _GEN7273 : _GEN10206;
wire  _GEN10208 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10209 = io_x[27] ? _GEN10208 : _GEN7271;
wire  _GEN10210 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10211 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10212 = io_x[27] ? _GEN10211 : _GEN10210;
wire  _GEN10213 = io_x[19] ? _GEN10212 : _GEN10209;
wire  _GEN10214 = io_x[23] ? _GEN10213 : _GEN10207;
wire  _GEN10215 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10216 = io_x[27] ? _GEN7271 : _GEN10215;
wire  _GEN10217 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10218 = io_x[27] ? _GEN10217 : _GEN7271;
wire  _GEN10219 = io_x[19] ? _GEN10218 : _GEN10216;
wire  _GEN10220 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10221 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10222 = io_x[27] ? _GEN10221 : _GEN10220;
wire  _GEN10223 = io_x[77] ? _GEN7269 : _GEN7268;
wire  _GEN10224 = io_x[77] ? _GEN7268 : _GEN7269;
wire  _GEN10225 = io_x[27] ? _GEN10224 : _GEN10223;
wire  _GEN10226 = io_x[19] ? _GEN10225 : _GEN10222;
wire  _GEN10227 = io_x[23] ? _GEN10226 : _GEN10219;
wire  _GEN10228 = io_x[18] ? _GEN10227 : _GEN10214;
wire  _GEN10229 = io_x[33] ? _GEN10228 : _GEN10205;
wire  _GEN10230 = io_x[31] ? _GEN10229 : _GEN10189;
wire  _GEN10231 = io_x[28] ? _GEN10230 : _GEN10151;
wire  _GEN10232 = io_x[26] ? _GEN10231 : _GEN10100;
wire  _GEN10233 = io_x[20] ? _GEN10232 : _GEN10005;
wire  _GEN10234 = io_x[24] ? _GEN10233 : _GEN9860;
wire  _GEN10235 = io_x[78] ? _GEN10234 : _GEN9603;
wire  _GEN10236 = io_x[72] ? _GEN10235 : _GEN8795;
assign io_y[9] = _GEN10236;
wire  _GEN10237 = 1'b1;
wire  _GEN10238 = 1'b0;
wire  _GEN10239 = 1'b1;
wire  _GEN10240 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10241 = 1'b1;
wire  _GEN10242 = io_x[26] ? _GEN10241 : _GEN10240;
wire  _GEN10243 = 1'b1;
wire  _GEN10244 = io_x[73] ? _GEN10243 : _GEN10242;
wire  _GEN10245 = io_x[33] ? _GEN10244 : _GEN10237;
wire  _GEN10246 = 1'b0;
wire  _GEN10247 = 1'b0;
wire  _GEN10248 = 1'b1;
wire  _GEN10249 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10250 = io_x[30] ? _GEN10249 : _GEN10239;
wire  _GEN10251 = io_x[26] ? _GEN10250 : _GEN10246;
wire  _GEN10252 = io_x[73] ? _GEN10243 : _GEN10251;
wire  _GEN10253 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10254 = io_x[30] ? _GEN10253 : _GEN10239;
wire  _GEN10255 = io_x[26] ? _GEN10254 : _GEN10246;
wire  _GEN10256 = io_x[73] ? _GEN10243 : _GEN10255;
wire  _GEN10257 = io_x[33] ? _GEN10256 : _GEN10252;
wire  _GEN10258 = io_x[28] ? _GEN10257 : _GEN10245;
wire  _GEN10259 = 1'b0;
wire  _GEN10260 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10261 = io_x[73] ? _GEN10260 : _GEN10259;
wire  _GEN10262 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10263 = io_x[30] ? _GEN10262 : _GEN10239;
wire  _GEN10264 = io_x[26] ? _GEN10263 : _GEN10246;
wire  _GEN10265 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10266 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10267 = io_x[30] ? _GEN10266 : _GEN10265;
wire  _GEN10268 = io_x[26] ? _GEN10246 : _GEN10267;
wire  _GEN10269 = io_x[73] ? _GEN10268 : _GEN10264;
wire  _GEN10270 = io_x[33] ? _GEN10269 : _GEN10261;
wire  _GEN10271 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10272 = io_x[26] ? _GEN10271 : _GEN10241;
wire  _GEN10273 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10274 = io_x[73] ? _GEN10273 : _GEN10272;
wire  _GEN10275 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10276 = io_x[30] ? _GEN10275 : _GEN10239;
wire  _GEN10277 = io_x[26] ? _GEN10276 : _GEN10241;
wire  _GEN10278 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10279 = io_x[30] ? _GEN10278 : _GEN10239;
wire  _GEN10280 = io_x[26] ? _GEN10246 : _GEN10279;
wire  _GEN10281 = io_x[73] ? _GEN10280 : _GEN10277;
wire  _GEN10282 = io_x[33] ? _GEN10281 : _GEN10274;
wire  _GEN10283 = io_x[28] ? _GEN10282 : _GEN10270;
wire  _GEN10284 = io_x[18] ? _GEN10283 : _GEN10258;
wire  _GEN10285 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10286 = io_x[26] ? _GEN10285 : _GEN10241;
wire  _GEN10287 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10288 = io_x[26] ? _GEN10287 : _GEN10241;
wire  _GEN10289 = io_x[73] ? _GEN10288 : _GEN10286;
wire  _GEN10290 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10291 = io_x[30] ? _GEN10290 : _GEN10238;
wire  _GEN10292 = io_x[26] ? _GEN10291 : _GEN10241;
wire  _GEN10293 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10294 = io_x[26] ? _GEN10293 : _GEN10241;
wire  _GEN10295 = io_x[73] ? _GEN10294 : _GEN10292;
wire  _GEN10296 = io_x[33] ? _GEN10295 : _GEN10289;
wire  _GEN10297 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10298 = io_x[30] ? _GEN10297 : _GEN10239;
wire  _GEN10299 = io_x[26] ? _GEN10298 : _GEN10246;
wire  _GEN10300 = io_x[73] ? _GEN10243 : _GEN10299;
wire  _GEN10301 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10302 = io_x[26] ? _GEN10301 : _GEN10246;
wire  _GEN10303 = io_x[73] ? _GEN10259 : _GEN10302;
wire  _GEN10304 = io_x[33] ? _GEN10303 : _GEN10300;
wire  _GEN10305 = io_x[28] ? _GEN10304 : _GEN10296;
wire  _GEN10306 = 1'b0;
wire  _GEN10307 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10308 = io_x[30] ? _GEN10307 : _GEN10239;
wire  _GEN10309 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10310 = io_x[30] ? _GEN10309 : _GEN10239;
wire  _GEN10311 = io_x[26] ? _GEN10310 : _GEN10308;
wire  _GEN10312 = io_x[73] ? _GEN10259 : _GEN10311;
wire  _GEN10313 = io_x[33] ? _GEN10312 : _GEN10306;
wire  _GEN10314 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10315 = io_x[30] ? _GEN10314 : _GEN10239;
wire  _GEN10316 = io_x[26] ? _GEN10315 : _GEN10241;
wire  _GEN10317 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10318 = io_x[73] ? _GEN10317 : _GEN10316;
wire  _GEN10319 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10320 = io_x[30] ? _GEN10319 : _GEN10238;
wire  _GEN10321 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10322 = io_x[26] ? _GEN10321 : _GEN10320;
wire  _GEN10323 = io_x[73] ? _GEN10322 : _GEN10259;
wire  _GEN10324 = io_x[33] ? _GEN10323 : _GEN10318;
wire  _GEN10325 = io_x[28] ? _GEN10324 : _GEN10313;
wire  _GEN10326 = io_x[18] ? _GEN10325 : _GEN10305;
wire  _GEN10327 = io_x[25] ? _GEN10326 : _GEN10284;
wire  _GEN10328 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10329 = io_x[73] ? _GEN10259 : _GEN10328;
wire  _GEN10330 = io_x[33] ? _GEN10329 : _GEN10306;
wire  _GEN10331 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10332 = io_x[30] ? _GEN10239 : _GEN10331;
wire  _GEN10333 = io_x[26] ? _GEN10246 : _GEN10332;
wire  _GEN10334 = io_x[73] ? _GEN10243 : _GEN10333;
wire  _GEN10335 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10336 = io_x[30] ? _GEN10239 : _GEN10335;
wire  _GEN10337 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10338 = io_x[26] ? _GEN10337 : _GEN10336;
wire  _GEN10339 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10340 = io_x[30] ? _GEN10339 : _GEN10239;
wire  _GEN10341 = io_x[26] ? _GEN10340 : _GEN10241;
wire  _GEN10342 = io_x[73] ? _GEN10341 : _GEN10338;
wire  _GEN10343 = io_x[33] ? _GEN10342 : _GEN10334;
wire  _GEN10344 = io_x[28] ? _GEN10343 : _GEN10330;
wire  _GEN10345 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10346 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN10347 = io_x[73] ? _GEN10346 : _GEN10345;
wire  _GEN10348 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10349 = io_x[26] ? _GEN10348 : _GEN10246;
wire  _GEN10350 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10351 = io_x[26] ? _GEN10350 : _GEN10241;
wire  _GEN10352 = io_x[73] ? _GEN10351 : _GEN10349;
wire  _GEN10353 = io_x[33] ? _GEN10352 : _GEN10347;
wire  _GEN10354 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10355 = io_x[26] ? _GEN10354 : _GEN10246;
wire  _GEN10356 = io_x[73] ? _GEN10355 : _GEN10259;
wire  _GEN10357 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10358 = io_x[30] ? _GEN10357 : _GEN10238;
wire  _GEN10359 = io_x[26] ? _GEN10358 : _GEN10241;
wire  _GEN10360 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10361 = io_x[26] ? _GEN10360 : _GEN10241;
wire  _GEN10362 = io_x[73] ? _GEN10361 : _GEN10359;
wire  _GEN10363 = io_x[33] ? _GEN10362 : _GEN10356;
wire  _GEN10364 = io_x[28] ? _GEN10363 : _GEN10353;
wire  _GEN10365 = io_x[18] ? _GEN10364 : _GEN10344;
wire  _GEN10366 = io_x[73] ? _GEN10259 : _GEN10243;
wire  _GEN10367 = io_x[33] ? _GEN10366 : _GEN10237;
wire  _GEN10368 = io_x[73] ? _GEN10243 : _GEN10259;
wire  _GEN10369 = io_x[33] ? _GEN10368 : _GEN10237;
wire  _GEN10370 = io_x[28] ? _GEN10369 : _GEN10367;
wire  _GEN10371 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10372 = io_x[26] ? _GEN10371 : _GEN10241;
wire  _GEN10373 = io_x[73] ? _GEN10259 : _GEN10372;
wire  _GEN10374 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10375 = io_x[30] ? _GEN10374 : _GEN10239;
wire  _GEN10376 = io_x[26] ? _GEN10246 : _GEN10375;
wire  _GEN10377 = io_x[73] ? _GEN10243 : _GEN10376;
wire  _GEN10378 = io_x[33] ? _GEN10377 : _GEN10373;
wire  _GEN10379 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10380 = io_x[30] ? _GEN10379 : _GEN10239;
wire  _GEN10381 = io_x[26] ? _GEN10380 : _GEN10241;
wire  _GEN10382 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10383 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10384 = io_x[26] ? _GEN10383 : _GEN10382;
wire  _GEN10385 = io_x[73] ? _GEN10384 : _GEN10381;
wire  _GEN10386 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10387 = io_x[30] ? _GEN10386 : _GEN10239;
wire  _GEN10388 = io_x[26] ? _GEN10387 : _GEN10241;
wire  _GEN10389 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10390 = io_x[30] ? _GEN10238 : _GEN10389;
wire  _GEN10391 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10392 = io_x[26] ? _GEN10391 : _GEN10390;
wire  _GEN10393 = io_x[73] ? _GEN10392 : _GEN10388;
wire  _GEN10394 = io_x[33] ? _GEN10393 : _GEN10385;
wire  _GEN10395 = io_x[28] ? _GEN10394 : _GEN10378;
wire  _GEN10396 = io_x[18] ? _GEN10395 : _GEN10370;
wire  _GEN10397 = io_x[25] ? _GEN10396 : _GEN10365;
wire  _GEN10398 = io_x[29] ? _GEN10397 : _GEN10327;
wire  _GEN10399 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10400 = io_x[73] ? _GEN10243 : _GEN10399;
wire  _GEN10401 = io_x[33] ? _GEN10400 : _GEN10237;
wire  _GEN10402 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10403 = io_x[73] ? _GEN10243 : _GEN10402;
wire  _GEN10404 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10405 = io_x[30] ? _GEN10404 : _GEN10239;
wire  _GEN10406 = io_x[26] ? _GEN10246 : _GEN10405;
wire  _GEN10407 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10408 = io_x[73] ? _GEN10407 : _GEN10406;
wire  _GEN10409 = io_x[33] ? _GEN10408 : _GEN10403;
wire  _GEN10410 = io_x[28] ? _GEN10409 : _GEN10401;
wire  _GEN10411 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10412 = io_x[30] ? _GEN10411 : _GEN10239;
wire  _GEN10413 = io_x[26] ? _GEN10412 : _GEN10246;
wire  _GEN10414 = io_x[73] ? _GEN10243 : _GEN10413;
wire  _GEN10415 = io_x[33] ? _GEN10306 : _GEN10414;
wire  _GEN10416 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10417 = io_x[26] ? _GEN10416 : _GEN10241;
wire  _GEN10418 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10419 = io_x[30] ? _GEN10238 : _GEN10418;
wire  _GEN10420 = io_x[26] ? _GEN10419 : _GEN10241;
wire  _GEN10421 = io_x[73] ? _GEN10420 : _GEN10417;
wire  _GEN10422 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10423 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10424 = io_x[30] ? _GEN10423 : _GEN10422;
wire  _GEN10425 = io_x[26] ? _GEN10424 : _GEN10241;
wire  _GEN10426 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10427 = io_x[30] ? _GEN10238 : _GEN10426;
wire  _GEN10428 = io_x[26] ? _GEN10427 : _GEN10246;
wire  _GEN10429 = io_x[73] ? _GEN10428 : _GEN10425;
wire  _GEN10430 = io_x[33] ? _GEN10429 : _GEN10421;
wire  _GEN10431 = io_x[28] ? _GEN10430 : _GEN10415;
wire  _GEN10432 = io_x[18] ? _GEN10431 : _GEN10410;
wire  _GEN10433 = 1'b1;
wire  _GEN10434 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN10435 = io_x[73] ? _GEN10434 : _GEN10243;
wire  _GEN10436 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10437 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10438 = io_x[30] ? _GEN10437 : _GEN10436;
wire  _GEN10439 = io_x[26] ? _GEN10438 : _GEN10241;
wire  _GEN10440 = io_x[73] ? _GEN10243 : _GEN10439;
wire  _GEN10441 = io_x[33] ? _GEN10440 : _GEN10435;
wire  _GEN10442 = io_x[28] ? _GEN10441 : _GEN10433;
wire  _GEN10443 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10444 = io_x[73] ? _GEN10243 : _GEN10443;
wire  _GEN10445 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10446 = io_x[73] ? _GEN10445 : _GEN10259;
wire  _GEN10447 = io_x[33] ? _GEN10446 : _GEN10444;
wire  _GEN10448 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10449 = io_x[30] ? _GEN10448 : _GEN10239;
wire  _GEN10450 = io_x[26] ? _GEN10246 : _GEN10449;
wire  _GEN10451 = io_x[73] ? _GEN10259 : _GEN10450;
wire  _GEN10452 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10453 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10454 = io_x[30] ? _GEN10238 : _GEN10453;
wire  _GEN10455 = io_x[26] ? _GEN10454 : _GEN10452;
wire  _GEN10456 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10457 = io_x[26] ? _GEN10246 : _GEN10456;
wire  _GEN10458 = io_x[73] ? _GEN10457 : _GEN10455;
wire  _GEN10459 = io_x[33] ? _GEN10458 : _GEN10451;
wire  _GEN10460 = io_x[28] ? _GEN10459 : _GEN10447;
wire  _GEN10461 = io_x[18] ? _GEN10460 : _GEN10442;
wire  _GEN10462 = io_x[25] ? _GEN10461 : _GEN10432;
wire  _GEN10463 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10464 = io_x[30] ? _GEN10238 : _GEN10463;
wire  _GEN10465 = io_x[26] ? _GEN10464 : _GEN10241;
wire  _GEN10466 = io_x[73] ? _GEN10243 : _GEN10465;
wire  _GEN10467 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10468 = io_x[26] ? _GEN10467 : _GEN10241;
wire  _GEN10469 = io_x[73] ? _GEN10243 : _GEN10468;
wire  _GEN10470 = io_x[33] ? _GEN10469 : _GEN10466;
wire  _GEN10471 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10472 = io_x[30] ? _GEN10238 : _GEN10471;
wire  _GEN10473 = io_x[26] ? _GEN10472 : _GEN10241;
wire  _GEN10474 = io_x[73] ? _GEN10259 : _GEN10473;
wire  _GEN10475 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10476 = io_x[30] ? _GEN10239 : _GEN10475;
wire  _GEN10477 = io_x[26] ? _GEN10476 : _GEN10241;
wire  _GEN10478 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10479 = io_x[30] ? _GEN10478 : _GEN10238;
wire  _GEN10480 = io_x[26] ? _GEN10479 : _GEN10246;
wire  _GEN10481 = io_x[73] ? _GEN10480 : _GEN10477;
wire  _GEN10482 = io_x[33] ? _GEN10481 : _GEN10474;
wire  _GEN10483 = io_x[28] ? _GEN10482 : _GEN10470;
wire  _GEN10484 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10485 = io_x[26] ? _GEN10484 : _GEN10246;
wire  _GEN10486 = io_x[73] ? _GEN10485 : _GEN10259;
wire  _GEN10487 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10488 = io_x[30] ? _GEN10487 : _GEN10238;
wire  _GEN10489 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10490 = io_x[26] ? _GEN10489 : _GEN10488;
wire  _GEN10491 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN10492 = io_x[73] ? _GEN10491 : _GEN10490;
wire  _GEN10493 = io_x[33] ? _GEN10492 : _GEN10486;
wire  _GEN10494 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10495 = io_x[30] ? _GEN10494 : _GEN10239;
wire  _GEN10496 = io_x[26] ? _GEN10495 : _GEN10241;
wire  _GEN10497 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10498 = io_x[30] ? _GEN10497 : _GEN10239;
wire  _GEN10499 = io_x[26] ? _GEN10498 : _GEN10241;
wire  _GEN10500 = io_x[73] ? _GEN10499 : _GEN10496;
wire  _GEN10501 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10502 = io_x[30] ? _GEN10501 : _GEN10239;
wire  _GEN10503 = io_x[26] ? _GEN10502 : _GEN10241;
wire  _GEN10504 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10505 = io_x[26] ? _GEN10241 : _GEN10504;
wire  _GEN10506 = io_x[73] ? _GEN10505 : _GEN10503;
wire  _GEN10507 = io_x[33] ? _GEN10506 : _GEN10500;
wire  _GEN10508 = io_x[28] ? _GEN10507 : _GEN10493;
wire  _GEN10509 = io_x[18] ? _GEN10508 : _GEN10483;
wire  _GEN10510 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10511 = io_x[30] ? _GEN10238 : _GEN10510;
wire  _GEN10512 = io_x[26] ? _GEN10246 : _GEN10511;
wire  _GEN10513 = io_x[73] ? _GEN10243 : _GEN10512;
wire  _GEN10514 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10515 = io_x[30] ? _GEN10238 : _GEN10514;
wire  _GEN10516 = io_x[26] ? _GEN10241 : _GEN10515;
wire  _GEN10517 = io_x[73] ? _GEN10243 : _GEN10516;
wire  _GEN10518 = io_x[33] ? _GEN10517 : _GEN10513;
wire  _GEN10519 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10520 = io_x[26] ? _GEN10519 : _GEN10246;
wire  _GEN10521 = io_x[73] ? _GEN10243 : _GEN10520;
wire  _GEN10522 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10523 = io_x[30] ? _GEN10522 : _GEN10238;
wire  _GEN10524 = io_x[26] ? _GEN10523 : _GEN10241;
wire  _GEN10525 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10526 = io_x[26] ? _GEN10246 : _GEN10525;
wire  _GEN10527 = io_x[73] ? _GEN10526 : _GEN10524;
wire  _GEN10528 = io_x[33] ? _GEN10527 : _GEN10521;
wire  _GEN10529 = io_x[28] ? _GEN10528 : _GEN10518;
wire  _GEN10530 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10531 = io_x[30] ? _GEN10530 : _GEN10239;
wire  _GEN10532 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10533 = io_x[30] ? _GEN10238 : _GEN10532;
wire  _GEN10534 = io_x[26] ? _GEN10533 : _GEN10531;
wire  _GEN10535 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10536 = io_x[26] ? _GEN10246 : _GEN10535;
wire  _GEN10537 = io_x[73] ? _GEN10536 : _GEN10534;
wire  _GEN10538 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10539 = io_x[26] ? _GEN10246 : _GEN10538;
wire  _GEN10540 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10541 = io_x[30] ? _GEN10239 : _GEN10540;
wire  _GEN10542 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10543 = io_x[26] ? _GEN10542 : _GEN10541;
wire  _GEN10544 = io_x[73] ? _GEN10543 : _GEN10539;
wire  _GEN10545 = io_x[33] ? _GEN10544 : _GEN10537;
wire  _GEN10546 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10547 = io_x[26] ? _GEN10546 : _GEN10241;
wire  _GEN10548 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10549 = io_x[30] ? _GEN10548 : _GEN10239;
wire  _GEN10550 = io_x[26] ? _GEN10549 : _GEN10246;
wire  _GEN10551 = io_x[73] ? _GEN10550 : _GEN10547;
wire  _GEN10552 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10553 = io_x[30] ? _GEN10552 : _GEN10239;
wire  _GEN10554 = io_x[26] ? _GEN10553 : _GEN10241;
wire  _GEN10555 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10556 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10557 = io_x[26] ? _GEN10556 : _GEN10555;
wire  _GEN10558 = io_x[73] ? _GEN10557 : _GEN10554;
wire  _GEN10559 = io_x[33] ? _GEN10558 : _GEN10551;
wire  _GEN10560 = io_x[28] ? _GEN10559 : _GEN10545;
wire  _GEN10561 = io_x[18] ? _GEN10560 : _GEN10529;
wire  _GEN10562 = io_x[25] ? _GEN10561 : _GEN10509;
wire  _GEN10563 = io_x[29] ? _GEN10562 : _GEN10462;
wire  _GEN10564 = io_x[23] ? _GEN10563 : _GEN10398;
wire  _GEN10565 = io_x[73] ? _GEN10243 : _GEN10259;
wire  _GEN10566 = io_x[33] ? _GEN10306 : _GEN10565;
wire  _GEN10567 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10568 = io_x[26] ? _GEN10241 : _GEN10567;
wire  _GEN10569 = io_x[73] ? _GEN10243 : _GEN10568;
wire  _GEN10570 = io_x[33] ? _GEN10306 : _GEN10569;
wire  _GEN10571 = io_x[28] ? _GEN10570 : _GEN10566;
wire  _GEN10572 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10573 = io_x[26] ? _GEN10572 : _GEN10241;
wire  _GEN10574 = io_x[73] ? _GEN10259 : _GEN10573;
wire  _GEN10575 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10576 = io_x[26] ? _GEN10246 : _GEN10575;
wire  _GEN10577 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10578 = io_x[30] ? _GEN10577 : _GEN10239;
wire  _GEN10579 = io_x[26] ? _GEN10578 : _GEN10246;
wire  _GEN10580 = io_x[73] ? _GEN10579 : _GEN10576;
wire  _GEN10581 = io_x[33] ? _GEN10580 : _GEN10574;
wire  _GEN10582 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10583 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10584 = io_x[30] ? _GEN10583 : _GEN10239;
wire  _GEN10585 = io_x[26] ? _GEN10584 : _GEN10582;
wire  _GEN10586 = io_x[73] ? _GEN10259 : _GEN10585;
wire  _GEN10587 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10588 = io_x[30] ? _GEN10239 : _GEN10587;
wire  _GEN10589 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10590 = io_x[30] ? _GEN10589 : _GEN10239;
wire  _GEN10591 = io_x[26] ? _GEN10590 : _GEN10588;
wire  _GEN10592 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10593 = io_x[26] ? _GEN10592 : _GEN10241;
wire  _GEN10594 = io_x[73] ? _GEN10593 : _GEN10591;
wire  _GEN10595 = io_x[33] ? _GEN10594 : _GEN10586;
wire  _GEN10596 = io_x[28] ? _GEN10595 : _GEN10581;
wire  _GEN10597 = io_x[18] ? _GEN10596 : _GEN10571;
wire  _GEN10598 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10599 = io_x[30] ? _GEN10598 : _GEN10239;
wire  _GEN10600 = io_x[26] ? _GEN10599 : _GEN10241;
wire  _GEN10601 = io_x[73] ? _GEN10259 : _GEN10600;
wire  _GEN10602 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10603 = io_x[30] ? _GEN10239 : _GEN10602;
wire  _GEN10604 = io_x[26] ? _GEN10603 : _GEN10241;
wire  _GEN10605 = io_x[73] ? _GEN10243 : _GEN10604;
wire  _GEN10606 = io_x[33] ? _GEN10605 : _GEN10601;
wire  _GEN10607 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10608 = io_x[30] ? _GEN10239 : _GEN10607;
wire  _GEN10609 = io_x[26] ? _GEN10246 : _GEN10608;
wire  _GEN10610 = io_x[73] ? _GEN10243 : _GEN10609;
wire  _GEN10611 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10612 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10613 = io_x[26] ? _GEN10612 : _GEN10611;
wire  _GEN10614 = io_x[73] ? _GEN10243 : _GEN10613;
wire  _GEN10615 = io_x[33] ? _GEN10614 : _GEN10610;
wire  _GEN10616 = io_x[28] ? _GEN10615 : _GEN10606;
wire  _GEN10617 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10618 = io_x[30] ? _GEN10617 : _GEN10239;
wire  _GEN10619 = io_x[26] ? _GEN10618 : _GEN10241;
wire  _GEN10620 = io_x[73] ? _GEN10619 : _GEN10243;
wire  _GEN10621 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10622 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10623 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10624 = io_x[30] ? _GEN10623 : _GEN10622;
wire  _GEN10625 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10626 = io_x[26] ? _GEN10625 : _GEN10624;
wire  _GEN10627 = io_x[73] ? _GEN10626 : _GEN10621;
wire  _GEN10628 = io_x[33] ? _GEN10627 : _GEN10620;
wire  _GEN10629 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10630 = io_x[26] ? _GEN10629 : _GEN10241;
wire  _GEN10631 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10632 = io_x[30] ? _GEN10631 : _GEN10239;
wire  _GEN10633 = io_x[26] ? _GEN10632 : _GEN10246;
wire  _GEN10634 = io_x[73] ? _GEN10633 : _GEN10630;
wire  _GEN10635 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10636 = io_x[30] ? _GEN10635 : _GEN10239;
wire  _GEN10637 = io_x[26] ? _GEN10636 : _GEN10241;
wire  _GEN10638 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10639 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10640 = io_x[30] ? _GEN10639 : _GEN10239;
wire  _GEN10641 = io_x[26] ? _GEN10640 : _GEN10638;
wire  _GEN10642 = io_x[73] ? _GEN10641 : _GEN10637;
wire  _GEN10643 = io_x[33] ? _GEN10642 : _GEN10634;
wire  _GEN10644 = io_x[28] ? _GEN10643 : _GEN10628;
wire  _GEN10645 = io_x[18] ? _GEN10644 : _GEN10616;
wire  _GEN10646 = io_x[25] ? _GEN10645 : _GEN10597;
wire  _GEN10647 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10648 = io_x[26] ? _GEN10241 : _GEN10647;
wire  _GEN10649 = io_x[73] ? _GEN10648 : _GEN10259;
wire  _GEN10650 = io_x[33] ? _GEN10649 : _GEN10237;
wire  _GEN10651 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10652 = io_x[30] ? _GEN10651 : _GEN10239;
wire  _GEN10653 = io_x[26] ? _GEN10652 : _GEN10241;
wire  _GEN10654 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10655 = io_x[73] ? _GEN10654 : _GEN10653;
wire  _GEN10656 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10657 = io_x[26] ? _GEN10656 : _GEN10241;
wire  _GEN10658 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10659 = io_x[30] ? _GEN10658 : _GEN10238;
wire  _GEN10660 = io_x[26] ? _GEN10659 : _GEN10241;
wire  _GEN10661 = io_x[73] ? _GEN10660 : _GEN10657;
wire  _GEN10662 = io_x[33] ? _GEN10661 : _GEN10655;
wire  _GEN10663 = io_x[28] ? _GEN10662 : _GEN10650;
wire  _GEN10664 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10665 = io_x[26] ? _GEN10664 : _GEN10241;
wire  _GEN10666 = io_x[73] ? _GEN10243 : _GEN10665;
wire  _GEN10667 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10668 = io_x[30] ? _GEN10667 : _GEN10239;
wire  _GEN10669 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10670 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10671 = io_x[30] ? _GEN10670 : _GEN10669;
wire  _GEN10672 = io_x[26] ? _GEN10671 : _GEN10668;
wire  _GEN10673 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10674 = io_x[26] ? _GEN10673 : _GEN10246;
wire  _GEN10675 = io_x[73] ? _GEN10674 : _GEN10672;
wire  _GEN10676 = io_x[33] ? _GEN10675 : _GEN10666;
wire  _GEN10677 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10678 = io_x[30] ? _GEN10239 : _GEN10677;
wire  _GEN10679 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10680 = io_x[30] ? _GEN10679 : _GEN10239;
wire  _GEN10681 = io_x[26] ? _GEN10680 : _GEN10678;
wire  _GEN10682 = io_x[73] ? _GEN10259 : _GEN10681;
wire  _GEN10683 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10684 = io_x[30] ? _GEN10683 : _GEN10238;
wire  _GEN10685 = io_x[26] ? _GEN10246 : _GEN10684;
wire  _GEN10686 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10687 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10688 = io_x[30] ? _GEN10687 : _GEN10239;
wire  _GEN10689 = io_x[26] ? _GEN10688 : _GEN10686;
wire  _GEN10690 = io_x[73] ? _GEN10689 : _GEN10685;
wire  _GEN10691 = io_x[33] ? _GEN10690 : _GEN10682;
wire  _GEN10692 = io_x[28] ? _GEN10691 : _GEN10676;
wire  _GEN10693 = io_x[18] ? _GEN10692 : _GEN10663;
wire  _GEN10694 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10695 = io_x[30] ? _GEN10694 : _GEN10239;
wire  _GEN10696 = io_x[26] ? _GEN10695 : _GEN10241;
wire  _GEN10697 = io_x[73] ? _GEN10259 : _GEN10696;
wire  _GEN10698 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10699 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10700 = io_x[30] ? _GEN10699 : _GEN10698;
wire  _GEN10701 = io_x[26] ? _GEN10700 : _GEN10246;
wire  _GEN10702 = io_x[73] ? _GEN10259 : _GEN10701;
wire  _GEN10703 = io_x[33] ? _GEN10702 : _GEN10697;
wire  _GEN10704 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10705 = io_x[73] ? _GEN10243 : _GEN10704;
wire  _GEN10706 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10707 = io_x[30] ? _GEN10706 : _GEN10239;
wire  _GEN10708 = io_x[26] ? _GEN10707 : _GEN10241;
wire  _GEN10709 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10710 = io_x[30] ? _GEN10709 : _GEN10238;
wire  _GEN10711 = io_x[26] ? _GEN10710 : _GEN10241;
wire  _GEN10712 = io_x[73] ? _GEN10711 : _GEN10708;
wire  _GEN10713 = io_x[33] ? _GEN10712 : _GEN10705;
wire  _GEN10714 = io_x[28] ? _GEN10713 : _GEN10703;
wire  _GEN10715 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN10716 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10717 = io_x[30] ? _GEN10239 : _GEN10716;
wire  _GEN10718 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10719 = io_x[30] ? _GEN10239 : _GEN10718;
wire  _GEN10720 = io_x[26] ? _GEN10719 : _GEN10717;
wire  _GEN10721 = io_x[73] ? _GEN10720 : _GEN10715;
wire  _GEN10722 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10723 = io_x[30] ? _GEN10239 : _GEN10722;
wire  _GEN10724 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10725 = io_x[30] ? _GEN10724 : _GEN10239;
wire  _GEN10726 = io_x[26] ? _GEN10725 : _GEN10723;
wire  _GEN10727 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10728 = io_x[30] ? _GEN10727 : _GEN10238;
wire  _GEN10729 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10730 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10731 = io_x[30] ? _GEN10730 : _GEN10729;
wire  _GEN10732 = io_x[26] ? _GEN10731 : _GEN10728;
wire  _GEN10733 = io_x[73] ? _GEN10732 : _GEN10726;
wire  _GEN10734 = io_x[33] ? _GEN10733 : _GEN10721;
wire  _GEN10735 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10736 = io_x[30] ? _GEN10735 : _GEN10239;
wire  _GEN10737 = io_x[26] ? _GEN10736 : _GEN10241;
wire  _GEN10738 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10739 = io_x[26] ? _GEN10738 : _GEN10241;
wire  _GEN10740 = io_x[73] ? _GEN10739 : _GEN10737;
wire  _GEN10741 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10742 = io_x[30] ? _GEN10741 : _GEN10238;
wire  _GEN10743 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10744 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10745 = io_x[30] ? _GEN10744 : _GEN10743;
wire  _GEN10746 = io_x[26] ? _GEN10745 : _GEN10742;
wire  _GEN10747 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10748 = io_x[30] ? _GEN10747 : _GEN10239;
wire  _GEN10749 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10750 = io_x[30] ? _GEN10749 : _GEN10239;
wire  _GEN10751 = io_x[26] ? _GEN10750 : _GEN10748;
wire  _GEN10752 = io_x[73] ? _GEN10751 : _GEN10746;
wire  _GEN10753 = io_x[33] ? _GEN10752 : _GEN10740;
wire  _GEN10754 = io_x[28] ? _GEN10753 : _GEN10734;
wire  _GEN10755 = io_x[18] ? _GEN10754 : _GEN10714;
wire  _GEN10756 = io_x[25] ? _GEN10755 : _GEN10693;
wire  _GEN10757 = io_x[29] ? _GEN10756 : _GEN10646;
wire  _GEN10758 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10759 = io_x[30] ? _GEN10758 : _GEN10239;
wire  _GEN10760 = io_x[26] ? _GEN10759 : _GEN10241;
wire  _GEN10761 = io_x[73] ? _GEN10243 : _GEN10760;
wire  _GEN10762 = io_x[33] ? _GEN10761 : _GEN10237;
wire  _GEN10763 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10764 = io_x[73] ? _GEN10763 : _GEN10243;
wire  _GEN10765 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10766 = io_x[30] ? _GEN10765 : _GEN10238;
wire  _GEN10767 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10768 = io_x[30] ? _GEN10239 : _GEN10767;
wire  _GEN10769 = io_x[26] ? _GEN10768 : _GEN10766;
wire  _GEN10770 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10771 = io_x[73] ? _GEN10770 : _GEN10769;
wire  _GEN10772 = io_x[33] ? _GEN10771 : _GEN10764;
wire  _GEN10773 = io_x[28] ? _GEN10772 : _GEN10762;
wire  _GEN10774 = io_x[73] ? _GEN10259 : _GEN10243;
wire  _GEN10775 = io_x[33] ? _GEN10774 : _GEN10237;
wire  _GEN10776 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10777 = io_x[30] ? _GEN10776 : _GEN10238;
wire  _GEN10778 = io_x[26] ? _GEN10777 : _GEN10241;
wire  _GEN10779 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10780 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10781 = io_x[30] ? _GEN10780 : _GEN10779;
wire  _GEN10782 = io_x[26] ? _GEN10781 : _GEN10246;
wire  _GEN10783 = io_x[73] ? _GEN10782 : _GEN10778;
wire  _GEN10784 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10785 = io_x[30] ? _GEN10784 : _GEN10238;
wire  _GEN10786 = io_x[26] ? _GEN10785 : _GEN10241;
wire  _GEN10787 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10788 = io_x[30] ? _GEN10239 : _GEN10787;
wire  _GEN10789 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10790 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10791 = io_x[30] ? _GEN10790 : _GEN10789;
wire  _GEN10792 = io_x[26] ? _GEN10791 : _GEN10788;
wire  _GEN10793 = io_x[73] ? _GEN10792 : _GEN10786;
wire  _GEN10794 = io_x[33] ? _GEN10793 : _GEN10783;
wire  _GEN10795 = io_x[28] ? _GEN10794 : _GEN10775;
wire  _GEN10796 = io_x[18] ? _GEN10795 : _GEN10773;
wire  _GEN10797 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10798 = io_x[73] ? _GEN10243 : _GEN10797;
wire  _GEN10799 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10800 = io_x[26] ? _GEN10799 : _GEN10246;
wire  _GEN10801 = io_x[73] ? _GEN10243 : _GEN10800;
wire  _GEN10802 = io_x[33] ? _GEN10801 : _GEN10798;
wire  _GEN10803 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN10804 = io_x[73] ? _GEN10243 : _GEN10803;
wire  _GEN10805 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10806 = io_x[30] ? _GEN10805 : _GEN10239;
wire  _GEN10807 = io_x[26] ? _GEN10806 : _GEN10241;
wire  _GEN10808 = io_x[73] ? _GEN10243 : _GEN10807;
wire  _GEN10809 = io_x[33] ? _GEN10808 : _GEN10804;
wire  _GEN10810 = io_x[28] ? _GEN10809 : _GEN10802;
wire  _GEN10811 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10812 = io_x[30] ? _GEN10238 : _GEN10811;
wire  _GEN10813 = io_x[26] ? _GEN10246 : _GEN10812;
wire  _GEN10814 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10815 = io_x[30] ? _GEN10814 : _GEN10239;
wire  _GEN10816 = io_x[26] ? _GEN10815 : _GEN10246;
wire  _GEN10817 = io_x[73] ? _GEN10816 : _GEN10813;
wire  _GEN10818 = io_x[33] ? _GEN10817 : _GEN10306;
wire  _GEN10819 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10820 = io_x[30] ? _GEN10819 : _GEN10239;
wire  _GEN10821 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10822 = io_x[30] ? _GEN10821 : _GEN10239;
wire  _GEN10823 = io_x[26] ? _GEN10822 : _GEN10820;
wire  _GEN10824 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10825 = io_x[30] ? _GEN10824 : _GEN10239;
wire  _GEN10826 = io_x[26] ? _GEN10825 : _GEN10241;
wire  _GEN10827 = io_x[73] ? _GEN10826 : _GEN10823;
wire  _GEN10828 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10829 = io_x[30] ? _GEN10828 : _GEN10239;
wire  _GEN10830 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10831 = io_x[30] ? _GEN10830 : _GEN10239;
wire  _GEN10832 = io_x[26] ? _GEN10831 : _GEN10829;
wire  _GEN10833 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10834 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10835 = io_x[30] ? _GEN10834 : _GEN10833;
wire  _GEN10836 = io_x[26] ? _GEN10835 : _GEN10241;
wire  _GEN10837 = io_x[73] ? _GEN10836 : _GEN10832;
wire  _GEN10838 = io_x[33] ? _GEN10837 : _GEN10827;
wire  _GEN10839 = io_x[28] ? _GEN10838 : _GEN10818;
wire  _GEN10840 = io_x[18] ? _GEN10839 : _GEN10810;
wire  _GEN10841 = io_x[25] ? _GEN10840 : _GEN10796;
wire  _GEN10842 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10843 = io_x[30] ? _GEN10842 : _GEN10239;
wire  _GEN10844 = io_x[26] ? _GEN10246 : _GEN10843;
wire  _GEN10845 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10846 = io_x[26] ? _GEN10241 : _GEN10845;
wire  _GEN10847 = io_x[73] ? _GEN10846 : _GEN10844;
wire  _GEN10848 = io_x[33] ? _GEN10847 : _GEN10237;
wire  _GEN10849 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10850 = io_x[73] ? _GEN10243 : _GEN10849;
wire  _GEN10851 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10852 = io_x[30] ? _GEN10851 : _GEN10239;
wire  _GEN10853 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10854 = io_x[30] ? _GEN10853 : _GEN10238;
wire  _GEN10855 = io_x[26] ? _GEN10854 : _GEN10852;
wire  _GEN10856 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN10857 = io_x[73] ? _GEN10856 : _GEN10855;
wire  _GEN10858 = io_x[33] ? _GEN10857 : _GEN10850;
wire  _GEN10859 = io_x[28] ? _GEN10858 : _GEN10848;
wire  _GEN10860 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10861 = io_x[30] ? _GEN10239 : _GEN10860;
wire  _GEN10862 = io_x[26] ? _GEN10861 : _GEN10241;
wire  _GEN10863 = io_x[73] ? _GEN10243 : _GEN10862;
wire  _GEN10864 = io_x[73] ? _GEN10243 : _GEN10259;
wire  _GEN10865 = io_x[33] ? _GEN10864 : _GEN10863;
wire  _GEN10866 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10867 = io_x[30] ? _GEN10238 : _GEN10866;
wire  _GEN10868 = io_x[26] ? _GEN10867 : _GEN10241;
wire  _GEN10869 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10870 = io_x[26] ? _GEN10869 : _GEN10241;
wire  _GEN10871 = io_x[73] ? _GEN10870 : _GEN10868;
wire  _GEN10872 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10873 = io_x[26] ? _GEN10872 : _GEN10241;
wire  _GEN10874 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10875 = io_x[26] ? _GEN10874 : _GEN10241;
wire  _GEN10876 = io_x[73] ? _GEN10875 : _GEN10873;
wire  _GEN10877 = io_x[33] ? _GEN10876 : _GEN10871;
wire  _GEN10878 = io_x[28] ? _GEN10877 : _GEN10865;
wire  _GEN10879 = io_x[18] ? _GEN10878 : _GEN10859;
wire  _GEN10880 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10881 = io_x[30] ? _GEN10239 : _GEN10880;
wire  _GEN10882 = io_x[26] ? _GEN10241 : _GEN10881;
wire  _GEN10883 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN10884 = io_x[73] ? _GEN10883 : _GEN10882;
wire  _GEN10885 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10886 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10887 = io_x[30] ? _GEN10886 : _GEN10885;
wire  _GEN10888 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10889 = io_x[30] ? _GEN10888 : _GEN10238;
wire  _GEN10890 = io_x[26] ? _GEN10889 : _GEN10887;
wire  _GEN10891 = io_x[73] ? _GEN10243 : _GEN10890;
wire  _GEN10892 = io_x[33] ? _GEN10891 : _GEN10884;
wire  _GEN10893 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10894 = io_x[30] ? _GEN10893 : _GEN10238;
wire  _GEN10895 = io_x[26] ? _GEN10894 : _GEN10241;
wire  _GEN10896 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10897 = io_x[26] ? _GEN10896 : _GEN10246;
wire  _GEN10898 = io_x[73] ? _GEN10897 : _GEN10895;
wire  _GEN10899 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10900 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10901 = io_x[30] ? _GEN10900 : _GEN10899;
wire  _GEN10902 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10903 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10904 = io_x[30] ? _GEN10903 : _GEN10902;
wire  _GEN10905 = io_x[26] ? _GEN10904 : _GEN10901;
wire  _GEN10906 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10907 = io_x[30] ? _GEN10906 : _GEN10239;
wire  _GEN10908 = io_x[26] ? _GEN10907 : _GEN10246;
wire  _GEN10909 = io_x[73] ? _GEN10908 : _GEN10905;
wire  _GEN10910 = io_x[33] ? _GEN10909 : _GEN10898;
wire  _GEN10911 = io_x[28] ? _GEN10910 : _GEN10892;
wire  _GEN10912 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10913 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10914 = io_x[30] ? _GEN10913 : _GEN10912;
wire  _GEN10915 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN10916 = io_x[26] ? _GEN10915 : _GEN10914;
wire  _GEN10917 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10918 = io_x[30] ? _GEN10239 : _GEN10917;
wire  _GEN10919 = io_x[26] ? _GEN10241 : _GEN10918;
wire  _GEN10920 = io_x[73] ? _GEN10919 : _GEN10916;
wire  _GEN10921 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10922 = io_x[30] ? _GEN10921 : _GEN10239;
wire  _GEN10923 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10924 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10925 = io_x[30] ? _GEN10924 : _GEN10923;
wire  _GEN10926 = io_x[26] ? _GEN10925 : _GEN10922;
wire  _GEN10927 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10928 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10929 = io_x[30] ? _GEN10928 : _GEN10927;
wire  _GEN10930 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10931 = io_x[30] ? _GEN10238 : _GEN10930;
wire  _GEN10932 = io_x[26] ? _GEN10931 : _GEN10929;
wire  _GEN10933 = io_x[73] ? _GEN10932 : _GEN10926;
wire  _GEN10934 = io_x[33] ? _GEN10933 : _GEN10920;
wire  _GEN10935 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10936 = io_x[30] ? _GEN10239 : _GEN10935;
wire  _GEN10937 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10938 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10939 = io_x[30] ? _GEN10938 : _GEN10937;
wire  _GEN10940 = io_x[26] ? _GEN10939 : _GEN10936;
wire  _GEN10941 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10942 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10943 = io_x[30] ? _GEN10942 : _GEN10941;
wire  _GEN10944 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10945 = io_x[30] ? _GEN10944 : _GEN10239;
wire  _GEN10946 = io_x[26] ? _GEN10945 : _GEN10943;
wire  _GEN10947 = io_x[73] ? _GEN10946 : _GEN10940;
wire  _GEN10948 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10949 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10950 = io_x[30] ? _GEN10949 : _GEN10948;
wire  _GEN10951 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10952 = io_x[30] ? _GEN10951 : _GEN10239;
wire  _GEN10953 = io_x[26] ? _GEN10952 : _GEN10950;
wire  _GEN10954 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10955 = io_x[30] ? _GEN10239 : _GEN10954;
wire  _GEN10956 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10957 = io_x[30] ? _GEN10956 : _GEN10239;
wire  _GEN10958 = io_x[26] ? _GEN10957 : _GEN10955;
wire  _GEN10959 = io_x[73] ? _GEN10958 : _GEN10953;
wire  _GEN10960 = io_x[33] ? _GEN10959 : _GEN10947;
wire  _GEN10961 = io_x[28] ? _GEN10960 : _GEN10934;
wire  _GEN10962 = io_x[18] ? _GEN10961 : _GEN10911;
wire  _GEN10963 = io_x[25] ? _GEN10962 : _GEN10879;
wire  _GEN10964 = io_x[29] ? _GEN10963 : _GEN10841;
wire  _GEN10965 = io_x[23] ? _GEN10964 : _GEN10757;
wire  _GEN10966 = io_x[31] ? _GEN10965 : _GEN10564;
wire  _GEN10967 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10968 = io_x[30] ? _GEN10967 : _GEN10239;
wire  _GEN10969 = io_x[26] ? _GEN10968 : _GEN10241;
wire  _GEN10970 = io_x[73] ? _GEN10243 : _GEN10969;
wire  _GEN10971 = io_x[33] ? _GEN10970 : _GEN10237;
wire  _GEN10972 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN10973 = io_x[73] ? _GEN10972 : _GEN10243;
wire  _GEN10974 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN10975 = io_x[26] ? _GEN10974 : _GEN10241;
wire  _GEN10976 = io_x[73] ? _GEN10259 : _GEN10975;
wire  _GEN10977 = io_x[33] ? _GEN10976 : _GEN10973;
wire  _GEN10978 = io_x[28] ? _GEN10977 : _GEN10971;
wire  _GEN10979 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10980 = io_x[30] ? _GEN10979 : _GEN10239;
wire  _GEN10981 = io_x[26] ? _GEN10980 : _GEN10241;
wire  _GEN10982 = io_x[73] ? _GEN10981 : _GEN10243;
wire  _GEN10983 = io_x[33] ? _GEN10982 : _GEN10306;
wire  _GEN10984 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10985 = io_x[30] ? _GEN10984 : _GEN10239;
wire  _GEN10986 = io_x[26] ? _GEN10985 : _GEN10241;
wire  _GEN10987 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN10988 = io_x[73] ? _GEN10987 : _GEN10986;
wire  _GEN10989 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10990 = io_x[30] ? _GEN10989 : _GEN10239;
wire  _GEN10991 = io_x[26] ? _GEN10246 : _GEN10990;
wire  _GEN10992 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN10993 = io_x[30] ? _GEN10992 : _GEN10239;
wire  _GEN10994 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN10995 = io_x[30] ? _GEN10994 : _GEN10238;
wire  _GEN10996 = io_x[26] ? _GEN10995 : _GEN10993;
wire  _GEN10997 = io_x[73] ? _GEN10996 : _GEN10991;
wire  _GEN10998 = io_x[33] ? _GEN10997 : _GEN10988;
wire  _GEN10999 = io_x[28] ? _GEN10998 : _GEN10983;
wire  _GEN11000 = io_x[18] ? _GEN10999 : _GEN10978;
wire  _GEN11001 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN11002 = io_x[73] ? _GEN11001 : _GEN10243;
wire  _GEN11003 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11004 = io_x[26] ? _GEN11003 : _GEN10241;
wire  _GEN11005 = io_x[73] ? _GEN10243 : _GEN11004;
wire  _GEN11006 = io_x[33] ? _GEN11005 : _GEN11002;
wire  _GEN11007 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11008 = io_x[26] ? _GEN11007 : _GEN10241;
wire  _GEN11009 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11010 = io_x[30] ? _GEN11009 : _GEN10239;
wire  _GEN11011 = io_x[26] ? _GEN10241 : _GEN11010;
wire  _GEN11012 = io_x[73] ? _GEN11011 : _GEN11008;
wire  _GEN11013 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11014 = io_x[30] ? _GEN11013 : _GEN10239;
wire  _GEN11015 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11016 = io_x[30] ? _GEN11015 : _GEN10238;
wire  _GEN11017 = io_x[26] ? _GEN11016 : _GEN11014;
wire  _GEN11018 = io_x[73] ? _GEN10243 : _GEN11017;
wire  _GEN11019 = io_x[33] ? _GEN11018 : _GEN11012;
wire  _GEN11020 = io_x[28] ? _GEN11019 : _GEN11006;
wire  _GEN11021 = 1'b0;
wire  _GEN11022 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11023 = io_x[30] ? _GEN11022 : _GEN10239;
wire  _GEN11024 = io_x[26] ? _GEN11023 : _GEN10246;
wire  _GEN11025 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11026 = io_x[26] ? _GEN11025 : _GEN10241;
wire  _GEN11027 = io_x[73] ? _GEN11026 : _GEN11024;
wire  _GEN11028 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11029 = io_x[30] ? _GEN11028 : _GEN10239;
wire  _GEN11030 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11031 = io_x[30] ? _GEN11030 : _GEN10239;
wire  _GEN11032 = io_x[26] ? _GEN11031 : _GEN11029;
wire  _GEN11033 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11034 = io_x[26] ? _GEN10241 : _GEN11033;
wire  _GEN11035 = io_x[73] ? _GEN11034 : _GEN11032;
wire  _GEN11036 = io_x[33] ? _GEN11035 : _GEN11027;
wire  _GEN11037 = io_x[28] ? _GEN11036 : _GEN11021;
wire  _GEN11038 = io_x[18] ? _GEN11037 : _GEN11020;
wire  _GEN11039 = io_x[25] ? _GEN11038 : _GEN11000;
wire  _GEN11040 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11041 = io_x[30] ? _GEN10239 : _GEN11040;
wire  _GEN11042 = io_x[26] ? _GEN11041 : _GEN10241;
wire  _GEN11043 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN11044 = io_x[73] ? _GEN11043 : _GEN11042;
wire  _GEN11045 = io_x[33] ? _GEN11044 : _GEN10237;
wire  _GEN11046 = io_x[73] ? _GEN10243 : _GEN10259;
wire  _GEN11047 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11048 = io_x[30] ? _GEN11047 : _GEN10239;
wire  _GEN11049 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11050 = io_x[26] ? _GEN11049 : _GEN11048;
wire  _GEN11051 = io_x[73] ? _GEN10259 : _GEN11050;
wire  _GEN11052 = io_x[33] ? _GEN11051 : _GEN11046;
wire  _GEN11053 = io_x[28] ? _GEN11052 : _GEN11045;
wire  _GEN11054 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11055 = io_x[26] ? _GEN11054 : _GEN10241;
wire  _GEN11056 = io_x[73] ? _GEN11055 : _GEN10259;
wire  _GEN11057 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11058 = io_x[30] ? _GEN11057 : _GEN10239;
wire  _GEN11059 = io_x[26] ? _GEN11058 : _GEN10246;
wire  _GEN11060 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11061 = io_x[30] ? _GEN10238 : _GEN11060;
wire  _GEN11062 = io_x[26] ? _GEN11061 : _GEN10241;
wire  _GEN11063 = io_x[73] ? _GEN11062 : _GEN11059;
wire  _GEN11064 = io_x[33] ? _GEN11063 : _GEN11056;
wire  _GEN11065 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11066 = io_x[26] ? _GEN11065 : _GEN10241;
wire  _GEN11067 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11068 = io_x[26] ? _GEN11067 : _GEN10241;
wire  _GEN11069 = io_x[73] ? _GEN11068 : _GEN11066;
wire  _GEN11070 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11071 = io_x[26] ? _GEN10246 : _GEN11070;
wire  _GEN11072 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11073 = io_x[26] ? _GEN11072 : _GEN10241;
wire  _GEN11074 = io_x[73] ? _GEN11073 : _GEN11071;
wire  _GEN11075 = io_x[33] ? _GEN11074 : _GEN11069;
wire  _GEN11076 = io_x[28] ? _GEN11075 : _GEN11064;
wire  _GEN11077 = io_x[18] ? _GEN11076 : _GEN11053;
wire  _GEN11078 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11079 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11080 = io_x[26] ? _GEN11079 : _GEN11078;
wire  _GEN11081 = io_x[73] ? _GEN11080 : _GEN10259;
wire  _GEN11082 = io_x[33] ? _GEN11081 : _GEN10306;
wire  _GEN11083 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11084 = io_x[26] ? _GEN11083 : _GEN10241;
wire  _GEN11085 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11086 = io_x[30] ? _GEN10238 : _GEN11085;
wire  _GEN11087 = io_x[26] ? _GEN11086 : _GEN10246;
wire  _GEN11088 = io_x[73] ? _GEN11087 : _GEN11084;
wire  _GEN11089 = io_x[33] ? _GEN11088 : _GEN10237;
wire  _GEN11090 = io_x[28] ? _GEN11089 : _GEN11082;
wire  _GEN11091 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11092 = io_x[26] ? _GEN10241 : _GEN11091;
wire  _GEN11093 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11094 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11095 = io_x[26] ? _GEN11094 : _GEN11093;
wire  _GEN11096 = io_x[73] ? _GEN11095 : _GEN11092;
wire  _GEN11097 = io_x[33] ? _GEN11096 : _GEN10237;
wire  _GEN11098 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11099 = io_x[30] ? _GEN11098 : _GEN10239;
wire  _GEN11100 = io_x[26] ? _GEN11099 : _GEN10241;
wire  _GEN11101 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11102 = io_x[30] ? _GEN10239 : _GEN11101;
wire  _GEN11103 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11104 = io_x[30] ? _GEN11103 : _GEN10239;
wire  _GEN11105 = io_x[26] ? _GEN11104 : _GEN11102;
wire  _GEN11106 = io_x[73] ? _GEN11105 : _GEN11100;
wire  _GEN11107 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11108 = io_x[30] ? _GEN11107 : _GEN10239;
wire  _GEN11109 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11110 = io_x[30] ? _GEN11109 : _GEN10238;
wire  _GEN11111 = io_x[26] ? _GEN11110 : _GEN11108;
wire  _GEN11112 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11113 = io_x[30] ? _GEN11112 : _GEN10239;
wire  _GEN11114 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11115 = io_x[30] ? _GEN11114 : _GEN10239;
wire  _GEN11116 = io_x[26] ? _GEN11115 : _GEN11113;
wire  _GEN11117 = io_x[73] ? _GEN11116 : _GEN11111;
wire  _GEN11118 = io_x[33] ? _GEN11117 : _GEN11106;
wire  _GEN11119 = io_x[28] ? _GEN11118 : _GEN11097;
wire  _GEN11120 = io_x[18] ? _GEN11119 : _GEN11090;
wire  _GEN11121 = io_x[25] ? _GEN11120 : _GEN11077;
wire  _GEN11122 = io_x[29] ? _GEN11121 : _GEN11039;
wire  _GEN11123 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN11124 = io_x[73] ? _GEN11123 : _GEN10243;
wire  _GEN11125 = io_x[33] ? _GEN11124 : _GEN10237;
wire  _GEN11126 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN11127 = io_x[73] ? _GEN10259 : _GEN11126;
wire  _GEN11128 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11129 = io_x[30] ? _GEN11128 : _GEN10239;
wire  _GEN11130 = io_x[26] ? _GEN11129 : _GEN10241;
wire  _GEN11131 = io_x[73] ? _GEN10243 : _GEN11130;
wire  _GEN11132 = io_x[33] ? _GEN11131 : _GEN11127;
wire  _GEN11133 = io_x[28] ? _GEN11132 : _GEN11125;
wire  _GEN11134 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN11135 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11136 = io_x[30] ? _GEN11135 : _GEN10239;
wire  _GEN11137 = io_x[26] ? _GEN10246 : _GEN11136;
wire  _GEN11138 = io_x[73] ? _GEN11137 : _GEN11134;
wire  _GEN11139 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11140 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11141 = io_x[30] ? _GEN11140 : _GEN10239;
wire  _GEN11142 = io_x[26] ? _GEN11141 : _GEN11139;
wire  _GEN11143 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11144 = io_x[30] ? _GEN11143 : _GEN10239;
wire  _GEN11145 = io_x[26] ? _GEN11144 : _GEN10241;
wire  _GEN11146 = io_x[73] ? _GEN11145 : _GEN11142;
wire  _GEN11147 = io_x[33] ? _GEN11146 : _GEN11138;
wire  _GEN11148 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11149 = io_x[26] ? _GEN11148 : _GEN10246;
wire  _GEN11150 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11151 = io_x[30] ? _GEN11150 : _GEN10239;
wire  _GEN11152 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11153 = io_x[30] ? _GEN11152 : _GEN10239;
wire  _GEN11154 = io_x[26] ? _GEN11153 : _GEN11151;
wire  _GEN11155 = io_x[73] ? _GEN11154 : _GEN11149;
wire  _GEN11156 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11157 = io_x[30] ? _GEN10239 : _GEN11156;
wire  _GEN11158 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11159 = io_x[30] ? _GEN11158 : _GEN10239;
wire  _GEN11160 = io_x[26] ? _GEN11159 : _GEN11157;
wire  _GEN11161 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11162 = io_x[30] ? _GEN10238 : _GEN11161;
wire  _GEN11163 = io_x[26] ? _GEN11162 : _GEN10241;
wire  _GEN11164 = io_x[73] ? _GEN11163 : _GEN11160;
wire  _GEN11165 = io_x[33] ? _GEN11164 : _GEN11155;
wire  _GEN11166 = io_x[28] ? _GEN11165 : _GEN11147;
wire  _GEN11167 = io_x[18] ? _GEN11166 : _GEN11133;
wire  _GEN11168 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11169 = io_x[30] ? _GEN10239 : _GEN11168;
wire  _GEN11170 = io_x[26] ? _GEN10241 : _GEN11169;
wire  _GEN11171 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11172 = io_x[30] ? _GEN11171 : _GEN10239;
wire  _GEN11173 = io_x[26] ? _GEN10241 : _GEN11172;
wire  _GEN11174 = io_x[73] ? _GEN11173 : _GEN11170;
wire  _GEN11175 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN11176 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11177 = io_x[30] ? _GEN11176 : _GEN10239;
wire  _GEN11178 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11179 = io_x[30] ? _GEN11178 : _GEN10239;
wire  _GEN11180 = io_x[26] ? _GEN11179 : _GEN11177;
wire  _GEN11181 = io_x[73] ? _GEN11180 : _GEN11175;
wire  _GEN11182 = io_x[33] ? _GEN11181 : _GEN11174;
wire  _GEN11183 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11184 = io_x[30] ? _GEN11183 : _GEN10238;
wire  _GEN11185 = io_x[26] ? _GEN11184 : _GEN10246;
wire  _GEN11186 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11187 = io_x[26] ? _GEN11186 : _GEN10246;
wire  _GEN11188 = io_x[73] ? _GEN11187 : _GEN11185;
wire  _GEN11189 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11190 = io_x[30] ? _GEN11189 : _GEN10238;
wire  _GEN11191 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11192 = io_x[30] ? _GEN11191 : _GEN10238;
wire  _GEN11193 = io_x[26] ? _GEN11192 : _GEN11190;
wire  _GEN11194 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11195 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11196 = io_x[26] ? _GEN11195 : _GEN11194;
wire  _GEN11197 = io_x[73] ? _GEN11196 : _GEN11193;
wire  _GEN11198 = io_x[33] ? _GEN11197 : _GEN11188;
wire  _GEN11199 = io_x[28] ? _GEN11198 : _GEN11182;
wire  _GEN11200 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11201 = io_x[30] ? _GEN11200 : _GEN10239;
wire  _GEN11202 = io_x[26] ? _GEN11201 : _GEN10241;
wire  _GEN11203 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11204 = io_x[30] ? _GEN11203 : _GEN10239;
wire  _GEN11205 = io_x[26] ? _GEN11204 : _GEN10241;
wire  _GEN11206 = io_x[73] ? _GEN11205 : _GEN11202;
wire  _GEN11207 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11208 = io_x[26] ? _GEN11207 : _GEN10241;
wire  _GEN11209 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11210 = io_x[30] ? _GEN11209 : _GEN10238;
wire  _GEN11211 = io_x[26] ? _GEN10246 : _GEN11210;
wire  _GEN11212 = io_x[73] ? _GEN11211 : _GEN11208;
wire  _GEN11213 = io_x[33] ? _GEN11212 : _GEN11206;
wire  _GEN11214 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11215 = io_x[30] ? _GEN11214 : _GEN10239;
wire  _GEN11216 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11217 = io_x[26] ? _GEN11216 : _GEN11215;
wire  _GEN11218 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11219 = io_x[30] ? _GEN10238 : _GEN11218;
wire  _GEN11220 = io_x[26] ? _GEN11219 : _GEN10241;
wire  _GEN11221 = io_x[73] ? _GEN11220 : _GEN11217;
wire  _GEN11222 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11223 = io_x[30] ? _GEN11222 : _GEN10238;
wire  _GEN11224 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11225 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11226 = io_x[30] ? _GEN11225 : _GEN11224;
wire  _GEN11227 = io_x[26] ? _GEN11226 : _GEN11223;
wire  _GEN11228 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11229 = io_x[30] ? _GEN10238 : _GEN11228;
wire  _GEN11230 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11231 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11232 = io_x[30] ? _GEN11231 : _GEN11230;
wire  _GEN11233 = io_x[26] ? _GEN11232 : _GEN11229;
wire  _GEN11234 = io_x[73] ? _GEN11233 : _GEN11227;
wire  _GEN11235 = io_x[33] ? _GEN11234 : _GEN11221;
wire  _GEN11236 = io_x[28] ? _GEN11235 : _GEN11213;
wire  _GEN11237 = io_x[18] ? _GEN11236 : _GEN11199;
wire  _GEN11238 = io_x[25] ? _GEN11237 : _GEN11167;
wire  _GEN11239 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11240 = io_x[30] ? _GEN10238 : _GEN11239;
wire  _GEN11241 = io_x[26] ? _GEN11240 : _GEN10241;
wire  _GEN11242 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11243 = io_x[26] ? _GEN10241 : _GEN11242;
wire  _GEN11244 = io_x[73] ? _GEN11243 : _GEN11241;
wire  _GEN11245 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11246 = io_x[30] ? _GEN11245 : _GEN10239;
wire  _GEN11247 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11248 = io_x[30] ? _GEN10239 : _GEN11247;
wire  _GEN11249 = io_x[26] ? _GEN11248 : _GEN11246;
wire  _GEN11250 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11251 = io_x[26] ? _GEN11250 : _GEN10246;
wire  _GEN11252 = io_x[73] ? _GEN11251 : _GEN11249;
wire  _GEN11253 = io_x[33] ? _GEN11252 : _GEN11244;
wire  _GEN11254 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11255 = io_x[26] ? _GEN11254 : _GEN10241;
wire  _GEN11256 = io_x[73] ? _GEN10243 : _GEN11255;
wire  _GEN11257 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11258 = io_x[30] ? _GEN11257 : _GEN10238;
wire  _GEN11259 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11260 = io_x[30] ? _GEN11259 : _GEN10239;
wire  _GEN11261 = io_x[26] ? _GEN11260 : _GEN11258;
wire  _GEN11262 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11263 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11264 = io_x[26] ? _GEN11263 : _GEN11262;
wire  _GEN11265 = io_x[73] ? _GEN11264 : _GEN11261;
wire  _GEN11266 = io_x[33] ? _GEN11265 : _GEN11256;
wire  _GEN11267 = io_x[28] ? _GEN11266 : _GEN11253;
wire  _GEN11268 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11269 = io_x[26] ? _GEN10241 : _GEN11268;
wire  _GEN11270 = io_x[73] ? _GEN11269 : _GEN10259;
wire  _GEN11271 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11272 = io_x[30] ? _GEN11271 : _GEN10239;
wire  _GEN11273 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11274 = io_x[26] ? _GEN11273 : _GEN11272;
wire  _GEN11275 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11276 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11277 = io_x[26] ? _GEN11276 : _GEN11275;
wire  _GEN11278 = io_x[73] ? _GEN11277 : _GEN11274;
wire  _GEN11279 = io_x[33] ? _GEN11278 : _GEN11270;
wire  _GEN11280 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11281 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11282 = io_x[30] ? _GEN11281 : _GEN11280;
wire  _GEN11283 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11284 = io_x[26] ? _GEN11283 : _GEN11282;
wire  _GEN11285 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN11286 = io_x[73] ? _GEN11285 : _GEN11284;
wire  _GEN11287 = io_x[33] ? _GEN11286 : _GEN10306;
wire  _GEN11288 = io_x[28] ? _GEN11287 : _GEN11279;
wire  _GEN11289 = io_x[18] ? _GEN11288 : _GEN11267;
wire  _GEN11290 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11291 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11292 = io_x[30] ? _GEN11291 : _GEN11290;
wire  _GEN11293 = io_x[26] ? _GEN10241 : _GEN11292;
wire  _GEN11294 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11295 = io_x[30] ? _GEN11294 : _GEN10239;
wire  _GEN11296 = io_x[26] ? _GEN11295 : _GEN10246;
wire  _GEN11297 = io_x[73] ? _GEN11296 : _GEN11293;
wire  _GEN11298 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11299 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11300 = io_x[30] ? _GEN11299 : _GEN11298;
wire  _GEN11301 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11302 = io_x[30] ? _GEN11301 : _GEN10239;
wire  _GEN11303 = io_x[26] ? _GEN11302 : _GEN11300;
wire  _GEN11304 = io_x[73] ? _GEN10259 : _GEN11303;
wire  _GEN11305 = io_x[33] ? _GEN11304 : _GEN11297;
wire  _GEN11306 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11307 = io_x[30] ? _GEN11306 : _GEN10239;
wire  _GEN11308 = io_x[26] ? _GEN11307 : _GEN10246;
wire  _GEN11309 = io_x[73] ? _GEN10243 : _GEN11308;
wire  _GEN11310 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11311 = io_x[30] ? _GEN11310 : _GEN10238;
wire  _GEN11312 = io_x[26] ? _GEN11311 : _GEN10246;
wire  _GEN11313 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11314 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11315 = io_x[30] ? _GEN11314 : _GEN11313;
wire  _GEN11316 = io_x[26] ? _GEN11315 : _GEN10241;
wire  _GEN11317 = io_x[73] ? _GEN11316 : _GEN11312;
wire  _GEN11318 = io_x[33] ? _GEN11317 : _GEN11309;
wire  _GEN11319 = io_x[28] ? _GEN11318 : _GEN11305;
wire  _GEN11320 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11321 = io_x[26] ? _GEN11320 : _GEN10241;
wire  _GEN11322 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11323 = io_x[30] ? _GEN10239 : _GEN11322;
wire  _GEN11324 = io_x[26] ? _GEN10241 : _GEN11323;
wire  _GEN11325 = io_x[73] ? _GEN11324 : _GEN11321;
wire  _GEN11326 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11327 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11328 = io_x[26] ? _GEN11327 : _GEN11326;
wire  _GEN11329 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11330 = io_x[26] ? _GEN11329 : _GEN10241;
wire  _GEN11331 = io_x[73] ? _GEN11330 : _GEN11328;
wire  _GEN11332 = io_x[33] ? _GEN11331 : _GEN11325;
wire  _GEN11333 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11334 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11335 = io_x[30] ? _GEN11334 : _GEN10239;
wire  _GEN11336 = io_x[26] ? _GEN11335 : _GEN11333;
wire  _GEN11337 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11338 = io_x[30] ? _GEN11337 : _GEN10238;
wire  _GEN11339 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11340 = io_x[30] ? _GEN11339 : _GEN10239;
wire  _GEN11341 = io_x[26] ? _GEN11340 : _GEN11338;
wire  _GEN11342 = io_x[73] ? _GEN11341 : _GEN11336;
wire  _GEN11343 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11344 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11345 = io_x[30] ? _GEN11344 : _GEN11343;
wire  _GEN11346 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11347 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11348 = io_x[30] ? _GEN11347 : _GEN11346;
wire  _GEN11349 = io_x[26] ? _GEN11348 : _GEN11345;
wire  _GEN11350 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11351 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11352 = io_x[30] ? _GEN11351 : _GEN11350;
wire  _GEN11353 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11354 = io_x[30] ? _GEN11353 : _GEN10239;
wire  _GEN11355 = io_x[26] ? _GEN11354 : _GEN11352;
wire  _GEN11356 = io_x[73] ? _GEN11355 : _GEN11349;
wire  _GEN11357 = io_x[33] ? _GEN11356 : _GEN11342;
wire  _GEN11358 = io_x[28] ? _GEN11357 : _GEN11332;
wire  _GEN11359 = io_x[18] ? _GEN11358 : _GEN11319;
wire  _GEN11360 = io_x[25] ? _GEN11359 : _GEN11289;
wire  _GEN11361 = io_x[29] ? _GEN11360 : _GEN11238;
wire  _GEN11362 = io_x[23] ? _GEN11361 : _GEN11122;
wire  _GEN11363 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11364 = io_x[26] ? _GEN11363 : _GEN10241;
wire  _GEN11365 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11366 = io_x[26] ? _GEN10241 : _GEN11365;
wire  _GEN11367 = io_x[73] ? _GEN11366 : _GEN11364;
wire  _GEN11368 = io_x[33] ? _GEN11367 : _GEN10237;
wire  _GEN11369 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11370 = io_x[26] ? _GEN11369 : _GEN10241;
wire  _GEN11371 = io_x[73] ? _GEN10243 : _GEN11370;
wire  _GEN11372 = io_x[33] ? _GEN11371 : _GEN10237;
wire  _GEN11373 = io_x[28] ? _GEN11372 : _GEN11368;
wire  _GEN11374 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11375 = io_x[26] ? _GEN11374 : _GEN10241;
wire  _GEN11376 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11377 = io_x[30] ? _GEN11376 : _GEN10239;
wire  _GEN11378 = io_x[26] ? _GEN10241 : _GEN11377;
wire  _GEN11379 = io_x[73] ? _GEN11378 : _GEN11375;
wire  _GEN11380 = io_x[33] ? _GEN11379 : _GEN10306;
wire  _GEN11381 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11382 = io_x[30] ? _GEN11381 : _GEN10239;
wire  _GEN11383 = io_x[26] ? _GEN11382 : _GEN10246;
wire  _GEN11384 = io_x[73] ? _GEN11383 : _GEN10259;
wire  _GEN11385 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11386 = io_x[30] ? _GEN10239 : _GEN11385;
wire  _GEN11387 = io_x[26] ? _GEN10246 : _GEN11386;
wire  _GEN11388 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11389 = io_x[30] ? _GEN11388 : _GEN10238;
wire  _GEN11390 = io_x[26] ? _GEN11389 : _GEN10241;
wire  _GEN11391 = io_x[73] ? _GEN11390 : _GEN11387;
wire  _GEN11392 = io_x[33] ? _GEN11391 : _GEN11384;
wire  _GEN11393 = io_x[28] ? _GEN11392 : _GEN11380;
wire  _GEN11394 = io_x[18] ? _GEN11393 : _GEN11373;
wire  _GEN11395 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11396 = io_x[26] ? _GEN10241 : _GEN11395;
wire  _GEN11397 = io_x[73] ? _GEN10243 : _GEN11396;
wire  _GEN11398 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11399 = io_x[30] ? _GEN11398 : _GEN10239;
wire  _GEN11400 = io_x[26] ? _GEN10241 : _GEN11399;
wire  _GEN11401 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11402 = io_x[26] ? _GEN10246 : _GEN11401;
wire  _GEN11403 = io_x[73] ? _GEN11402 : _GEN11400;
wire  _GEN11404 = io_x[33] ? _GEN11403 : _GEN11397;
wire  _GEN11405 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11406 = io_x[26] ? _GEN10241 : _GEN11405;
wire  _GEN11407 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11408 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11409 = io_x[30] ? _GEN11408 : _GEN10239;
wire  _GEN11410 = io_x[26] ? _GEN11409 : _GEN11407;
wire  _GEN11411 = io_x[73] ? _GEN11410 : _GEN11406;
wire  _GEN11412 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11413 = io_x[30] ? _GEN11412 : _GEN10239;
wire  _GEN11414 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11415 = io_x[30] ? _GEN11414 : _GEN10238;
wire  _GEN11416 = io_x[26] ? _GEN11415 : _GEN11413;
wire  _GEN11417 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11418 = io_x[30] ? _GEN10238 : _GEN11417;
wire  _GEN11419 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11420 = io_x[30] ? _GEN11419 : _GEN10239;
wire  _GEN11421 = io_x[26] ? _GEN11420 : _GEN11418;
wire  _GEN11422 = io_x[73] ? _GEN11421 : _GEN11416;
wire  _GEN11423 = io_x[33] ? _GEN11422 : _GEN11411;
wire  _GEN11424 = io_x[28] ? _GEN11423 : _GEN11404;
wire  _GEN11425 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN11426 = io_x[73] ? _GEN10243 : _GEN11425;
wire  _GEN11427 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11428 = io_x[26] ? _GEN10246 : _GEN11427;
wire  _GEN11429 = io_x[73] ? _GEN11428 : _GEN10243;
wire  _GEN11430 = io_x[33] ? _GEN11429 : _GEN11426;
wire  _GEN11431 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11432 = io_x[30] ? _GEN10239 : _GEN11431;
wire  _GEN11433 = io_x[26] ? _GEN10246 : _GEN11432;
wire  _GEN11434 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11435 = io_x[30] ? _GEN11434 : _GEN10239;
wire  _GEN11436 = io_x[26] ? _GEN11435 : _GEN10241;
wire  _GEN11437 = io_x[73] ? _GEN11436 : _GEN11433;
wire  _GEN11438 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11439 = io_x[26] ? _GEN11438 : _GEN10241;
wire  _GEN11440 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11441 = io_x[30] ? _GEN10239 : _GEN11440;
wire  _GEN11442 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11443 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11444 = io_x[30] ? _GEN11443 : _GEN11442;
wire  _GEN11445 = io_x[26] ? _GEN11444 : _GEN11441;
wire  _GEN11446 = io_x[73] ? _GEN11445 : _GEN11439;
wire  _GEN11447 = io_x[33] ? _GEN11446 : _GEN11437;
wire  _GEN11448 = io_x[28] ? _GEN11447 : _GEN11430;
wire  _GEN11449 = io_x[18] ? _GEN11448 : _GEN11424;
wire  _GEN11450 = io_x[25] ? _GEN11449 : _GEN11394;
wire  _GEN11451 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11452 = io_x[30] ? _GEN11451 : _GEN10238;
wire  _GEN11453 = io_x[26] ? _GEN11452 : _GEN10241;
wire  _GEN11454 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11455 = io_x[30] ? _GEN10239 : _GEN11454;
wire  _GEN11456 = io_x[26] ? _GEN11455 : _GEN10241;
wire  _GEN11457 = io_x[73] ? _GEN11456 : _GEN11453;
wire  _GEN11458 = io_x[33] ? _GEN11457 : _GEN10237;
wire  _GEN11459 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN11460 = io_x[73] ? _GEN10243 : _GEN11459;
wire  _GEN11461 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11462 = io_x[30] ? _GEN11461 : _GEN10238;
wire  _GEN11463 = io_x[26] ? _GEN11462 : _GEN10246;
wire  _GEN11464 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11465 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11466 = io_x[30] ? _GEN11465 : _GEN11464;
wire  _GEN11467 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11468 = io_x[26] ? _GEN11467 : _GEN11466;
wire  _GEN11469 = io_x[73] ? _GEN11468 : _GEN11463;
wire  _GEN11470 = io_x[33] ? _GEN11469 : _GEN11460;
wire  _GEN11471 = io_x[28] ? _GEN11470 : _GEN11458;
wire  _GEN11472 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11473 = io_x[26] ? _GEN11472 : _GEN10241;
wire  _GEN11474 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11475 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11476 = io_x[30] ? _GEN10238 : _GEN11475;
wire  _GEN11477 = io_x[26] ? _GEN11476 : _GEN11474;
wire  _GEN11478 = io_x[73] ? _GEN11477 : _GEN11473;
wire  _GEN11479 = io_x[33] ? _GEN11478 : _GEN10237;
wire  _GEN11480 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11481 = io_x[30] ? _GEN11480 : _GEN10239;
wire  _GEN11482 = io_x[26] ? _GEN11481 : _GEN10246;
wire  _GEN11483 = io_x[73] ? _GEN11482 : _GEN10243;
wire  _GEN11484 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11485 = io_x[30] ? _GEN11484 : _GEN10239;
wire  _GEN11486 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11487 = io_x[30] ? _GEN11486 : _GEN10239;
wire  _GEN11488 = io_x[26] ? _GEN11487 : _GEN11485;
wire  _GEN11489 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11490 = io_x[30] ? _GEN11489 : _GEN10239;
wire  _GEN11491 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11492 = io_x[30] ? _GEN10238 : _GEN11491;
wire  _GEN11493 = io_x[26] ? _GEN11492 : _GEN11490;
wire  _GEN11494 = io_x[73] ? _GEN11493 : _GEN11488;
wire  _GEN11495 = io_x[33] ? _GEN11494 : _GEN11483;
wire  _GEN11496 = io_x[28] ? _GEN11495 : _GEN11479;
wire  _GEN11497 = io_x[18] ? _GEN11496 : _GEN11471;
wire  _GEN11498 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11499 = io_x[30] ? _GEN11498 : _GEN10239;
wire  _GEN11500 = io_x[26] ? _GEN11499 : _GEN10246;
wire  _GEN11501 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11502 = io_x[26] ? _GEN10241 : _GEN11501;
wire  _GEN11503 = io_x[73] ? _GEN11502 : _GEN11500;
wire  _GEN11504 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11505 = io_x[30] ? _GEN10239 : _GEN11504;
wire  _GEN11506 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11507 = io_x[30] ? _GEN11506 : _GEN10239;
wire  _GEN11508 = io_x[26] ? _GEN11507 : _GEN11505;
wire  _GEN11509 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11510 = io_x[30] ? _GEN10239 : _GEN11509;
wire  _GEN11511 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11512 = io_x[26] ? _GEN11511 : _GEN11510;
wire  _GEN11513 = io_x[73] ? _GEN11512 : _GEN11508;
wire  _GEN11514 = io_x[33] ? _GEN11513 : _GEN11503;
wire  _GEN11515 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11516 = io_x[30] ? _GEN11515 : _GEN10239;
wire  _GEN11517 = io_x[26] ? _GEN11516 : _GEN10241;
wire  _GEN11518 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11519 = io_x[30] ? _GEN10239 : _GEN11518;
wire  _GEN11520 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11521 = io_x[26] ? _GEN11520 : _GEN11519;
wire  _GEN11522 = io_x[73] ? _GEN11521 : _GEN11517;
wire  _GEN11523 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11524 = io_x[30] ? _GEN11523 : _GEN10239;
wire  _GEN11525 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11526 = io_x[30] ? _GEN11525 : _GEN10238;
wire  _GEN11527 = io_x[26] ? _GEN11526 : _GEN11524;
wire  _GEN11528 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11529 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11530 = io_x[30] ? _GEN11529 : _GEN11528;
wire  _GEN11531 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11532 = io_x[30] ? _GEN11531 : _GEN10238;
wire  _GEN11533 = io_x[26] ? _GEN11532 : _GEN11530;
wire  _GEN11534 = io_x[73] ? _GEN11533 : _GEN11527;
wire  _GEN11535 = io_x[33] ? _GEN11534 : _GEN11522;
wire  _GEN11536 = io_x[28] ? _GEN11535 : _GEN11514;
wire  _GEN11537 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11538 = io_x[30] ? _GEN10239 : _GEN11537;
wire  _GEN11539 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11540 = io_x[30] ? _GEN11539 : _GEN10239;
wire  _GEN11541 = io_x[26] ? _GEN11540 : _GEN11538;
wire  _GEN11542 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11543 = io_x[30] ? _GEN11542 : _GEN10238;
wire  _GEN11544 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11545 = io_x[30] ? _GEN11544 : _GEN10239;
wire  _GEN11546 = io_x[26] ? _GEN11545 : _GEN11543;
wire  _GEN11547 = io_x[73] ? _GEN11546 : _GEN11541;
wire  _GEN11548 = io_x[33] ? _GEN11547 : _GEN10306;
wire  _GEN11549 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11550 = io_x[30] ? _GEN11549 : _GEN10239;
wire  _GEN11551 = io_x[26] ? _GEN11550 : _GEN10246;
wire  _GEN11552 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11553 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11554 = io_x[30] ? _GEN11553 : _GEN10239;
wire  _GEN11555 = io_x[26] ? _GEN11554 : _GEN11552;
wire  _GEN11556 = io_x[73] ? _GEN11555 : _GEN11551;
wire  _GEN11557 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11558 = io_x[30] ? _GEN11557 : _GEN10238;
wire  _GEN11559 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11560 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11561 = io_x[30] ? _GEN11560 : _GEN11559;
wire  _GEN11562 = io_x[26] ? _GEN11561 : _GEN11558;
wire  _GEN11563 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11564 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11565 = io_x[30] ? _GEN11564 : _GEN11563;
wire  _GEN11566 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11567 = io_x[30] ? _GEN11566 : _GEN10239;
wire  _GEN11568 = io_x[26] ? _GEN11567 : _GEN11565;
wire  _GEN11569 = io_x[73] ? _GEN11568 : _GEN11562;
wire  _GEN11570 = io_x[33] ? _GEN11569 : _GEN11556;
wire  _GEN11571 = io_x[28] ? _GEN11570 : _GEN11548;
wire  _GEN11572 = io_x[18] ? _GEN11571 : _GEN11536;
wire  _GEN11573 = io_x[25] ? _GEN11572 : _GEN11497;
wire  _GEN11574 = io_x[29] ? _GEN11573 : _GEN11450;
wire  _GEN11575 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11576 = io_x[30] ? _GEN10239 : _GEN11575;
wire  _GEN11577 = io_x[26] ? _GEN10246 : _GEN11576;
wire  _GEN11578 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11579 = io_x[30] ? _GEN11578 : _GEN10239;
wire  _GEN11580 = io_x[26] ? _GEN11579 : _GEN10241;
wire  _GEN11581 = io_x[73] ? _GEN11580 : _GEN11577;
wire  _GEN11582 = io_x[33] ? _GEN11581 : _GEN10306;
wire  _GEN11583 = io_x[73] ? _GEN10243 : _GEN10259;
wire  _GEN11584 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11585 = io_x[30] ? _GEN11584 : _GEN10239;
wire  _GEN11586 = io_x[26] ? _GEN11585 : _GEN10246;
wire  _GEN11587 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11588 = io_x[30] ? _GEN10239 : _GEN11587;
wire  _GEN11589 = io_x[26] ? _GEN11588 : _GEN10246;
wire  _GEN11590 = io_x[73] ? _GEN11589 : _GEN11586;
wire  _GEN11591 = io_x[33] ? _GEN11590 : _GEN11583;
wire  _GEN11592 = io_x[28] ? _GEN11591 : _GEN11582;
wire  _GEN11593 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11594 = io_x[26] ? _GEN11593 : _GEN10246;
wire  _GEN11595 = io_x[73] ? _GEN11594 : _GEN10243;
wire  _GEN11596 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11597 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11598 = io_x[30] ? _GEN11597 : _GEN11596;
wire  _GEN11599 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11600 = io_x[26] ? _GEN11599 : _GEN11598;
wire  _GEN11601 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11602 = io_x[26] ? _GEN11601 : _GEN10246;
wire  _GEN11603 = io_x[73] ? _GEN11602 : _GEN11600;
wire  _GEN11604 = io_x[33] ? _GEN11603 : _GEN11595;
wire  _GEN11605 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11606 = io_x[30] ? _GEN11605 : _GEN10239;
wire  _GEN11607 = io_x[26] ? _GEN11606 : _GEN10246;
wire  _GEN11608 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11609 = io_x[26] ? _GEN11608 : _GEN10246;
wire  _GEN11610 = io_x[73] ? _GEN11609 : _GEN11607;
wire  _GEN11611 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11612 = io_x[30] ? _GEN11611 : _GEN10238;
wire  _GEN11613 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11614 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11615 = io_x[30] ? _GEN11614 : _GEN11613;
wire  _GEN11616 = io_x[26] ? _GEN11615 : _GEN11612;
wire  _GEN11617 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11618 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11619 = io_x[30] ? _GEN11618 : _GEN11617;
wire  _GEN11620 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11621 = io_x[26] ? _GEN11620 : _GEN11619;
wire  _GEN11622 = io_x[73] ? _GEN11621 : _GEN11616;
wire  _GEN11623 = io_x[33] ? _GEN11622 : _GEN11610;
wire  _GEN11624 = io_x[28] ? _GEN11623 : _GEN11604;
wire  _GEN11625 = io_x[18] ? _GEN11624 : _GEN11592;
wire  _GEN11626 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11627 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11628 = io_x[30] ? _GEN11627 : _GEN11626;
wire  _GEN11629 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11630 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11631 = io_x[30] ? _GEN11630 : _GEN11629;
wire  _GEN11632 = io_x[26] ? _GEN11631 : _GEN11628;
wire  _GEN11633 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11634 = io_x[30] ? _GEN11633 : _GEN10239;
wire  _GEN11635 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11636 = io_x[26] ? _GEN11635 : _GEN11634;
wire  _GEN11637 = io_x[73] ? _GEN11636 : _GEN11632;
wire  _GEN11638 = io_x[33] ? _GEN11637 : _GEN10306;
wire  _GEN11639 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11640 = io_x[30] ? _GEN10239 : _GEN11639;
wire  _GEN11641 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11642 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11643 = io_x[30] ? _GEN11642 : _GEN11641;
wire  _GEN11644 = io_x[26] ? _GEN11643 : _GEN11640;
wire  _GEN11645 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11646 = io_x[26] ? _GEN11645 : _GEN10241;
wire  _GEN11647 = io_x[73] ? _GEN11646 : _GEN11644;
wire  _GEN11648 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11649 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11650 = io_x[30] ? _GEN11649 : _GEN11648;
wire  _GEN11651 = io_x[26] ? _GEN11650 : _GEN10246;
wire  _GEN11652 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN11653 = io_x[73] ? _GEN11652 : _GEN11651;
wire  _GEN11654 = io_x[33] ? _GEN11653 : _GEN11647;
wire  _GEN11655 = io_x[28] ? _GEN11654 : _GEN11638;
wire  _GEN11656 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11657 = io_x[30] ? _GEN11656 : _GEN10239;
wire  _GEN11658 = io_x[26] ? _GEN11657 : _GEN10246;
wire  _GEN11659 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11660 = io_x[30] ? _GEN11659 : _GEN10239;
wire  _GEN11661 = io_x[26] ? _GEN11660 : _GEN10241;
wire  _GEN11662 = io_x[73] ? _GEN11661 : _GEN11658;
wire  _GEN11663 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11664 = io_x[30] ? _GEN11663 : _GEN10239;
wire  _GEN11665 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11666 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11667 = io_x[30] ? _GEN11666 : _GEN11665;
wire  _GEN11668 = io_x[26] ? _GEN11667 : _GEN11664;
wire  _GEN11669 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11670 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11671 = io_x[30] ? _GEN10238 : _GEN11670;
wire  _GEN11672 = io_x[26] ? _GEN11671 : _GEN11669;
wire  _GEN11673 = io_x[73] ? _GEN11672 : _GEN11668;
wire  _GEN11674 = io_x[33] ? _GEN11673 : _GEN11662;
wire  _GEN11675 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11676 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11677 = io_x[30] ? _GEN11676 : _GEN11675;
wire  _GEN11678 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11679 = io_x[30] ? _GEN11678 : _GEN10239;
wire  _GEN11680 = io_x[26] ? _GEN11679 : _GEN11677;
wire  _GEN11681 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11682 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11683 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11684 = io_x[30] ? _GEN11683 : _GEN11682;
wire  _GEN11685 = io_x[26] ? _GEN11684 : _GEN11681;
wire  _GEN11686 = io_x[73] ? _GEN11685 : _GEN11680;
wire  _GEN11687 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11688 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11689 = io_x[30] ? _GEN11688 : _GEN11687;
wire  _GEN11690 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11691 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11692 = io_x[30] ? _GEN11691 : _GEN11690;
wire  _GEN11693 = io_x[26] ? _GEN11692 : _GEN11689;
wire  _GEN11694 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11695 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11696 = io_x[30] ? _GEN11695 : _GEN11694;
wire  _GEN11697 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11698 = io_x[30] ? _GEN11697 : _GEN10239;
wire  _GEN11699 = io_x[26] ? _GEN11698 : _GEN11696;
wire  _GEN11700 = io_x[73] ? _GEN11699 : _GEN11693;
wire  _GEN11701 = io_x[33] ? _GEN11700 : _GEN11686;
wire  _GEN11702 = io_x[28] ? _GEN11701 : _GEN11674;
wire  _GEN11703 = io_x[18] ? _GEN11702 : _GEN11655;
wire  _GEN11704 = io_x[25] ? _GEN11703 : _GEN11625;
wire  _GEN11705 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11706 = io_x[30] ? _GEN10239 : _GEN11705;
wire  _GEN11707 = io_x[26] ? _GEN11706 : _GEN10241;
wire  _GEN11708 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN11709 = io_x[73] ? _GEN11708 : _GEN11707;
wire  _GEN11710 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11711 = io_x[30] ? _GEN11710 : _GEN10238;
wire  _GEN11712 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11713 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11714 = io_x[30] ? _GEN11713 : _GEN11712;
wire  _GEN11715 = io_x[26] ? _GEN11714 : _GEN11711;
wire  _GEN11716 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11717 = io_x[30] ? _GEN11716 : _GEN10239;
wire  _GEN11718 = io_x[26] ? _GEN11717 : _GEN10246;
wire  _GEN11719 = io_x[73] ? _GEN11718 : _GEN11715;
wire  _GEN11720 = io_x[33] ? _GEN11719 : _GEN11709;
wire  _GEN11721 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11722 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11723 = io_x[30] ? _GEN11722 : _GEN11721;
wire  _GEN11724 = io_x[26] ? _GEN11723 : _GEN10241;
wire  _GEN11725 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11726 = io_x[30] ? _GEN11725 : _GEN10239;
wire  _GEN11727 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11728 = io_x[30] ? _GEN11727 : _GEN10238;
wire  _GEN11729 = io_x[26] ? _GEN11728 : _GEN11726;
wire  _GEN11730 = io_x[73] ? _GEN11729 : _GEN11724;
wire  _GEN11731 = io_x[33] ? _GEN11730 : _GEN10237;
wire  _GEN11732 = io_x[28] ? _GEN11731 : _GEN11720;
wire  _GEN11733 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11734 = io_x[30] ? _GEN10238 : _GEN11733;
wire  _GEN11735 = io_x[26] ? _GEN11734 : _GEN10241;
wire  _GEN11736 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11737 = io_x[30] ? _GEN10239 : _GEN11736;
wire  _GEN11738 = io_x[26] ? _GEN11737 : _GEN10246;
wire  _GEN11739 = io_x[73] ? _GEN11738 : _GEN11735;
wire  _GEN11740 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11741 = io_x[30] ? _GEN11740 : _GEN10238;
wire  _GEN11742 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11743 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11744 = io_x[30] ? _GEN11743 : _GEN11742;
wire  _GEN11745 = io_x[26] ? _GEN11744 : _GEN11741;
wire  _GEN11746 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11747 = io_x[26] ? _GEN10246 : _GEN11746;
wire  _GEN11748 = io_x[73] ? _GEN11747 : _GEN11745;
wire  _GEN11749 = io_x[33] ? _GEN11748 : _GEN11739;
wire  _GEN11750 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11751 = io_x[30] ? _GEN11750 : _GEN10238;
wire  _GEN11752 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11753 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11754 = io_x[30] ? _GEN11753 : _GEN11752;
wire  _GEN11755 = io_x[26] ? _GEN11754 : _GEN11751;
wire  _GEN11756 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11757 = io_x[30] ? _GEN11756 : _GEN10239;
wire  _GEN11758 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11759 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11760 = io_x[30] ? _GEN11759 : _GEN11758;
wire  _GEN11761 = io_x[26] ? _GEN11760 : _GEN11757;
wire  _GEN11762 = io_x[73] ? _GEN11761 : _GEN11755;
wire  _GEN11763 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11764 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11765 = io_x[30] ? _GEN11764 : _GEN11763;
wire  _GEN11766 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11767 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11768 = io_x[30] ? _GEN11767 : _GEN11766;
wire  _GEN11769 = io_x[26] ? _GEN11768 : _GEN11765;
wire  _GEN11770 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11771 = io_x[30] ? _GEN11770 : _GEN10239;
wire  _GEN11772 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11773 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11774 = io_x[30] ? _GEN11773 : _GEN11772;
wire  _GEN11775 = io_x[26] ? _GEN11774 : _GEN11771;
wire  _GEN11776 = io_x[73] ? _GEN11775 : _GEN11769;
wire  _GEN11777 = io_x[33] ? _GEN11776 : _GEN11762;
wire  _GEN11778 = io_x[28] ? _GEN11777 : _GEN11749;
wire  _GEN11779 = io_x[18] ? _GEN11778 : _GEN11732;
wire  _GEN11780 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11781 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11782 = io_x[30] ? _GEN10238 : _GEN11781;
wire  _GEN11783 = io_x[26] ? _GEN11782 : _GEN11780;
wire  _GEN11784 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11785 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11786 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11787 = io_x[30] ? _GEN11786 : _GEN11785;
wire  _GEN11788 = io_x[26] ? _GEN11787 : _GEN11784;
wire  _GEN11789 = io_x[73] ? _GEN11788 : _GEN11783;
wire  _GEN11790 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11791 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11792 = io_x[30] ? _GEN11791 : _GEN11790;
wire  _GEN11793 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11794 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11795 = io_x[30] ? _GEN11794 : _GEN11793;
wire  _GEN11796 = io_x[26] ? _GEN11795 : _GEN11792;
wire  _GEN11797 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11798 = io_x[30] ? _GEN10239 : _GEN11797;
wire  _GEN11799 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11800 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11801 = io_x[30] ? _GEN11800 : _GEN11799;
wire  _GEN11802 = io_x[26] ? _GEN11801 : _GEN11798;
wire  _GEN11803 = io_x[73] ? _GEN11802 : _GEN11796;
wire  _GEN11804 = io_x[33] ? _GEN11803 : _GEN11789;
wire  _GEN11805 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11806 = io_x[30] ? _GEN11805 : _GEN10238;
wire  _GEN11807 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11808 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11809 = io_x[30] ? _GEN11808 : _GEN11807;
wire  _GEN11810 = io_x[26] ? _GEN11809 : _GEN11806;
wire  _GEN11811 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11812 = io_x[30] ? _GEN10239 : _GEN11811;
wire  _GEN11813 = io_x[26] ? _GEN11812 : _GEN10246;
wire  _GEN11814 = io_x[73] ? _GEN11813 : _GEN11810;
wire  _GEN11815 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11816 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11817 = io_x[30] ? _GEN11816 : _GEN11815;
wire  _GEN11818 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11819 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11820 = io_x[30] ? _GEN11819 : _GEN11818;
wire  _GEN11821 = io_x[26] ? _GEN11820 : _GEN11817;
wire  _GEN11822 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11823 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11824 = io_x[30] ? _GEN11823 : _GEN11822;
wire  _GEN11825 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11826 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11827 = io_x[30] ? _GEN11826 : _GEN11825;
wire  _GEN11828 = io_x[26] ? _GEN11827 : _GEN11824;
wire  _GEN11829 = io_x[73] ? _GEN11828 : _GEN11821;
wire  _GEN11830 = io_x[33] ? _GEN11829 : _GEN11814;
wire  _GEN11831 = io_x[28] ? _GEN11830 : _GEN11804;
wire  _GEN11832 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11833 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11834 = io_x[30] ? _GEN11833 : _GEN11832;
wire  _GEN11835 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11836 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11837 = io_x[30] ? _GEN11836 : _GEN11835;
wire  _GEN11838 = io_x[26] ? _GEN11837 : _GEN11834;
wire  _GEN11839 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11840 = io_x[30] ? _GEN10238 : _GEN11839;
wire  _GEN11841 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11842 = io_x[30] ? _GEN11841 : _GEN10239;
wire  _GEN11843 = io_x[26] ? _GEN11842 : _GEN11840;
wire  _GEN11844 = io_x[73] ? _GEN11843 : _GEN11838;
wire  _GEN11845 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11846 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11847 = io_x[30] ? _GEN11846 : _GEN11845;
wire  _GEN11848 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11849 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11850 = io_x[30] ? _GEN11849 : _GEN11848;
wire  _GEN11851 = io_x[26] ? _GEN11850 : _GEN11847;
wire  _GEN11852 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11853 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11854 = io_x[30] ? _GEN11853 : _GEN11852;
wire  _GEN11855 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11856 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11857 = io_x[30] ? _GEN11856 : _GEN11855;
wire  _GEN11858 = io_x[26] ? _GEN11857 : _GEN11854;
wire  _GEN11859 = io_x[73] ? _GEN11858 : _GEN11851;
wire  _GEN11860 = io_x[33] ? _GEN11859 : _GEN11844;
wire  _GEN11861 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11862 = io_x[30] ? _GEN11861 : _GEN10239;
wire  _GEN11863 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11864 = io_x[30] ? _GEN11863 : _GEN10239;
wire  _GEN11865 = io_x[26] ? _GEN11864 : _GEN11862;
wire  _GEN11866 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11867 = io_x[30] ? _GEN11866 : _GEN10239;
wire  _GEN11868 = io_x[26] ? _GEN11867 : _GEN10241;
wire  _GEN11869 = io_x[73] ? _GEN11868 : _GEN11865;
wire  _GEN11870 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11871 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11872 = io_x[30] ? _GEN11871 : _GEN11870;
wire  _GEN11873 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11874 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11875 = io_x[30] ? _GEN11874 : _GEN11873;
wire  _GEN11876 = io_x[26] ? _GEN11875 : _GEN11872;
wire  _GEN11877 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11878 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11879 = io_x[30] ? _GEN11878 : _GEN11877;
wire  _GEN11880 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11881 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11882 = io_x[30] ? _GEN11881 : _GEN11880;
wire  _GEN11883 = io_x[26] ? _GEN11882 : _GEN11879;
wire  _GEN11884 = io_x[73] ? _GEN11883 : _GEN11876;
wire  _GEN11885 = io_x[33] ? _GEN11884 : _GEN11869;
wire  _GEN11886 = io_x[28] ? _GEN11885 : _GEN11860;
wire  _GEN11887 = io_x[18] ? _GEN11886 : _GEN11831;
wire  _GEN11888 = io_x[25] ? _GEN11887 : _GEN11779;
wire  _GEN11889 = io_x[29] ? _GEN11888 : _GEN11704;
wire  _GEN11890 = io_x[23] ? _GEN11889 : _GEN11574;
wire  _GEN11891 = io_x[31] ? _GEN11890 : _GEN11362;
wire  _GEN11892 = io_x[19] ? _GEN11891 : _GEN10966;
wire  _GEN11893 = io_x[73] ? _GEN10243 : _GEN10259;
wire  _GEN11894 = io_x[33] ? _GEN11893 : _GEN10237;
wire  _GEN11895 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11896 = io_x[26] ? _GEN10246 : _GEN11895;
wire  _GEN11897 = io_x[73] ? _GEN11896 : _GEN10259;
wire  _GEN11898 = io_x[73] ? _GEN10243 : _GEN10259;
wire  _GEN11899 = io_x[33] ? _GEN11898 : _GEN11897;
wire  _GEN11900 = io_x[28] ? _GEN11899 : _GEN11894;
wire  _GEN11901 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN11902 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11903 = io_x[30] ? _GEN11902 : _GEN10239;
wire  _GEN11904 = io_x[26] ? _GEN11903 : _GEN10241;
wire  _GEN11905 = io_x[73] ? _GEN11904 : _GEN11901;
wire  _GEN11906 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11907 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11908 = io_x[30] ? _GEN11907 : _GEN10239;
wire  _GEN11909 = io_x[26] ? _GEN11908 : _GEN11906;
wire  _GEN11910 = io_x[73] ? _GEN11909 : _GEN10243;
wire  _GEN11911 = io_x[33] ? _GEN11910 : _GEN11905;
wire  _GEN11912 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11913 = io_x[30] ? _GEN11912 : _GEN10239;
wire  _GEN11914 = io_x[26] ? _GEN11913 : _GEN10246;
wire  _GEN11915 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN11916 = io_x[73] ? _GEN11915 : _GEN11914;
wire  _GEN11917 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11918 = io_x[30] ? _GEN11917 : _GEN10239;
wire  _GEN11919 = io_x[26] ? _GEN11918 : _GEN10246;
wire  _GEN11920 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN11921 = io_x[73] ? _GEN11920 : _GEN11919;
wire  _GEN11922 = io_x[33] ? _GEN11921 : _GEN11916;
wire  _GEN11923 = io_x[28] ? _GEN11922 : _GEN11911;
wire  _GEN11924 = io_x[18] ? _GEN11923 : _GEN11900;
wire  _GEN11925 = io_x[73] ? _GEN10259 : _GEN10243;
wire  _GEN11926 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11927 = io_x[30] ? _GEN11926 : _GEN10239;
wire  _GEN11928 = io_x[26] ? _GEN11927 : _GEN10241;
wire  _GEN11929 = io_x[73] ? _GEN11928 : _GEN10243;
wire  _GEN11930 = io_x[33] ? _GEN11929 : _GEN11925;
wire  _GEN11931 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11932 = io_x[26] ? _GEN11931 : _GEN10246;
wire  _GEN11933 = io_x[73] ? _GEN11932 : _GEN10243;
wire  _GEN11934 = io_x[33] ? _GEN11933 : _GEN10306;
wire  _GEN11935 = io_x[28] ? _GEN11934 : _GEN11930;
wire  _GEN11936 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN11937 = io_x[73] ? _GEN10259 : _GEN11936;
wire  _GEN11938 = io_x[33] ? _GEN11937 : _GEN10306;
wire  _GEN11939 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11940 = io_x[30] ? _GEN10239 : _GEN11939;
wire  _GEN11941 = io_x[26] ? _GEN11940 : _GEN10246;
wire  _GEN11942 = io_x[73] ? _GEN10243 : _GEN11941;
wire  _GEN11943 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11944 = io_x[30] ? _GEN11943 : _GEN10239;
wire  _GEN11945 = io_x[26] ? _GEN11944 : _GEN10241;
wire  _GEN11946 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11947 = io_x[30] ? _GEN11946 : _GEN10238;
wire  _GEN11948 = io_x[26] ? _GEN11947 : _GEN10246;
wire  _GEN11949 = io_x[73] ? _GEN11948 : _GEN11945;
wire  _GEN11950 = io_x[33] ? _GEN11949 : _GEN11942;
wire  _GEN11951 = io_x[28] ? _GEN11950 : _GEN11938;
wire  _GEN11952 = io_x[18] ? _GEN11951 : _GEN11935;
wire  _GEN11953 = io_x[25] ? _GEN11952 : _GEN11924;
wire  _GEN11954 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11955 = io_x[30] ? _GEN11954 : _GEN10239;
wire  _GEN11956 = io_x[26] ? _GEN10241 : _GEN11955;
wire  _GEN11957 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN11958 = io_x[73] ? _GEN11957 : _GEN11956;
wire  _GEN11959 = io_x[33] ? _GEN11958 : _GEN10237;
wire  _GEN11960 = io_x[28] ? _GEN11021 : _GEN11959;
wire  _GEN11961 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11962 = io_x[26] ? _GEN11961 : _GEN10241;
wire  _GEN11963 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11964 = io_x[26] ? _GEN11963 : _GEN10241;
wire  _GEN11965 = io_x[73] ? _GEN11964 : _GEN11962;
wire  _GEN11966 = io_x[33] ? _GEN11965 : _GEN10306;
wire  _GEN11967 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN11968 = io_x[26] ? _GEN11967 : _GEN10241;
wire  _GEN11969 = io_x[73] ? _GEN10243 : _GEN11968;
wire  _GEN11970 = io_x[33] ? _GEN10237 : _GEN11969;
wire  _GEN11971 = io_x[28] ? _GEN11970 : _GEN11966;
wire  _GEN11972 = io_x[18] ? _GEN11971 : _GEN11960;
wire  _GEN11973 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11974 = io_x[26] ? _GEN11973 : _GEN10241;
wire  _GEN11975 = io_x[73] ? _GEN10259 : _GEN11974;
wire  _GEN11976 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN11977 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN11978 = io_x[73] ? _GEN11977 : _GEN11976;
wire  _GEN11979 = io_x[33] ? _GEN11978 : _GEN11975;
wire  _GEN11980 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN11981 = io_x[73] ? _GEN10243 : _GEN11980;
wire  _GEN11982 = io_x[33] ? _GEN11981 : _GEN10237;
wire  _GEN11983 = io_x[28] ? _GEN11982 : _GEN11979;
wire  _GEN11984 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11985 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11986 = io_x[30] ? _GEN11985 : _GEN11984;
wire  _GEN11987 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11988 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11989 = io_x[30] ? _GEN11988 : _GEN11987;
wire  _GEN11990 = io_x[26] ? _GEN11989 : _GEN11986;
wire  _GEN11991 = io_x[73] ? _GEN10259 : _GEN11990;
wire  _GEN11992 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN11993 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11994 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN11995 = io_x[30] ? _GEN11994 : _GEN11993;
wire  _GEN11996 = io_x[26] ? _GEN11995 : _GEN11992;
wire  _GEN11997 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN11998 = io_x[30] ? _GEN10239 : _GEN11997;
wire  _GEN11999 = io_x[26] ? _GEN11998 : _GEN10246;
wire  _GEN12000 = io_x[73] ? _GEN11999 : _GEN11996;
wire  _GEN12001 = io_x[33] ? _GEN12000 : _GEN11991;
wire  _GEN12002 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN12003 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN12004 = io_x[73] ? _GEN12003 : _GEN12002;
wire  _GEN12005 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN12006 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12007 = io_x[30] ? _GEN10239 : _GEN12006;
wire  _GEN12008 = io_x[26] ? _GEN12007 : _GEN10246;
wire  _GEN12009 = io_x[73] ? _GEN12008 : _GEN12005;
wire  _GEN12010 = io_x[33] ? _GEN12009 : _GEN12004;
wire  _GEN12011 = io_x[28] ? _GEN12010 : _GEN12001;
wire  _GEN12012 = io_x[18] ? _GEN12011 : _GEN11983;
wire  _GEN12013 = io_x[25] ? _GEN12012 : _GEN11972;
wire  _GEN12014 = io_x[29] ? _GEN12013 : _GEN11953;
wire  _GEN12015 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12016 = io_x[30] ? _GEN12015 : _GEN10239;
wire  _GEN12017 = io_x[26] ? _GEN12016 : _GEN10241;
wire  _GEN12018 = io_x[73] ? _GEN10259 : _GEN12017;
wire  _GEN12019 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12020 = io_x[26] ? _GEN12019 : _GEN10246;
wire  _GEN12021 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN12022 = io_x[73] ? _GEN12021 : _GEN12020;
wire  _GEN12023 = io_x[33] ? _GEN12022 : _GEN12018;
wire  _GEN12024 = io_x[28] ? _GEN12023 : _GEN10433;
wire  _GEN12025 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12026 = io_x[30] ? _GEN12025 : _GEN10238;
wire  _GEN12027 = io_x[26] ? _GEN10246 : _GEN12026;
wire  _GEN12028 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN12029 = io_x[73] ? _GEN12028 : _GEN12027;
wire  _GEN12030 = io_x[33] ? _GEN12029 : _GEN10306;
wire  _GEN12031 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12032 = io_x[30] ? _GEN12031 : _GEN10239;
wire  _GEN12033 = io_x[26] ? _GEN12032 : _GEN10241;
wire  _GEN12034 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12035 = io_x[30] ? _GEN12034 : _GEN10239;
wire  _GEN12036 = io_x[26] ? _GEN12035 : _GEN10241;
wire  _GEN12037 = io_x[73] ? _GEN12036 : _GEN12033;
wire  _GEN12038 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12039 = io_x[30] ? _GEN12038 : _GEN10239;
wire  _GEN12040 = io_x[26] ? _GEN12039 : _GEN10246;
wire  _GEN12041 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12042 = io_x[30] ? _GEN12041 : _GEN10239;
wire  _GEN12043 = io_x[26] ? _GEN12042 : _GEN10241;
wire  _GEN12044 = io_x[73] ? _GEN12043 : _GEN12040;
wire  _GEN12045 = io_x[33] ? _GEN12044 : _GEN12037;
wire  _GEN12046 = io_x[28] ? _GEN12045 : _GEN12030;
wire  _GEN12047 = io_x[18] ? _GEN12046 : _GEN12024;
wire  _GEN12048 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12049 = io_x[26] ? _GEN10246 : _GEN12048;
wire  _GEN12050 = io_x[73] ? _GEN12049 : _GEN10259;
wire  _GEN12051 = io_x[33] ? _GEN12050 : _GEN10306;
wire  _GEN12052 = io_x[28] ? _GEN12051 : _GEN11021;
wire  _GEN12053 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12054 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12055 = io_x[30] ? _GEN12054 : _GEN10239;
wire  _GEN12056 = io_x[26] ? _GEN12055 : _GEN12053;
wire  _GEN12057 = io_x[73] ? _GEN10243 : _GEN12056;
wire  _GEN12058 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN12059 = io_x[73] ? _GEN10243 : _GEN12058;
wire  _GEN12060 = io_x[33] ? _GEN12059 : _GEN12057;
wire  _GEN12061 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12062 = io_x[30] ? _GEN12061 : _GEN10238;
wire  _GEN12063 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12064 = io_x[30] ? _GEN12063 : _GEN10239;
wire  _GEN12065 = io_x[26] ? _GEN12064 : _GEN12062;
wire  _GEN12066 = io_x[73] ? _GEN10243 : _GEN12065;
wire  _GEN12067 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12068 = io_x[30] ? _GEN12067 : _GEN10238;
wire  _GEN12069 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12070 = io_x[30] ? _GEN12069 : _GEN10239;
wire  _GEN12071 = io_x[26] ? _GEN12070 : _GEN12068;
wire  _GEN12072 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12073 = io_x[30] ? _GEN12072 : _GEN10238;
wire  _GEN12074 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12075 = io_x[30] ? _GEN12074 : _GEN10239;
wire  _GEN12076 = io_x[26] ? _GEN12075 : _GEN12073;
wire  _GEN12077 = io_x[73] ? _GEN12076 : _GEN12071;
wire  _GEN12078 = io_x[33] ? _GEN12077 : _GEN12066;
wire  _GEN12079 = io_x[28] ? _GEN12078 : _GEN12060;
wire  _GEN12080 = io_x[18] ? _GEN12079 : _GEN12052;
wire  _GEN12081 = io_x[25] ? _GEN12080 : _GEN12047;
wire  _GEN12082 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12083 = io_x[30] ? _GEN10239 : _GEN12082;
wire  _GEN12084 = io_x[26] ? _GEN12083 : _GEN10241;
wire  _GEN12085 = io_x[73] ? _GEN10259 : _GEN12084;
wire  _GEN12086 = io_x[33] ? _GEN12085 : _GEN10306;
wire  _GEN12087 = io_x[28] ? _GEN10433 : _GEN12086;
wire  _GEN12088 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12089 = io_x[30] ? _GEN10239 : _GEN12088;
wire  _GEN12090 = io_x[26] ? _GEN12089 : _GEN10241;
wire  _GEN12091 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12092 = io_x[26] ? _GEN12091 : _GEN10241;
wire  _GEN12093 = io_x[73] ? _GEN12092 : _GEN12090;
wire  _GEN12094 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12095 = io_x[30] ? _GEN10239 : _GEN12094;
wire  _GEN12096 = io_x[26] ? _GEN12095 : _GEN10241;
wire  _GEN12097 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12098 = io_x[30] ? _GEN10239 : _GEN12097;
wire  _GEN12099 = io_x[26] ? _GEN12098 : _GEN10241;
wire  _GEN12100 = io_x[73] ? _GEN12099 : _GEN12096;
wire  _GEN12101 = io_x[33] ? _GEN12100 : _GEN12093;
wire  _GEN12102 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12103 = io_x[30] ? _GEN12102 : _GEN10239;
wire  _GEN12104 = io_x[26] ? _GEN10246 : _GEN12103;
wire  _GEN12105 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12106 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12107 = io_x[30] ? _GEN12106 : _GEN10239;
wire  _GEN12108 = io_x[26] ? _GEN12107 : _GEN12105;
wire  _GEN12109 = io_x[73] ? _GEN12108 : _GEN12104;
wire  _GEN12110 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12111 = io_x[30] ? _GEN10239 : _GEN12110;
wire  _GEN12112 = io_x[26] ? _GEN10246 : _GEN12111;
wire  _GEN12113 = io_x[73] ? _GEN12112 : _GEN10243;
wire  _GEN12114 = io_x[33] ? _GEN12113 : _GEN12109;
wire  _GEN12115 = io_x[28] ? _GEN12114 : _GEN12101;
wire  _GEN12116 = io_x[18] ? _GEN12115 : _GEN12087;
wire  _GEN12117 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12118 = io_x[30] ? _GEN12117 : _GEN10239;
wire  _GEN12119 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12120 = io_x[30] ? _GEN12119 : _GEN10239;
wire  _GEN12121 = io_x[26] ? _GEN12120 : _GEN12118;
wire  _GEN12122 = io_x[73] ? _GEN10259 : _GEN12121;
wire  _GEN12123 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12124 = io_x[30] ? _GEN12123 : _GEN10239;
wire  _GEN12125 = io_x[26] ? _GEN10241 : _GEN12124;
wire  _GEN12126 = io_x[73] ? _GEN10259 : _GEN12125;
wire  _GEN12127 = io_x[33] ? _GEN12126 : _GEN12122;
wire  _GEN12128 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12129 = io_x[26] ? _GEN10241 : _GEN12128;
wire  _GEN12130 = io_x[73] ? _GEN10243 : _GEN12129;
wire  _GEN12131 = io_x[73] ? _GEN10259 : _GEN10243;
wire  _GEN12132 = io_x[33] ? _GEN12131 : _GEN12130;
wire  _GEN12133 = io_x[28] ? _GEN12132 : _GEN12127;
wire  _GEN12134 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12135 = io_x[26] ? _GEN10241 : _GEN12134;
wire  _GEN12136 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12137 = io_x[30] ? _GEN12136 : _GEN10239;
wire  _GEN12138 = io_x[26] ? _GEN10241 : _GEN12137;
wire  _GEN12139 = io_x[73] ? _GEN12138 : _GEN12135;
wire  _GEN12140 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12141 = io_x[30] ? _GEN12140 : _GEN10239;
wire  _GEN12142 = io_x[26] ? _GEN10241 : _GEN12141;
wire  _GEN12143 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12144 = io_x[30] ? _GEN12143 : _GEN10239;
wire  _GEN12145 = io_x[26] ? _GEN10241 : _GEN12144;
wire  _GEN12146 = io_x[73] ? _GEN12145 : _GEN12142;
wire  _GEN12147 = io_x[33] ? _GEN12146 : _GEN12139;
wire  _GEN12148 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12149 = io_x[30] ? _GEN12148 : _GEN10239;
wire  _GEN12150 = io_x[26] ? _GEN12149 : _GEN10246;
wire  _GEN12151 = io_x[73] ? _GEN10259 : _GEN12150;
wire  _GEN12152 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12153 = io_x[30] ? _GEN12152 : _GEN10238;
wire  _GEN12154 = io_x[26] ? _GEN12153 : _GEN10246;
wire  _GEN12155 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12156 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12157 = io_x[30] ? _GEN12156 : _GEN10239;
wire  _GEN12158 = io_x[26] ? _GEN12157 : _GEN12155;
wire  _GEN12159 = io_x[73] ? _GEN12158 : _GEN12154;
wire  _GEN12160 = io_x[33] ? _GEN12159 : _GEN12151;
wire  _GEN12161 = io_x[28] ? _GEN12160 : _GEN12147;
wire  _GEN12162 = io_x[18] ? _GEN12161 : _GEN12133;
wire  _GEN12163 = io_x[25] ? _GEN12162 : _GEN12116;
wire  _GEN12164 = io_x[29] ? _GEN12163 : _GEN12081;
wire  _GEN12165 = io_x[23] ? _GEN12164 : _GEN12014;
wire  _GEN12166 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12167 = io_x[30] ? _GEN10239 : _GEN12166;
wire  _GEN12168 = io_x[26] ? _GEN12167 : _GEN10241;
wire  _GEN12169 = io_x[73] ? _GEN12168 : _GEN10243;
wire  _GEN12170 = io_x[33] ? _GEN12169 : _GEN10237;
wire  _GEN12171 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12172 = io_x[26] ? _GEN12171 : _GEN10241;
wire  _GEN12173 = io_x[73] ? _GEN10243 : _GEN12172;
wire  _GEN12174 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12175 = io_x[26] ? _GEN12174 : _GEN10241;
wire  _GEN12176 = io_x[73] ? _GEN10243 : _GEN12175;
wire  _GEN12177 = io_x[33] ? _GEN12176 : _GEN12173;
wire  _GEN12178 = io_x[28] ? _GEN12177 : _GEN12170;
wire  _GEN12179 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12180 = io_x[26] ? _GEN12179 : _GEN10241;
wire  _GEN12181 = io_x[73] ? _GEN10243 : _GEN12180;
wire  _GEN12182 = io_x[33] ? _GEN12181 : _GEN10237;
wire  _GEN12183 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12184 = io_x[26] ? _GEN12183 : _GEN10241;
wire  _GEN12185 = io_x[73] ? _GEN12184 : _GEN10259;
wire  _GEN12186 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12187 = io_x[30] ? _GEN12186 : _GEN10238;
wire  _GEN12188 = io_x[26] ? _GEN12187 : _GEN10241;
wire  _GEN12189 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12190 = io_x[30] ? _GEN12189 : _GEN10238;
wire  _GEN12191 = io_x[26] ? _GEN12190 : _GEN10241;
wire  _GEN12192 = io_x[73] ? _GEN12191 : _GEN12188;
wire  _GEN12193 = io_x[33] ? _GEN12192 : _GEN12185;
wire  _GEN12194 = io_x[28] ? _GEN12193 : _GEN12182;
wire  _GEN12195 = io_x[18] ? _GEN12194 : _GEN12178;
wire  _GEN12196 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12197 = io_x[30] ? _GEN12196 : _GEN10239;
wire  _GEN12198 = io_x[26] ? _GEN12197 : _GEN10241;
wire  _GEN12199 = io_x[73] ? _GEN12198 : _GEN10243;
wire  _GEN12200 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12201 = io_x[30] ? _GEN12200 : _GEN10238;
wire  _GEN12202 = io_x[26] ? _GEN12201 : _GEN10241;
wire  _GEN12203 = io_x[73] ? _GEN12202 : _GEN10243;
wire  _GEN12204 = io_x[33] ? _GEN12203 : _GEN12199;
wire  _GEN12205 = io_x[28] ? _GEN11021 : _GEN12204;
wire  _GEN12206 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12207 = io_x[30] ? _GEN12206 : _GEN10238;
wire  _GEN12208 = io_x[26] ? _GEN10241 : _GEN12207;
wire  _GEN12209 = io_x[73] ? _GEN10259 : _GEN12208;
wire  _GEN12210 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN12211 = io_x[73] ? _GEN10243 : _GEN12210;
wire  _GEN12212 = io_x[33] ? _GEN12211 : _GEN12209;
wire  _GEN12213 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12214 = io_x[30] ? _GEN10239 : _GEN12213;
wire  _GEN12215 = io_x[26] ? _GEN10246 : _GEN12214;
wire  _GEN12216 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12217 = io_x[30] ? _GEN10238 : _GEN12216;
wire  _GEN12218 = io_x[26] ? _GEN10241 : _GEN12217;
wire  _GEN12219 = io_x[73] ? _GEN12218 : _GEN12215;
wire  _GEN12220 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12221 = io_x[30] ? _GEN10238 : _GEN12220;
wire  _GEN12222 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12223 = io_x[30] ? _GEN12222 : _GEN10238;
wire  _GEN12224 = io_x[26] ? _GEN12223 : _GEN12221;
wire  _GEN12225 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12226 = io_x[30] ? _GEN12225 : _GEN10239;
wire  _GEN12227 = io_x[26] ? _GEN12226 : _GEN10246;
wire  _GEN12228 = io_x[73] ? _GEN12227 : _GEN12224;
wire  _GEN12229 = io_x[33] ? _GEN12228 : _GEN12219;
wire  _GEN12230 = io_x[28] ? _GEN12229 : _GEN12212;
wire  _GEN12231 = io_x[18] ? _GEN12230 : _GEN12205;
wire  _GEN12232 = io_x[25] ? _GEN12231 : _GEN12195;
wire  _GEN12233 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12234 = io_x[26] ? _GEN12233 : _GEN10246;
wire  _GEN12235 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12236 = io_x[30] ? _GEN12235 : _GEN10239;
wire  _GEN12237 = io_x[26] ? _GEN12236 : _GEN10241;
wire  _GEN12238 = io_x[73] ? _GEN12237 : _GEN12234;
wire  _GEN12239 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12240 = io_x[26] ? _GEN12239 : _GEN10246;
wire  _GEN12241 = io_x[73] ? _GEN10243 : _GEN12240;
wire  _GEN12242 = io_x[33] ? _GEN12241 : _GEN12238;
wire  _GEN12243 = io_x[73] ? _GEN10259 : _GEN10243;
wire  _GEN12244 = io_x[33] ? _GEN10237 : _GEN12243;
wire  _GEN12245 = io_x[28] ? _GEN12244 : _GEN12242;
wire  _GEN12246 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12247 = io_x[26] ? _GEN12246 : _GEN10246;
wire  _GEN12248 = io_x[73] ? _GEN10243 : _GEN12247;
wire  _GEN12249 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12250 = io_x[30] ? _GEN12249 : _GEN10239;
wire  _GEN12251 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12252 = io_x[26] ? _GEN12251 : _GEN12250;
wire  _GEN12253 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12254 = io_x[30] ? _GEN12253 : _GEN10238;
wire  _GEN12255 = io_x[26] ? _GEN12254 : _GEN10241;
wire  _GEN12256 = io_x[73] ? _GEN12255 : _GEN12252;
wire  _GEN12257 = io_x[33] ? _GEN12256 : _GEN12248;
wire  _GEN12258 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12259 = io_x[30] ? _GEN10239 : _GEN12258;
wire  _GEN12260 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12261 = io_x[26] ? _GEN12260 : _GEN12259;
wire  _GEN12262 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN12263 = io_x[73] ? _GEN12262 : _GEN12261;
wire  _GEN12264 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12265 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12266 = io_x[30] ? _GEN12265 : _GEN12264;
wire  _GEN12267 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12268 = io_x[26] ? _GEN12267 : _GEN12266;
wire  _GEN12269 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12270 = io_x[30] ? _GEN10239 : _GEN12269;
wire  _GEN12271 = io_x[26] ? _GEN10246 : _GEN12270;
wire  _GEN12272 = io_x[73] ? _GEN12271 : _GEN12268;
wire  _GEN12273 = io_x[33] ? _GEN12272 : _GEN12263;
wire  _GEN12274 = io_x[28] ? _GEN12273 : _GEN12257;
wire  _GEN12275 = io_x[18] ? _GEN12274 : _GEN12245;
wire  _GEN12276 = io_x[73] ? _GEN10259 : _GEN10243;
wire  _GEN12277 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12278 = io_x[30] ? _GEN12277 : _GEN10239;
wire  _GEN12279 = io_x[26] ? _GEN12278 : _GEN10241;
wire  _GEN12280 = io_x[73] ? _GEN10243 : _GEN12279;
wire  _GEN12281 = io_x[33] ? _GEN12280 : _GEN12276;
wire  _GEN12282 = io_x[73] ? _GEN10243 : _GEN10259;
wire  _GEN12283 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12284 = io_x[30] ? _GEN12283 : _GEN10238;
wire  _GEN12285 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12286 = io_x[30] ? _GEN12285 : _GEN10239;
wire  _GEN12287 = io_x[26] ? _GEN12286 : _GEN12284;
wire  _GEN12288 = io_x[73] ? _GEN12287 : _GEN10259;
wire  _GEN12289 = io_x[33] ? _GEN12288 : _GEN12282;
wire  _GEN12290 = io_x[28] ? _GEN12289 : _GEN12281;
wire  _GEN12291 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12292 = io_x[30] ? _GEN10238 : _GEN12291;
wire  _GEN12293 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12294 = io_x[30] ? _GEN12293 : _GEN10239;
wire  _GEN12295 = io_x[26] ? _GEN12294 : _GEN12292;
wire  _GEN12296 = io_x[73] ? _GEN10243 : _GEN12295;
wire  _GEN12297 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12298 = io_x[30] ? _GEN12297 : _GEN10239;
wire  _GEN12299 = io_x[26] ? _GEN12298 : _GEN10241;
wire  _GEN12300 = io_x[73] ? _GEN10259 : _GEN12299;
wire  _GEN12301 = io_x[33] ? _GEN12300 : _GEN12296;
wire  _GEN12302 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12303 = io_x[26] ? _GEN10241 : _GEN12302;
wire  _GEN12304 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN12305 = io_x[73] ? _GEN12304 : _GEN12303;
wire  _GEN12306 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12307 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12308 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12309 = io_x[30] ? _GEN12308 : _GEN12307;
wire  _GEN12310 = io_x[26] ? _GEN12309 : _GEN12306;
wire  _GEN12311 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12312 = io_x[30] ? _GEN12311 : _GEN10239;
wire  _GEN12313 = io_x[26] ? _GEN12312 : _GEN10246;
wire  _GEN12314 = io_x[73] ? _GEN12313 : _GEN12310;
wire  _GEN12315 = io_x[33] ? _GEN12314 : _GEN12305;
wire  _GEN12316 = io_x[28] ? _GEN12315 : _GEN12301;
wire  _GEN12317 = io_x[18] ? _GEN12316 : _GEN12290;
wire  _GEN12318 = io_x[25] ? _GEN12317 : _GEN12275;
wire  _GEN12319 = io_x[29] ? _GEN12318 : _GEN12232;
wire  _GEN12320 = io_x[33] ? _GEN10306 : _GEN10237;
wire  _GEN12321 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12322 = io_x[30] ? _GEN12321 : _GEN10239;
wire  _GEN12323 = io_x[26] ? _GEN10241 : _GEN12322;
wire  _GEN12324 = io_x[73] ? _GEN10259 : _GEN12323;
wire  _GEN12325 = io_x[33] ? _GEN10237 : _GEN12324;
wire  _GEN12326 = io_x[28] ? _GEN12325 : _GEN12320;
wire  _GEN12327 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12328 = io_x[26] ? _GEN10241 : _GEN12327;
wire  _GEN12329 = io_x[73] ? _GEN10243 : _GEN12328;
wire  _GEN12330 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12331 = io_x[26] ? _GEN10241 : _GEN12330;
wire  _GEN12332 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12333 = io_x[30] ? _GEN12332 : _GEN10238;
wire  _GEN12334 = io_x[26] ? _GEN12333 : _GEN10246;
wire  _GEN12335 = io_x[73] ? _GEN12334 : _GEN12331;
wire  _GEN12336 = io_x[33] ? _GEN12335 : _GEN12329;
wire  _GEN12337 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12338 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12339 = io_x[30] ? _GEN12338 : _GEN12337;
wire  _GEN12340 = io_x[26] ? _GEN12339 : _GEN10241;
wire  _GEN12341 = io_x[73] ? _GEN12340 : _GEN10259;
wire  _GEN12342 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12343 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12344 = io_x[30] ? _GEN12343 : _GEN12342;
wire  _GEN12345 = io_x[26] ? _GEN12344 : _GEN10241;
wire  _GEN12346 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12347 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12348 = io_x[30] ? _GEN12347 : _GEN12346;
wire  _GEN12349 = io_x[26] ? _GEN12348 : _GEN10246;
wire  _GEN12350 = io_x[73] ? _GEN12349 : _GEN12345;
wire  _GEN12351 = io_x[33] ? _GEN12350 : _GEN12341;
wire  _GEN12352 = io_x[28] ? _GEN12351 : _GEN12336;
wire  _GEN12353 = io_x[18] ? _GEN12352 : _GEN12326;
wire  _GEN12354 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12355 = io_x[30] ? _GEN12354 : _GEN10238;
wire  _GEN12356 = io_x[26] ? _GEN12355 : _GEN10246;
wire  _GEN12357 = io_x[73] ? _GEN10259 : _GEN12356;
wire  _GEN12358 = io_x[33] ? _GEN12357 : _GEN10306;
wire  _GEN12359 = io_x[28] ? _GEN12358 : _GEN10433;
wire  _GEN12360 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN12361 = io_x[73] ? _GEN10243 : _GEN12360;
wire  _GEN12362 = io_x[33] ? _GEN10237 : _GEN12361;
wire  _GEN12363 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12364 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12365 = io_x[30] ? _GEN12364 : _GEN12363;
wire  _GEN12366 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12367 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12368 = io_x[30] ? _GEN12367 : _GEN12366;
wire  _GEN12369 = io_x[26] ? _GEN12368 : _GEN12365;
wire  _GEN12370 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12371 = io_x[30] ? _GEN12370 : _GEN10239;
wire  _GEN12372 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12373 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12374 = io_x[30] ? _GEN12373 : _GEN12372;
wire  _GEN12375 = io_x[26] ? _GEN12374 : _GEN12371;
wire  _GEN12376 = io_x[73] ? _GEN12375 : _GEN12369;
wire  _GEN12377 = io_x[33] ? _GEN12376 : _GEN10237;
wire  _GEN12378 = io_x[28] ? _GEN12377 : _GEN12362;
wire  _GEN12379 = io_x[18] ? _GEN12378 : _GEN12359;
wire  _GEN12380 = io_x[25] ? _GEN12379 : _GEN12353;
wire  _GEN12381 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12382 = io_x[30] ? _GEN12381 : _GEN10239;
wire  _GEN12383 = io_x[26] ? _GEN12382 : _GEN10241;
wire  _GEN12384 = io_x[73] ? _GEN12383 : _GEN10243;
wire  _GEN12385 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12386 = io_x[30] ? _GEN12385 : _GEN10238;
wire  _GEN12387 = io_x[26] ? _GEN12386 : _GEN10241;
wire  _GEN12388 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12389 = io_x[30] ? _GEN12388 : _GEN10238;
wire  _GEN12390 = io_x[26] ? _GEN12389 : _GEN10241;
wire  _GEN12391 = io_x[73] ? _GEN12390 : _GEN12387;
wire  _GEN12392 = io_x[33] ? _GEN12391 : _GEN12384;
wire  _GEN12393 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12394 = io_x[26] ? _GEN12393 : _GEN10241;
wire  _GEN12395 = io_x[73] ? _GEN10259 : _GEN12394;
wire  _GEN12396 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12397 = io_x[30] ? _GEN10239 : _GEN12396;
wire  _GEN12398 = io_x[26] ? _GEN12397 : _GEN10241;
wire  _GEN12399 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12400 = io_x[30] ? _GEN10239 : _GEN12399;
wire  _GEN12401 = io_x[26] ? _GEN12400 : _GEN10241;
wire  _GEN12402 = io_x[73] ? _GEN12401 : _GEN12398;
wire  _GEN12403 = io_x[33] ? _GEN12402 : _GEN12395;
wire  _GEN12404 = io_x[28] ? _GEN12403 : _GEN12392;
wire  _GEN12405 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12406 = io_x[26] ? _GEN12405 : _GEN10241;
wire  _GEN12407 = io_x[73] ? _GEN10259 : _GEN12406;
wire  _GEN12408 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12409 = io_x[30] ? _GEN12408 : _GEN10239;
wire  _GEN12410 = io_x[26] ? _GEN12409 : _GEN10246;
wire  _GEN12411 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12412 = io_x[30] ? _GEN12411 : _GEN10238;
wire  _GEN12413 = io_x[26] ? _GEN12412 : _GEN10241;
wire  _GEN12414 = io_x[73] ? _GEN12413 : _GEN12410;
wire  _GEN12415 = io_x[33] ? _GEN12414 : _GEN12407;
wire  _GEN12416 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12417 = io_x[30] ? _GEN10239 : _GEN12416;
wire  _GEN12418 = io_x[26] ? _GEN12417 : _GEN10241;
wire  _GEN12419 = io_x[73] ? _GEN10259 : _GEN12418;
wire  _GEN12420 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12421 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12422 = io_x[30] ? _GEN12421 : _GEN12420;
wire  _GEN12423 = io_x[26] ? _GEN12422 : _GEN10241;
wire  _GEN12424 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12425 = io_x[30] ? _GEN10238 : _GEN12424;
wire  _GEN12426 = io_x[26] ? _GEN12425 : _GEN10241;
wire  _GEN12427 = io_x[73] ? _GEN12426 : _GEN12423;
wire  _GEN12428 = io_x[33] ? _GEN12427 : _GEN12419;
wire  _GEN12429 = io_x[28] ? _GEN12428 : _GEN12415;
wire  _GEN12430 = io_x[18] ? _GEN12429 : _GEN12404;
wire  _GEN12431 = io_x[73] ? _GEN10259 : _GEN10243;
wire  _GEN12432 = io_x[73] ? _GEN10259 : _GEN10243;
wire  _GEN12433 = io_x[33] ? _GEN12432 : _GEN12431;
wire  _GEN12434 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12435 = io_x[30] ? _GEN12434 : _GEN10239;
wire  _GEN12436 = io_x[26] ? _GEN12435 : _GEN10241;
wire  _GEN12437 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12438 = io_x[30] ? _GEN12437 : _GEN10239;
wire  _GEN12439 = io_x[26] ? _GEN12438 : _GEN10246;
wire  _GEN12440 = io_x[73] ? _GEN12439 : _GEN12436;
wire  _GEN12441 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12442 = io_x[26] ? _GEN10241 : _GEN12441;
wire  _GEN12443 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12444 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12445 = io_x[30] ? _GEN12444 : _GEN10239;
wire  _GEN12446 = io_x[26] ? _GEN12445 : _GEN12443;
wire  _GEN12447 = io_x[73] ? _GEN12446 : _GEN12442;
wire  _GEN12448 = io_x[33] ? _GEN12447 : _GEN12440;
wire  _GEN12449 = io_x[28] ? _GEN12448 : _GEN12433;
wire  _GEN12450 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12451 = io_x[30] ? _GEN10239 : _GEN12450;
wire  _GEN12452 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12453 = io_x[26] ? _GEN12452 : _GEN12451;
wire  _GEN12454 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12455 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12456 = io_x[30] ? _GEN12455 : _GEN12454;
wire  _GEN12457 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12458 = io_x[26] ? _GEN12457 : _GEN12456;
wire  _GEN12459 = io_x[73] ? _GEN12458 : _GEN12453;
wire  _GEN12460 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12461 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12462 = io_x[30] ? _GEN12461 : _GEN12460;
wire  _GEN12463 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12464 = io_x[26] ? _GEN12463 : _GEN12462;
wire  _GEN12465 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12466 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12467 = io_x[30] ? _GEN12466 : _GEN12465;
wire  _GEN12468 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12469 = io_x[26] ? _GEN12468 : _GEN12467;
wire  _GEN12470 = io_x[73] ? _GEN12469 : _GEN12464;
wire  _GEN12471 = io_x[33] ? _GEN12470 : _GEN12459;
wire  _GEN12472 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12473 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12474 = io_x[30] ? _GEN12473 : _GEN12472;
wire  _GEN12475 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12476 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12477 = io_x[30] ? _GEN12476 : _GEN12475;
wire  _GEN12478 = io_x[26] ? _GEN12477 : _GEN12474;
wire  _GEN12479 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12480 = io_x[30] ? _GEN12479 : _GEN10239;
wire  _GEN12481 = io_x[26] ? _GEN12480 : _GEN10246;
wire  _GEN12482 = io_x[73] ? _GEN12481 : _GEN12478;
wire  _GEN12483 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12484 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12485 = io_x[30] ? _GEN12484 : _GEN12483;
wire  _GEN12486 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12487 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12488 = io_x[30] ? _GEN12487 : _GEN12486;
wire  _GEN12489 = io_x[26] ? _GEN12488 : _GEN12485;
wire  _GEN12490 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12491 = io_x[30] ? _GEN10238 : _GEN12490;
wire  _GEN12492 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12493 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12494 = io_x[30] ? _GEN12493 : _GEN12492;
wire  _GEN12495 = io_x[26] ? _GEN12494 : _GEN12491;
wire  _GEN12496 = io_x[73] ? _GEN12495 : _GEN12489;
wire  _GEN12497 = io_x[33] ? _GEN12496 : _GEN12482;
wire  _GEN12498 = io_x[28] ? _GEN12497 : _GEN12471;
wire  _GEN12499 = io_x[18] ? _GEN12498 : _GEN12449;
wire  _GEN12500 = io_x[25] ? _GEN12499 : _GEN12430;
wire  _GEN12501 = io_x[29] ? _GEN12500 : _GEN12380;
wire  _GEN12502 = io_x[23] ? _GEN12501 : _GEN12319;
wire  _GEN12503 = io_x[31] ? _GEN12502 : _GEN12165;
wire  _GEN12504 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN12505 = io_x[73] ? _GEN10243 : _GEN12504;
wire  _GEN12506 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12507 = io_x[30] ? _GEN12506 : _GEN10238;
wire  _GEN12508 = io_x[26] ? _GEN10241 : _GEN12507;
wire  _GEN12509 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12510 = io_x[30] ? _GEN12509 : _GEN10239;
wire  _GEN12511 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12512 = io_x[26] ? _GEN12511 : _GEN12510;
wire  _GEN12513 = io_x[73] ? _GEN12512 : _GEN12508;
wire  _GEN12514 = io_x[33] ? _GEN12513 : _GEN12505;
wire  _GEN12515 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12516 = io_x[30] ? _GEN12515 : _GEN10238;
wire  _GEN12517 = io_x[26] ? _GEN12516 : _GEN10241;
wire  _GEN12518 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN12519 = io_x[73] ? _GEN12518 : _GEN12517;
wire  _GEN12520 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12521 = io_x[30] ? _GEN12520 : _GEN10238;
wire  _GEN12522 = io_x[26] ? _GEN12521 : _GEN10241;
wire  _GEN12523 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN12524 = io_x[73] ? _GEN12523 : _GEN12522;
wire  _GEN12525 = io_x[33] ? _GEN12524 : _GEN12519;
wire  _GEN12526 = io_x[28] ? _GEN12525 : _GEN12514;
wire  _GEN12527 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12528 = io_x[30] ? _GEN12527 : _GEN10239;
wire  _GEN12529 = io_x[26] ? _GEN10241 : _GEN12528;
wire  _GEN12530 = io_x[73] ? _GEN10243 : _GEN12529;
wire  _GEN12531 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12532 = io_x[30] ? _GEN12531 : _GEN10238;
wire  _GEN12533 = io_x[26] ? _GEN10241 : _GEN12532;
wire  _GEN12534 = io_x[73] ? _GEN10243 : _GEN12533;
wire  _GEN12535 = io_x[33] ? _GEN12534 : _GEN12530;
wire  _GEN12536 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12537 = io_x[30] ? _GEN12536 : _GEN10239;
wire  _GEN12538 = io_x[26] ? _GEN12537 : _GEN10246;
wire  _GEN12539 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12540 = io_x[30] ? _GEN12539 : _GEN10239;
wire  _GEN12541 = io_x[26] ? _GEN10241 : _GEN12540;
wire  _GEN12542 = io_x[73] ? _GEN12541 : _GEN12538;
wire  _GEN12543 = io_x[33] ? _GEN12542 : _GEN10237;
wire  _GEN12544 = io_x[28] ? _GEN12543 : _GEN12535;
wire  _GEN12545 = io_x[18] ? _GEN12544 : _GEN12526;
wire  _GEN12546 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12547 = io_x[26] ? _GEN12546 : _GEN10241;
wire  _GEN12548 = io_x[73] ? _GEN12547 : _GEN10259;
wire  _GEN12549 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12550 = io_x[26] ? _GEN12549 : _GEN10241;
wire  _GEN12551 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12552 = io_x[30] ? _GEN12551 : _GEN10239;
wire  _GEN12553 = io_x[26] ? _GEN12552 : _GEN10246;
wire  _GEN12554 = io_x[73] ? _GEN12553 : _GEN12550;
wire  _GEN12555 = io_x[33] ? _GEN12554 : _GEN12548;
wire  _GEN12556 = io_x[28] ? _GEN12555 : _GEN10433;
wire  _GEN12557 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12558 = io_x[30] ? _GEN12557 : _GEN10239;
wire  _GEN12559 = io_x[26] ? _GEN12558 : _GEN10241;
wire  _GEN12560 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12561 = io_x[26] ? _GEN12560 : _GEN10241;
wire  _GEN12562 = io_x[73] ? _GEN12561 : _GEN12559;
wire  _GEN12563 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12564 = io_x[30] ? _GEN12563 : _GEN10239;
wire  _GEN12565 = io_x[26] ? _GEN12564 : _GEN10246;
wire  _GEN12566 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN12567 = io_x[73] ? _GEN12566 : _GEN12565;
wire  _GEN12568 = io_x[33] ? _GEN12567 : _GEN12562;
wire  _GEN12569 = io_x[28] ? _GEN12568 : _GEN11021;
wire  _GEN12570 = io_x[18] ? _GEN12569 : _GEN12556;
wire  _GEN12571 = io_x[25] ? _GEN12570 : _GEN12545;
wire  _GEN12572 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12573 = io_x[26] ? _GEN12572 : _GEN10241;
wire  _GEN12574 = io_x[73] ? _GEN12573 : _GEN10243;
wire  _GEN12575 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12576 = io_x[30] ? _GEN12575 : _GEN10239;
wire  _GEN12577 = io_x[26] ? _GEN12576 : _GEN10241;
wire  _GEN12578 = io_x[73] ? _GEN10243 : _GEN12577;
wire  _GEN12579 = io_x[33] ? _GEN12578 : _GEN12574;
wire  _GEN12580 = io_x[73] ? _GEN10259 : _GEN10243;
wire  _GEN12581 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12582 = io_x[30] ? _GEN12581 : _GEN10238;
wire  _GEN12583 = io_x[26] ? _GEN10246 : _GEN12582;
wire  _GEN12584 = io_x[73] ? _GEN12583 : _GEN10243;
wire  _GEN12585 = io_x[33] ? _GEN12584 : _GEN12580;
wire  _GEN12586 = io_x[28] ? _GEN12585 : _GEN12579;
wire  _GEN12587 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12588 = io_x[30] ? _GEN10239 : _GEN12587;
wire  _GEN12589 = io_x[26] ? _GEN12588 : _GEN10241;
wire  _GEN12590 = io_x[73] ? _GEN10259 : _GEN12589;
wire  _GEN12591 = io_x[33] ? _GEN12590 : _GEN10306;
wire  _GEN12592 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12593 = io_x[26] ? _GEN12592 : _GEN10241;
wire  _GEN12594 = io_x[73] ? _GEN10243 : _GEN12593;
wire  _GEN12595 = io_x[33] ? _GEN12594 : _GEN10237;
wire  _GEN12596 = io_x[28] ? _GEN12595 : _GEN12591;
wire  _GEN12597 = io_x[18] ? _GEN12596 : _GEN12586;
wire  _GEN12598 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12599 = io_x[26] ? _GEN12598 : _GEN10241;
wire  _GEN12600 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12601 = io_x[26] ? _GEN12600 : _GEN10241;
wire  _GEN12602 = io_x[73] ? _GEN12601 : _GEN12599;
wire  _GEN12603 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12604 = io_x[30] ? _GEN12603 : _GEN10239;
wire  _GEN12605 = io_x[26] ? _GEN12604 : _GEN10241;
wire  _GEN12606 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12607 = io_x[30] ? _GEN12606 : _GEN10239;
wire  _GEN12608 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12609 = io_x[30] ? _GEN10238 : _GEN12608;
wire  _GEN12610 = io_x[26] ? _GEN12609 : _GEN12607;
wire  _GEN12611 = io_x[73] ? _GEN12610 : _GEN12605;
wire  _GEN12612 = io_x[33] ? _GEN12611 : _GEN12602;
wire  _GEN12613 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12614 = io_x[30] ? _GEN12613 : _GEN10238;
wire  _GEN12615 = io_x[26] ? _GEN12614 : _GEN10241;
wire  _GEN12616 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12617 = io_x[30] ? _GEN12616 : _GEN10239;
wire  _GEN12618 = io_x[26] ? _GEN12617 : _GEN10241;
wire  _GEN12619 = io_x[73] ? _GEN12618 : _GEN12615;
wire  _GEN12620 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12621 = io_x[30] ? _GEN12620 : _GEN10238;
wire  _GEN12622 = io_x[26] ? _GEN12621 : _GEN10241;
wire  _GEN12623 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12624 = io_x[30] ? _GEN12623 : _GEN10239;
wire  _GEN12625 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12626 = io_x[30] ? _GEN12625 : _GEN10239;
wire  _GEN12627 = io_x[26] ? _GEN12626 : _GEN12624;
wire  _GEN12628 = io_x[73] ? _GEN12627 : _GEN12622;
wire  _GEN12629 = io_x[33] ? _GEN12628 : _GEN12619;
wire  _GEN12630 = io_x[28] ? _GEN12629 : _GEN12612;
wire  _GEN12631 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12632 = io_x[30] ? _GEN10239 : _GEN12631;
wire  _GEN12633 = io_x[26] ? _GEN12632 : _GEN10241;
wire  _GEN12634 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12635 = io_x[30] ? _GEN12634 : _GEN10238;
wire  _GEN12636 = io_x[26] ? _GEN10241 : _GEN12635;
wire  _GEN12637 = io_x[73] ? _GEN12636 : _GEN12633;
wire  _GEN12638 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12639 = io_x[30] ? _GEN10239 : _GEN12638;
wire  _GEN12640 = io_x[26] ? _GEN12639 : _GEN10246;
wire  _GEN12641 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12642 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12643 = io_x[30] ? _GEN12642 : _GEN12641;
wire  _GEN12644 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12645 = io_x[30] ? _GEN10239 : _GEN12644;
wire  _GEN12646 = io_x[26] ? _GEN12645 : _GEN12643;
wire  _GEN12647 = io_x[73] ? _GEN12646 : _GEN12640;
wire  _GEN12648 = io_x[33] ? _GEN12647 : _GEN12637;
wire  _GEN12649 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN12650 = io_x[73] ? _GEN10243 : _GEN12649;
wire  _GEN12651 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN12652 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12653 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12654 = io_x[30] ? _GEN12653 : _GEN10239;
wire  _GEN12655 = io_x[26] ? _GEN12654 : _GEN12652;
wire  _GEN12656 = io_x[73] ? _GEN12655 : _GEN12651;
wire  _GEN12657 = io_x[33] ? _GEN12656 : _GEN12650;
wire  _GEN12658 = io_x[28] ? _GEN12657 : _GEN12648;
wire  _GEN12659 = io_x[18] ? _GEN12658 : _GEN12630;
wire  _GEN12660 = io_x[25] ? _GEN12659 : _GEN12597;
wire  _GEN12661 = io_x[29] ? _GEN12660 : _GEN12571;
wire  _GEN12662 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12663 = io_x[30] ? _GEN12662 : _GEN10239;
wire  _GEN12664 = io_x[26] ? _GEN12663 : _GEN10241;
wire  _GEN12665 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12666 = io_x[30] ? _GEN12665 : _GEN10239;
wire  _GEN12667 = io_x[26] ? _GEN12666 : _GEN10241;
wire  _GEN12668 = io_x[73] ? _GEN12667 : _GEN12664;
wire  _GEN12669 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12670 = io_x[30] ? _GEN12669 : _GEN10239;
wire  _GEN12671 = io_x[26] ? _GEN12670 : _GEN10241;
wire  _GEN12672 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12673 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12674 = io_x[30] ? _GEN12673 : _GEN10239;
wire  _GEN12675 = io_x[26] ? _GEN12674 : _GEN12672;
wire  _GEN12676 = io_x[73] ? _GEN12675 : _GEN12671;
wire  _GEN12677 = io_x[33] ? _GEN12676 : _GEN12668;
wire  _GEN12678 = io_x[28] ? _GEN12677 : _GEN11021;
wire  _GEN12679 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12680 = io_x[30] ? _GEN12679 : _GEN10239;
wire  _GEN12681 = io_x[26] ? _GEN12680 : _GEN10246;
wire  _GEN12682 = io_x[73] ? _GEN10243 : _GEN12681;
wire  _GEN12683 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12684 = io_x[30] ? _GEN12683 : _GEN10238;
wire  _GEN12685 = io_x[26] ? _GEN12684 : _GEN10241;
wire  _GEN12686 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12687 = io_x[30] ? _GEN12686 : _GEN10239;
wire  _GEN12688 = io_x[26] ? _GEN12687 : _GEN10241;
wire  _GEN12689 = io_x[73] ? _GEN12688 : _GEN12685;
wire  _GEN12690 = io_x[33] ? _GEN12689 : _GEN12682;
wire  _GEN12691 = io_x[28] ? _GEN12690 : _GEN11021;
wire  _GEN12692 = io_x[18] ? _GEN12691 : _GEN12678;
wire  _GEN12693 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12694 = io_x[30] ? _GEN12693 : _GEN10239;
wire  _GEN12695 = io_x[26] ? _GEN10241 : _GEN12694;
wire  _GEN12696 = io_x[73] ? _GEN12695 : _GEN10243;
wire  _GEN12697 = io_x[33] ? _GEN10237 : _GEN12696;
wire  _GEN12698 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN12699 = io_x[73] ? _GEN12698 : _GEN10259;
wire  _GEN12700 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12701 = io_x[30] ? _GEN12700 : _GEN10239;
wire  _GEN12702 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12703 = io_x[30] ? _GEN12702 : _GEN10239;
wire  _GEN12704 = io_x[26] ? _GEN12703 : _GEN12701;
wire  _GEN12705 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12706 = io_x[30] ? _GEN12705 : _GEN10238;
wire  _GEN12707 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12708 = io_x[26] ? _GEN12707 : _GEN12706;
wire  _GEN12709 = io_x[73] ? _GEN12708 : _GEN12704;
wire  _GEN12710 = io_x[33] ? _GEN12709 : _GEN12699;
wire  _GEN12711 = io_x[28] ? _GEN12710 : _GEN12697;
wire  _GEN12712 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12713 = io_x[30] ? _GEN12712 : _GEN10239;
wire  _GEN12714 = io_x[26] ? _GEN12713 : _GEN10246;
wire  _GEN12715 = io_x[73] ? _GEN10243 : _GEN12714;
wire  _GEN12716 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12717 = io_x[30] ? _GEN12716 : _GEN10239;
wire  _GEN12718 = io_x[26] ? _GEN12717 : _GEN10241;
wire  _GEN12719 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12720 = io_x[30] ? _GEN12719 : _GEN10239;
wire  _GEN12721 = io_x[26] ? _GEN10241 : _GEN12720;
wire  _GEN12722 = io_x[73] ? _GEN12721 : _GEN12718;
wire  _GEN12723 = io_x[33] ? _GEN12722 : _GEN12715;
wire  _GEN12724 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12725 = io_x[30] ? _GEN12724 : _GEN10239;
wire  _GEN12726 = io_x[26] ? _GEN10241 : _GEN12725;
wire  _GEN12727 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN12728 = io_x[73] ? _GEN12727 : _GEN12726;
wire  _GEN12729 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12730 = io_x[30] ? _GEN12729 : _GEN10239;
wire  _GEN12731 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12732 = io_x[26] ? _GEN12731 : _GEN12730;
wire  _GEN12733 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12734 = io_x[30] ? _GEN12733 : _GEN10239;
wire  _GEN12735 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12736 = io_x[30] ? _GEN12735 : _GEN10239;
wire  _GEN12737 = io_x[26] ? _GEN12736 : _GEN12734;
wire  _GEN12738 = io_x[73] ? _GEN12737 : _GEN12732;
wire  _GEN12739 = io_x[33] ? _GEN12738 : _GEN12728;
wire  _GEN12740 = io_x[28] ? _GEN12739 : _GEN12723;
wire  _GEN12741 = io_x[18] ? _GEN12740 : _GEN12711;
wire  _GEN12742 = io_x[25] ? _GEN12741 : _GEN12692;
wire  _GEN12743 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12744 = io_x[30] ? _GEN10239 : _GEN12743;
wire  _GEN12745 = io_x[26] ? _GEN12744 : _GEN10241;
wire  _GEN12746 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12747 = io_x[30] ? _GEN10239 : _GEN12746;
wire  _GEN12748 = io_x[26] ? _GEN12747 : _GEN10241;
wire  _GEN12749 = io_x[73] ? _GEN12748 : _GEN12745;
wire  _GEN12750 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12751 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12752 = io_x[30] ? _GEN12751 : _GEN12750;
wire  _GEN12753 = io_x[26] ? _GEN12752 : _GEN10241;
wire  _GEN12754 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12755 = io_x[30] ? _GEN10239 : _GEN12754;
wire  _GEN12756 = io_x[26] ? _GEN12755 : _GEN10241;
wire  _GEN12757 = io_x[73] ? _GEN12756 : _GEN12753;
wire  _GEN12758 = io_x[33] ? _GEN12757 : _GEN12749;
wire  _GEN12759 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12760 = io_x[30] ? _GEN12759 : _GEN10239;
wire  _GEN12761 = io_x[26] ? _GEN10246 : _GEN12760;
wire  _GEN12762 = io_x[73] ? _GEN10259 : _GEN12761;
wire  _GEN12763 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN12764 = io_x[73] ? _GEN10259 : _GEN12763;
wire  _GEN12765 = io_x[33] ? _GEN12764 : _GEN12762;
wire  _GEN12766 = io_x[28] ? _GEN12765 : _GEN12758;
wire  _GEN12767 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12768 = io_x[30] ? _GEN10239 : _GEN12767;
wire  _GEN12769 = io_x[26] ? _GEN12768 : _GEN10241;
wire  _GEN12770 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN12771 = io_x[73] ? _GEN12770 : _GEN12769;
wire  _GEN12772 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12773 = io_x[30] ? _GEN10239 : _GEN12772;
wire  _GEN12774 = io_x[26] ? _GEN12773 : _GEN10246;
wire  _GEN12775 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN12776 = io_x[73] ? _GEN12775 : _GEN12774;
wire  _GEN12777 = io_x[33] ? _GEN12776 : _GEN12771;
wire  _GEN12778 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN12779 = io_x[73] ? _GEN12778 : _GEN10243;
wire  _GEN12780 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12781 = io_x[26] ? _GEN10241 : _GEN12780;
wire  _GEN12782 = io_x[73] ? _GEN12781 : _GEN10243;
wire  _GEN12783 = io_x[33] ? _GEN12782 : _GEN12779;
wire  _GEN12784 = io_x[28] ? _GEN12783 : _GEN12777;
wire  _GEN12785 = io_x[18] ? _GEN12784 : _GEN12766;
wire  _GEN12786 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12787 = io_x[30] ? _GEN12786 : _GEN10238;
wire  _GEN12788 = io_x[26] ? _GEN10241 : _GEN12787;
wire  _GEN12789 = io_x[73] ? _GEN12788 : _GEN10243;
wire  _GEN12790 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12791 = io_x[30] ? _GEN12790 : _GEN10239;
wire  _GEN12792 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12793 = io_x[30] ? _GEN10238 : _GEN12792;
wire  _GEN12794 = io_x[26] ? _GEN12793 : _GEN12791;
wire  _GEN12795 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12796 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12797 = io_x[30] ? _GEN12796 : _GEN12795;
wire  _GEN12798 = io_x[26] ? _GEN10241 : _GEN12797;
wire  _GEN12799 = io_x[73] ? _GEN12798 : _GEN12794;
wire  _GEN12800 = io_x[33] ? _GEN12799 : _GEN12789;
wire  _GEN12801 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12802 = io_x[30] ? _GEN12801 : _GEN10239;
wire  _GEN12803 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12804 = io_x[30] ? _GEN12803 : _GEN10239;
wire  _GEN12805 = io_x[26] ? _GEN12804 : _GEN12802;
wire  _GEN12806 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12807 = io_x[30] ? _GEN12806 : _GEN10239;
wire  _GEN12808 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12809 = io_x[30] ? _GEN12808 : _GEN10238;
wire  _GEN12810 = io_x[26] ? _GEN12809 : _GEN12807;
wire  _GEN12811 = io_x[73] ? _GEN12810 : _GEN12805;
wire  _GEN12812 = io_x[33] ? _GEN12811 : _GEN10237;
wire  _GEN12813 = io_x[28] ? _GEN12812 : _GEN12800;
wire  _GEN12814 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12815 = io_x[30] ? _GEN12814 : _GEN10239;
wire  _GEN12816 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12817 = io_x[30] ? _GEN10239 : _GEN12816;
wire  _GEN12818 = io_x[26] ? _GEN12817 : _GEN12815;
wire  _GEN12819 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12820 = io_x[26] ? _GEN10246 : _GEN12819;
wire  _GEN12821 = io_x[73] ? _GEN12820 : _GEN12818;
wire  _GEN12822 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12823 = io_x[30] ? _GEN12822 : _GEN10238;
wire  _GEN12824 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12825 = io_x[26] ? _GEN12824 : _GEN12823;
wire  _GEN12826 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12827 = io_x[30] ? _GEN12826 : _GEN10239;
wire  _GEN12828 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12829 = io_x[26] ? _GEN12828 : _GEN12827;
wire  _GEN12830 = io_x[73] ? _GEN12829 : _GEN12825;
wire  _GEN12831 = io_x[33] ? _GEN12830 : _GEN12821;
wire  _GEN12832 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12833 = io_x[30] ? _GEN10238 : _GEN12832;
wire  _GEN12834 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12835 = io_x[30] ? _GEN12834 : _GEN10239;
wire  _GEN12836 = io_x[26] ? _GEN12835 : _GEN12833;
wire  _GEN12837 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12838 = io_x[30] ? _GEN12837 : _GEN10239;
wire  _GEN12839 = io_x[26] ? _GEN12838 : _GEN10241;
wire  _GEN12840 = io_x[73] ? _GEN12839 : _GEN12836;
wire  _GEN12841 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12842 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12843 = io_x[30] ? _GEN12842 : _GEN12841;
wire  _GEN12844 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12845 = io_x[30] ? _GEN12844 : _GEN10238;
wire  _GEN12846 = io_x[26] ? _GEN12845 : _GEN12843;
wire  _GEN12847 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12848 = io_x[30] ? _GEN12847 : _GEN10239;
wire  _GEN12849 = io_x[26] ? _GEN12848 : _GEN10246;
wire  _GEN12850 = io_x[73] ? _GEN12849 : _GEN12846;
wire  _GEN12851 = io_x[33] ? _GEN12850 : _GEN12840;
wire  _GEN12852 = io_x[28] ? _GEN12851 : _GEN12831;
wire  _GEN12853 = io_x[18] ? _GEN12852 : _GEN12813;
wire  _GEN12854 = io_x[25] ? _GEN12853 : _GEN12785;
wire  _GEN12855 = io_x[29] ? _GEN12854 : _GEN12742;
wire  _GEN12856 = io_x[23] ? _GEN12855 : _GEN12661;
wire  _GEN12857 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12858 = io_x[30] ? _GEN12857 : _GEN10239;
wire  _GEN12859 = io_x[26] ? _GEN10241 : _GEN12858;
wire  _GEN12860 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12861 = io_x[30] ? _GEN12860 : _GEN10239;
wire  _GEN12862 = io_x[26] ? _GEN10241 : _GEN12861;
wire  _GEN12863 = io_x[73] ? _GEN12862 : _GEN12859;
wire  _GEN12864 = io_x[33] ? _GEN12863 : _GEN10237;
wire  _GEN12865 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12866 = io_x[30] ? _GEN10239 : _GEN12865;
wire  _GEN12867 = io_x[26] ? _GEN12866 : _GEN10241;
wire  _GEN12868 = io_x[73] ? _GEN10259 : _GEN12867;
wire  _GEN12869 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12870 = io_x[30] ? _GEN10239 : _GEN12869;
wire  _GEN12871 = io_x[26] ? _GEN12870 : _GEN10241;
wire  _GEN12872 = io_x[73] ? _GEN10259 : _GEN12871;
wire  _GEN12873 = io_x[33] ? _GEN12872 : _GEN12868;
wire  _GEN12874 = io_x[28] ? _GEN12873 : _GEN12864;
wire  _GEN12875 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12876 = io_x[30] ? _GEN12875 : _GEN10239;
wire  _GEN12877 = io_x[26] ? _GEN10241 : _GEN12876;
wire  _GEN12878 = io_x[73] ? _GEN10243 : _GEN12877;
wire  _GEN12879 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12880 = io_x[30] ? _GEN12879 : _GEN10239;
wire  _GEN12881 = io_x[26] ? _GEN10241 : _GEN12880;
wire  _GEN12882 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN12883 = io_x[73] ? _GEN12882 : _GEN12881;
wire  _GEN12884 = io_x[33] ? _GEN12883 : _GEN12878;
wire  _GEN12885 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12886 = io_x[30] ? _GEN10239 : _GEN12885;
wire  _GEN12887 = io_x[26] ? _GEN12886 : _GEN10241;
wire  _GEN12888 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12889 = io_x[26] ? _GEN12888 : _GEN10241;
wire  _GEN12890 = io_x[73] ? _GEN12889 : _GEN12887;
wire  _GEN12891 = io_x[33] ? _GEN12890 : _GEN10237;
wire  _GEN12892 = io_x[28] ? _GEN12891 : _GEN12884;
wire  _GEN12893 = io_x[18] ? _GEN12892 : _GEN12874;
wire  _GEN12894 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12895 = io_x[26] ? _GEN10241 : _GEN12894;
wire  _GEN12896 = io_x[73] ? _GEN12895 : _GEN10243;
wire  _GEN12897 = io_x[33] ? _GEN12896 : _GEN10237;
wire  _GEN12898 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12899 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12900 = io_x[26] ? _GEN12899 : _GEN12898;
wire  _GEN12901 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12902 = io_x[26] ? _GEN12901 : _GEN10246;
wire  _GEN12903 = io_x[73] ? _GEN12902 : _GEN12900;
wire  _GEN12904 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12905 = io_x[30] ? _GEN12904 : _GEN10239;
wire  _GEN12906 = io_x[26] ? _GEN12905 : _GEN10246;
wire  _GEN12907 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12908 = io_x[30] ? _GEN12907 : _GEN10238;
wire  _GEN12909 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12910 = io_x[26] ? _GEN12909 : _GEN12908;
wire  _GEN12911 = io_x[73] ? _GEN12910 : _GEN12906;
wire  _GEN12912 = io_x[33] ? _GEN12911 : _GEN12903;
wire  _GEN12913 = io_x[28] ? _GEN12912 : _GEN12897;
wire  _GEN12914 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12915 = io_x[30] ? _GEN12914 : _GEN10238;
wire  _GEN12916 = io_x[26] ? _GEN10241 : _GEN12915;
wire  _GEN12917 = io_x[73] ? _GEN12916 : _GEN10259;
wire  _GEN12918 = io_x[33] ? _GEN12917 : _GEN10306;
wire  _GEN12919 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12920 = io_x[30] ? _GEN12919 : _GEN10238;
wire  _GEN12921 = io_x[26] ? _GEN12920 : _GEN10241;
wire  _GEN12922 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12923 = io_x[26] ? _GEN10246 : _GEN12922;
wire  _GEN12924 = io_x[73] ? _GEN12923 : _GEN12921;
wire  _GEN12925 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12926 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12927 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12928 = io_x[30] ? _GEN12927 : _GEN12926;
wire  _GEN12929 = io_x[26] ? _GEN12928 : _GEN12925;
wire  _GEN12930 = io_x[73] ? _GEN10243 : _GEN12929;
wire  _GEN12931 = io_x[33] ? _GEN12930 : _GEN12924;
wire  _GEN12932 = io_x[28] ? _GEN12931 : _GEN12918;
wire  _GEN12933 = io_x[18] ? _GEN12932 : _GEN12913;
wire  _GEN12934 = io_x[25] ? _GEN12933 : _GEN12893;
wire  _GEN12935 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12936 = io_x[30] ? _GEN10238 : _GEN12935;
wire  _GEN12937 = io_x[26] ? _GEN12936 : _GEN10241;
wire  _GEN12938 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12939 = io_x[26] ? _GEN12938 : _GEN10246;
wire  _GEN12940 = io_x[73] ? _GEN12939 : _GEN12937;
wire  _GEN12941 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12942 = io_x[30] ? _GEN10238 : _GEN12941;
wire  _GEN12943 = io_x[26] ? _GEN12942 : _GEN10241;
wire  _GEN12944 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12945 = io_x[26] ? _GEN12944 : _GEN10246;
wire  _GEN12946 = io_x[73] ? _GEN12945 : _GEN12943;
wire  _GEN12947 = io_x[33] ? _GEN12946 : _GEN12940;
wire  _GEN12948 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12949 = io_x[30] ? _GEN10239 : _GEN12948;
wire  _GEN12950 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12951 = io_x[26] ? _GEN12950 : _GEN12949;
wire  _GEN12952 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12953 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12954 = io_x[30] ? _GEN12953 : _GEN12952;
wire  _GEN12955 = io_x[26] ? _GEN10241 : _GEN12954;
wire  _GEN12956 = io_x[73] ? _GEN12955 : _GEN12951;
wire  _GEN12957 = io_x[33] ? _GEN12956 : _GEN10306;
wire  _GEN12958 = io_x[28] ? _GEN12957 : _GEN12947;
wire  _GEN12959 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12960 = io_x[26] ? _GEN12959 : _GEN10241;
wire  _GEN12961 = io_x[73] ? _GEN10243 : _GEN12960;
wire  _GEN12962 = io_x[33] ? _GEN12961 : _GEN10306;
wire  _GEN12963 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12964 = io_x[30] ? _GEN10238 : _GEN12963;
wire  _GEN12965 = io_x[26] ? _GEN10246 : _GEN12964;
wire  _GEN12966 = io_x[73] ? _GEN10259 : _GEN12965;
wire  _GEN12967 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12968 = io_x[30] ? _GEN10238 : _GEN12967;
wire  _GEN12969 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN12970 = io_x[26] ? _GEN12969 : _GEN12968;
wire  _GEN12971 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12972 = io_x[30] ? _GEN12971 : _GEN10239;
wire  _GEN12973 = io_x[26] ? _GEN10246 : _GEN12972;
wire  _GEN12974 = io_x[73] ? _GEN12973 : _GEN12970;
wire  _GEN12975 = io_x[33] ? _GEN12974 : _GEN12966;
wire  _GEN12976 = io_x[28] ? _GEN12975 : _GEN12962;
wire  _GEN12977 = io_x[18] ? _GEN12976 : _GEN12958;
wire  _GEN12978 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12979 = io_x[26] ? _GEN10241 : _GEN12978;
wire  _GEN12980 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12981 = io_x[30] ? _GEN10239 : _GEN12980;
wire  _GEN12982 = io_x[26] ? _GEN12981 : _GEN10246;
wire  _GEN12983 = io_x[73] ? _GEN12982 : _GEN12979;
wire  _GEN12984 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN12985 = io_x[30] ? _GEN12984 : _GEN10239;
wire  _GEN12986 = io_x[26] ? _GEN12985 : _GEN10241;
wire  _GEN12987 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12988 = io_x[30] ? _GEN10238 : _GEN12987;
wire  _GEN12989 = io_x[26] ? _GEN12988 : _GEN10246;
wire  _GEN12990 = io_x[73] ? _GEN12989 : _GEN12986;
wire  _GEN12991 = io_x[33] ? _GEN12990 : _GEN12983;
wire  _GEN12992 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12993 = io_x[30] ? _GEN10239 : _GEN12992;
wire  _GEN12994 = io_x[26] ? _GEN12993 : _GEN10241;
wire  _GEN12995 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN12996 = io_x[26] ? _GEN12995 : _GEN10241;
wire  _GEN12997 = io_x[73] ? _GEN12996 : _GEN12994;
wire  _GEN12998 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN12999 = io_x[30] ? _GEN12998 : _GEN10238;
wire  _GEN13000 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13001 = io_x[30] ? _GEN13000 : _GEN10239;
wire  _GEN13002 = io_x[26] ? _GEN13001 : _GEN12999;
wire  _GEN13003 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN13004 = io_x[26] ? _GEN13003 : _GEN10241;
wire  _GEN13005 = io_x[73] ? _GEN13004 : _GEN13002;
wire  _GEN13006 = io_x[33] ? _GEN13005 : _GEN12997;
wire  _GEN13007 = io_x[28] ? _GEN13006 : _GEN12991;
wire  _GEN13008 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13009 = io_x[30] ? _GEN13008 : _GEN10238;
wire  _GEN13010 = io_x[26] ? _GEN13009 : _GEN10241;
wire  _GEN13011 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13012 = io_x[30] ? _GEN10239 : _GEN13011;
wire  _GEN13013 = io_x[26] ? _GEN10246 : _GEN13012;
wire  _GEN13014 = io_x[73] ? _GEN13013 : _GEN13010;
wire  _GEN13015 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13016 = io_x[30] ? _GEN13015 : _GEN10238;
wire  _GEN13017 = io_x[26] ? _GEN13016 : _GEN10246;
wire  _GEN13018 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13019 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13020 = io_x[30] ? _GEN13019 : _GEN13018;
wire  _GEN13021 = io_x[26] ? _GEN10246 : _GEN13020;
wire  _GEN13022 = io_x[73] ? _GEN13021 : _GEN13017;
wire  _GEN13023 = io_x[33] ? _GEN13022 : _GEN13014;
wire  _GEN13024 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN13025 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13026 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13027 = io_x[30] ? _GEN13026 : _GEN13025;
wire  _GEN13028 = io_x[26] ? _GEN13027 : _GEN13024;
wire  _GEN13029 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13030 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13031 = io_x[30] ? _GEN13030 : _GEN13029;
wire  _GEN13032 = io_x[26] ? _GEN13031 : _GEN10241;
wire  _GEN13033 = io_x[73] ? _GEN13032 : _GEN13028;
wire  _GEN13034 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN13035 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13036 = io_x[30] ? _GEN13035 : _GEN10239;
wire  _GEN13037 = io_x[26] ? _GEN13036 : _GEN13034;
wire  _GEN13038 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13039 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13040 = io_x[30] ? _GEN13039 : _GEN13038;
wire  _GEN13041 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13042 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13043 = io_x[30] ? _GEN13042 : _GEN13041;
wire  _GEN13044 = io_x[26] ? _GEN13043 : _GEN13040;
wire  _GEN13045 = io_x[73] ? _GEN13044 : _GEN13037;
wire  _GEN13046 = io_x[33] ? _GEN13045 : _GEN13033;
wire  _GEN13047 = io_x[28] ? _GEN13046 : _GEN13023;
wire  _GEN13048 = io_x[18] ? _GEN13047 : _GEN13007;
wire  _GEN13049 = io_x[25] ? _GEN13048 : _GEN12977;
wire  _GEN13050 = io_x[29] ? _GEN13049 : _GEN12934;
wire  _GEN13051 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13052 = io_x[30] ? _GEN13051 : _GEN10239;
wire  _GEN13053 = io_x[26] ? _GEN13052 : _GEN10241;
wire  _GEN13054 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN13055 = io_x[73] ? _GEN13054 : _GEN13053;
wire  _GEN13056 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13057 = io_x[30] ? _GEN13056 : _GEN10239;
wire  _GEN13058 = io_x[26] ? _GEN13057 : _GEN10246;
wire  _GEN13059 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13060 = io_x[30] ? _GEN13059 : _GEN10239;
wire  _GEN13061 = io_x[26] ? _GEN13060 : _GEN10246;
wire  _GEN13062 = io_x[73] ? _GEN13061 : _GEN13058;
wire  _GEN13063 = io_x[33] ? _GEN13062 : _GEN13055;
wire  _GEN13064 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13065 = io_x[30] ? _GEN13064 : _GEN10239;
wire  _GEN13066 = io_x[26] ? _GEN13065 : _GEN10246;
wire  _GEN13067 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13068 = io_x[30] ? _GEN13067 : _GEN10239;
wire  _GEN13069 = io_x[26] ? _GEN13068 : _GEN10241;
wire  _GEN13070 = io_x[73] ? _GEN13069 : _GEN13066;
wire  _GEN13071 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13072 = io_x[30] ? _GEN13071 : _GEN10238;
wire  _GEN13073 = io_x[26] ? _GEN13072 : _GEN10246;
wire  _GEN13074 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13075 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13076 = io_x[30] ? _GEN13075 : _GEN13074;
wire  _GEN13077 = io_x[26] ? _GEN13076 : _GEN10241;
wire  _GEN13078 = io_x[73] ? _GEN13077 : _GEN13073;
wire  _GEN13079 = io_x[33] ? _GEN13078 : _GEN13070;
wire  _GEN13080 = io_x[28] ? _GEN13079 : _GEN13063;
wire  _GEN13081 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13082 = io_x[30] ? _GEN13081 : _GEN10238;
wire  _GEN13083 = io_x[26] ? _GEN13082 : _GEN10246;
wire  _GEN13084 = io_x[73] ? _GEN13083 : _GEN10243;
wire  _GEN13085 = io_x[33] ? _GEN13084 : _GEN10306;
wire  _GEN13086 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13087 = io_x[30] ? _GEN13086 : _GEN10239;
wire  _GEN13088 = io_x[26] ? _GEN13087 : _GEN10241;
wire  _GEN13089 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN13090 = io_x[73] ? _GEN13089 : _GEN13088;
wire  _GEN13091 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13092 = io_x[30] ? _GEN10239 : _GEN13091;
wire  _GEN13093 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13094 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13095 = io_x[30] ? _GEN13094 : _GEN13093;
wire  _GEN13096 = io_x[26] ? _GEN13095 : _GEN13092;
wire  _GEN13097 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13098 = io_x[30] ? _GEN13097 : _GEN10238;
wire  _GEN13099 = io_x[26] ? _GEN13098 : _GEN10246;
wire  _GEN13100 = io_x[73] ? _GEN13099 : _GEN13096;
wire  _GEN13101 = io_x[33] ? _GEN13100 : _GEN13090;
wire  _GEN13102 = io_x[28] ? _GEN13101 : _GEN13085;
wire  _GEN13103 = io_x[18] ? _GEN13102 : _GEN13080;
wire  _GEN13104 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13105 = io_x[30] ? _GEN13104 : _GEN10238;
wire  _GEN13106 = io_x[26] ? _GEN10241 : _GEN13105;
wire  _GEN13107 = io_x[73] ? _GEN10243 : _GEN13106;
wire  _GEN13108 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13109 = io_x[30] ? _GEN13108 : _GEN10238;
wire  _GEN13110 = io_x[26] ? _GEN10241 : _GEN13109;
wire  _GEN13111 = io_x[73] ? _GEN10243 : _GEN13110;
wire  _GEN13112 = io_x[33] ? _GEN13111 : _GEN13107;
wire  _GEN13113 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13114 = io_x[30] ? _GEN10239 : _GEN13113;
wire  _GEN13115 = io_x[26] ? _GEN10246 : _GEN13114;
wire  _GEN13116 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13117 = io_x[30] ? _GEN13116 : _GEN10239;
wire  _GEN13118 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13119 = io_x[30] ? _GEN13118 : _GEN10238;
wire  _GEN13120 = io_x[26] ? _GEN13119 : _GEN13117;
wire  _GEN13121 = io_x[73] ? _GEN13120 : _GEN13115;
wire  _GEN13122 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN13123 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13124 = io_x[30] ? _GEN10238 : _GEN13123;
wire  _GEN13125 = io_x[26] ? _GEN13124 : _GEN13122;
wire  _GEN13126 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN13127 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN13128 = io_x[26] ? _GEN13127 : _GEN13126;
wire  _GEN13129 = io_x[73] ? _GEN13128 : _GEN13125;
wire  _GEN13130 = io_x[33] ? _GEN13129 : _GEN13121;
wire  _GEN13131 = io_x[28] ? _GEN13130 : _GEN13112;
wire  _GEN13132 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13133 = io_x[30] ? _GEN13132 : _GEN10239;
wire  _GEN13134 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13135 = io_x[30] ? _GEN13134 : _GEN10239;
wire  _GEN13136 = io_x[26] ? _GEN13135 : _GEN13133;
wire  _GEN13137 = io_x[73] ? _GEN10243 : _GEN13136;
wire  _GEN13138 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13139 = io_x[30] ? _GEN13138 : _GEN10239;
wire  _GEN13140 = io_x[30] ? _GEN10239 : _GEN10238;
wire  _GEN13141 = io_x[26] ? _GEN13140 : _GEN13139;
wire  _GEN13142 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13143 = io_x[30] ? _GEN13142 : _GEN10239;
wire  _GEN13144 = io_x[26] ? _GEN10246 : _GEN13143;
wire  _GEN13145 = io_x[73] ? _GEN13144 : _GEN13141;
wire  _GEN13146 = io_x[33] ? _GEN13145 : _GEN13137;
wire  _GEN13147 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13148 = io_x[30] ? _GEN13147 : _GEN10238;
wire  _GEN13149 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13150 = io_x[30] ? _GEN10239 : _GEN13149;
wire  _GEN13151 = io_x[26] ? _GEN13150 : _GEN13148;
wire  _GEN13152 = io_x[73] ? _GEN10259 : _GEN13151;
wire  _GEN13153 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13154 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13155 = io_x[30] ? _GEN13154 : _GEN13153;
wire  _GEN13156 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13157 = io_x[30] ? _GEN10239 : _GEN13156;
wire  _GEN13158 = io_x[26] ? _GEN13157 : _GEN13155;
wire  _GEN13159 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13160 = io_x[30] ? _GEN10238 : _GEN13159;
wire  _GEN13161 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13162 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13163 = io_x[30] ? _GEN13162 : _GEN13161;
wire  _GEN13164 = io_x[26] ? _GEN13163 : _GEN13160;
wire  _GEN13165 = io_x[73] ? _GEN13164 : _GEN13158;
wire  _GEN13166 = io_x[33] ? _GEN13165 : _GEN13152;
wire  _GEN13167 = io_x[28] ? _GEN13166 : _GEN13146;
wire  _GEN13168 = io_x[18] ? _GEN13167 : _GEN13131;
wire  _GEN13169 = io_x[25] ? _GEN13168 : _GEN13103;
wire  _GEN13170 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13171 = io_x[30] ? _GEN13170 : _GEN10238;
wire  _GEN13172 = io_x[26] ? _GEN13171 : _GEN10241;
wire  _GEN13173 = io_x[73] ? _GEN13172 : _GEN10259;
wire  _GEN13174 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13175 = io_x[30] ? _GEN13174 : _GEN10238;
wire  _GEN13176 = io_x[26] ? _GEN13175 : _GEN10241;
wire  _GEN13177 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13178 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13179 = io_x[30] ? _GEN13178 : _GEN13177;
wire  _GEN13180 = io_x[26] ? _GEN13179 : _GEN10246;
wire  _GEN13181 = io_x[73] ? _GEN13180 : _GEN13176;
wire  _GEN13182 = io_x[33] ? _GEN13181 : _GEN13173;
wire  _GEN13183 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13184 = io_x[30] ? _GEN10239 : _GEN13183;
wire  _GEN13185 = io_x[26] ? _GEN13184 : _GEN10241;
wire  _GEN13186 = io_x[73] ? _GEN13185 : _GEN10243;
wire  _GEN13187 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13188 = io_x[30] ? _GEN10238 : _GEN13187;
wire  _GEN13189 = io_x[26] ? _GEN13188 : _GEN10241;
wire  _GEN13190 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13191 = io_x[30] ? _GEN10239 : _GEN13190;
wire  _GEN13192 = io_x[26] ? _GEN13191 : _GEN10241;
wire  _GEN13193 = io_x[73] ? _GEN13192 : _GEN13189;
wire  _GEN13194 = io_x[33] ? _GEN13193 : _GEN13186;
wire  _GEN13195 = io_x[28] ? _GEN13194 : _GEN13182;
wire  _GEN13196 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13197 = io_x[30] ? _GEN13196 : _GEN10239;
wire  _GEN13198 = io_x[26] ? _GEN13197 : _GEN10241;
wire  _GEN13199 = io_x[26] ? _GEN10241 : _GEN10246;
wire  _GEN13200 = io_x[73] ? _GEN13199 : _GEN13198;
wire  _GEN13201 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13202 = io_x[30] ? _GEN10239 : _GEN13201;
wire  _GEN13203 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13204 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13205 = io_x[30] ? _GEN13204 : _GEN13203;
wire  _GEN13206 = io_x[26] ? _GEN13205 : _GEN13202;
wire  _GEN13207 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13208 = io_x[30] ? _GEN13207 : _GEN10239;
wire  _GEN13209 = io_x[26] ? _GEN13208 : _GEN10241;
wire  _GEN13210 = io_x[73] ? _GEN13209 : _GEN13206;
wire  _GEN13211 = io_x[33] ? _GEN13210 : _GEN13200;
wire  _GEN13212 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13213 = io_x[30] ? _GEN13212 : _GEN10239;
wire  _GEN13214 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13215 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13216 = io_x[30] ? _GEN13215 : _GEN13214;
wire  _GEN13217 = io_x[26] ? _GEN13216 : _GEN13213;
wire  _GEN13218 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13219 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13220 = io_x[30] ? _GEN13219 : _GEN13218;
wire  _GEN13221 = io_x[26] ? _GEN13220 : _GEN10241;
wire  _GEN13222 = io_x[73] ? _GEN13221 : _GEN13217;
wire  _GEN13223 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN13224 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13225 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13226 = io_x[30] ? _GEN13225 : _GEN13224;
wire  _GEN13227 = io_x[26] ? _GEN13226 : _GEN13223;
wire  _GEN13228 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13229 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13230 = io_x[30] ? _GEN13229 : _GEN13228;
wire  _GEN13231 = io_x[26] ? _GEN13230 : _GEN10246;
wire  _GEN13232 = io_x[73] ? _GEN13231 : _GEN13227;
wire  _GEN13233 = io_x[33] ? _GEN13232 : _GEN13222;
wire  _GEN13234 = io_x[28] ? _GEN13233 : _GEN13211;
wire  _GEN13235 = io_x[18] ? _GEN13234 : _GEN13195;
wire  _GEN13236 = io_x[30] ? _GEN10238 : _GEN10239;
wire  _GEN13237 = io_x[26] ? _GEN10246 : _GEN13236;
wire  _GEN13238 = io_x[73] ? _GEN13237 : _GEN10259;
wire  _GEN13239 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13240 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13241 = io_x[30] ? _GEN13240 : _GEN13239;
wire  _GEN13242 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13243 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13244 = io_x[30] ? _GEN13243 : _GEN13242;
wire  _GEN13245 = io_x[26] ? _GEN13244 : _GEN13241;
wire  _GEN13246 = io_x[26] ? _GEN10246 : _GEN10241;
wire  _GEN13247 = io_x[73] ? _GEN13246 : _GEN13245;
wire  _GEN13248 = io_x[33] ? _GEN13247 : _GEN13238;
wire  _GEN13249 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13250 = io_x[30] ? _GEN13249 : _GEN10239;
wire  _GEN13251 = io_x[26] ? _GEN13250 : _GEN10246;
wire  _GEN13252 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13253 = io_x[30] ? _GEN10239 : _GEN13252;
wire  _GEN13254 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13255 = io_x[30] ? _GEN13254 : _GEN10238;
wire  _GEN13256 = io_x[26] ? _GEN13255 : _GEN13253;
wire  _GEN13257 = io_x[73] ? _GEN13256 : _GEN13251;
wire  _GEN13258 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13259 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13260 = io_x[30] ? _GEN13259 : _GEN13258;
wire  _GEN13261 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13262 = io_x[30] ? _GEN13261 : _GEN10239;
wire  _GEN13263 = io_x[26] ? _GEN13262 : _GEN13260;
wire  _GEN13264 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13265 = io_x[30] ? _GEN10238 : _GEN13264;
wire  _GEN13266 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13267 = io_x[30] ? _GEN13266 : _GEN10238;
wire  _GEN13268 = io_x[26] ? _GEN13267 : _GEN13265;
wire  _GEN13269 = io_x[73] ? _GEN13268 : _GEN13263;
wire  _GEN13270 = io_x[33] ? _GEN13269 : _GEN13257;
wire  _GEN13271 = io_x[28] ? _GEN13270 : _GEN13248;
wire  _GEN13272 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13273 = io_x[30] ? _GEN13272 : _GEN10238;
wire  _GEN13274 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13275 = io_x[30] ? _GEN13274 : _GEN10239;
wire  _GEN13276 = io_x[26] ? _GEN13275 : _GEN13273;
wire  _GEN13277 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13278 = io_x[30] ? _GEN10238 : _GEN13277;
wire  _GEN13279 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13280 = io_x[30] ? _GEN10239 : _GEN13279;
wire  _GEN13281 = io_x[26] ? _GEN13280 : _GEN13278;
wire  _GEN13282 = io_x[73] ? _GEN13281 : _GEN13276;
wire  _GEN13283 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13284 = io_x[30] ? _GEN10239 : _GEN13283;
wire  _GEN13285 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13286 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13287 = io_x[30] ? _GEN13286 : _GEN13285;
wire  _GEN13288 = io_x[26] ? _GEN13287 : _GEN13284;
wire  _GEN13289 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13290 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13291 = io_x[30] ? _GEN13290 : _GEN13289;
wire  _GEN13292 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13293 = io_x[30] ? _GEN13292 : _GEN10239;
wire  _GEN13294 = io_x[26] ? _GEN13293 : _GEN13291;
wire  _GEN13295 = io_x[73] ? _GEN13294 : _GEN13288;
wire  _GEN13296 = io_x[33] ? _GEN13295 : _GEN13282;
wire  _GEN13297 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13298 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13299 = io_x[30] ? _GEN13298 : _GEN13297;
wire  _GEN13300 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13301 = io_x[30] ? _GEN13300 : _GEN10238;
wire  _GEN13302 = io_x[26] ? _GEN13301 : _GEN13299;
wire  _GEN13303 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13304 = io_x[30] ? _GEN10238 : _GEN13303;
wire  _GEN13305 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13306 = io_x[30] ? _GEN13305 : _GEN10238;
wire  _GEN13307 = io_x[26] ? _GEN13306 : _GEN13304;
wire  _GEN13308 = io_x[73] ? _GEN13307 : _GEN13302;
wire  _GEN13309 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13310 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13311 = io_x[30] ? _GEN13310 : _GEN13309;
wire  _GEN13312 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13313 = io_x[30] ? _GEN13312 : _GEN10238;
wire  _GEN13314 = io_x[26] ? _GEN13313 : _GEN13311;
wire  _GEN13315 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13316 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13317 = io_x[30] ? _GEN13316 : _GEN13315;
wire  _GEN13318 = io_x[22] ? _GEN10247 : _GEN10248;
wire  _GEN13319 = io_x[22] ? _GEN10248 : _GEN10247;
wire  _GEN13320 = io_x[30] ? _GEN13319 : _GEN13318;
wire  _GEN13321 = io_x[26] ? _GEN13320 : _GEN13317;
wire  _GEN13322 = io_x[73] ? _GEN13321 : _GEN13314;
wire  _GEN13323 = io_x[33] ? _GEN13322 : _GEN13308;
wire  _GEN13324 = io_x[28] ? _GEN13323 : _GEN13296;
wire  _GEN13325 = io_x[18] ? _GEN13324 : _GEN13271;
wire  _GEN13326 = io_x[25] ? _GEN13325 : _GEN13235;
wire  _GEN13327 = io_x[29] ? _GEN13326 : _GEN13169;
wire  _GEN13328 = io_x[23] ? _GEN13327 : _GEN13050;
wire  _GEN13329 = io_x[31] ? _GEN13328 : _GEN12856;
wire  _GEN13330 = io_x[19] ? _GEN13329 : _GEN12503;
wire  _GEN13331 = io_x[76] ? _GEN13330 : _GEN11892;
assign io_y[8] = _GEN13331;
wire  _GEN13332 = 1'b0;
wire  _GEN13333 = 1'b1;
wire  _GEN13334 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13335 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13336 = io_x[25] ? _GEN13335 : _GEN13334;
wire  _GEN13337 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13338 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13339 = io_x[25] ? _GEN13338 : _GEN13337;
wire  _GEN13340 = io_x[73] ? _GEN13339 : _GEN13336;
wire  _GEN13341 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13342 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13343 = io_x[25] ? _GEN13342 : _GEN13341;
wire  _GEN13344 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13345 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13346 = io_x[25] ? _GEN13345 : _GEN13344;
wire  _GEN13347 = io_x[73] ? _GEN13346 : _GEN13343;
wire  _GEN13348 = io_x[75] ? _GEN13347 : _GEN13340;
wire  _GEN13349 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13350 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13351 = io_x[25] ? _GEN13350 : _GEN13349;
wire  _GEN13352 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13353 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13354 = io_x[25] ? _GEN13353 : _GEN13352;
wire  _GEN13355 = io_x[73] ? _GEN13354 : _GEN13351;
wire  _GEN13356 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13357 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13358 = io_x[25] ? _GEN13357 : _GEN13356;
wire  _GEN13359 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13360 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13361 = io_x[25] ? _GEN13360 : _GEN13359;
wire  _GEN13362 = io_x[73] ? _GEN13361 : _GEN13358;
wire  _GEN13363 = io_x[75] ? _GEN13362 : _GEN13355;
wire  _GEN13364 = io_x[21] ? _GEN13363 : _GEN13348;
wire  _GEN13365 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13366 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13367 = io_x[25] ? _GEN13366 : _GEN13365;
wire  _GEN13368 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13369 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13370 = io_x[25] ? _GEN13369 : _GEN13368;
wire  _GEN13371 = io_x[73] ? _GEN13370 : _GEN13367;
wire  _GEN13372 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13373 = 1'b1;
wire  _GEN13374 = io_x[25] ? _GEN13373 : _GEN13372;
wire  _GEN13375 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13376 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13377 = io_x[25] ? _GEN13376 : _GEN13375;
wire  _GEN13378 = io_x[73] ? _GEN13377 : _GEN13374;
wire  _GEN13379 = io_x[75] ? _GEN13378 : _GEN13371;
wire  _GEN13380 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13381 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13382 = io_x[25] ? _GEN13381 : _GEN13380;
wire  _GEN13383 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13384 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13385 = io_x[25] ? _GEN13384 : _GEN13383;
wire  _GEN13386 = io_x[73] ? _GEN13385 : _GEN13382;
wire  _GEN13387 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13388 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13389 = io_x[25] ? _GEN13388 : _GEN13387;
wire  _GEN13390 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13391 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13392 = io_x[25] ? _GEN13391 : _GEN13390;
wire  _GEN13393 = io_x[73] ? _GEN13392 : _GEN13389;
wire  _GEN13394 = io_x[75] ? _GEN13393 : _GEN13386;
wire  _GEN13395 = io_x[21] ? _GEN13394 : _GEN13379;
wire  _GEN13396 = io_x[71] ? _GEN13395 : _GEN13364;
wire  _GEN13397 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13398 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13399 = io_x[25] ? _GEN13398 : _GEN13397;
wire  _GEN13400 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13401 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13402 = io_x[25] ? _GEN13401 : _GEN13400;
wire  _GEN13403 = io_x[73] ? _GEN13402 : _GEN13399;
wire  _GEN13404 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13405 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13406 = io_x[25] ? _GEN13405 : _GEN13404;
wire  _GEN13407 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13408 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13409 = io_x[25] ? _GEN13408 : _GEN13407;
wire  _GEN13410 = io_x[73] ? _GEN13409 : _GEN13406;
wire  _GEN13411 = io_x[75] ? _GEN13410 : _GEN13403;
wire  _GEN13412 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13413 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13414 = io_x[25] ? _GEN13413 : _GEN13412;
wire  _GEN13415 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13416 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13417 = io_x[25] ? _GEN13416 : _GEN13415;
wire  _GEN13418 = io_x[73] ? _GEN13417 : _GEN13414;
wire  _GEN13419 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13420 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13421 = io_x[25] ? _GEN13420 : _GEN13419;
wire  _GEN13422 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13423 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13424 = io_x[25] ? _GEN13423 : _GEN13422;
wire  _GEN13425 = io_x[73] ? _GEN13424 : _GEN13421;
wire  _GEN13426 = io_x[75] ? _GEN13425 : _GEN13418;
wire  _GEN13427 = io_x[21] ? _GEN13426 : _GEN13411;
wire  _GEN13428 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13429 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13430 = io_x[25] ? _GEN13429 : _GEN13428;
wire  _GEN13431 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13432 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13433 = io_x[25] ? _GEN13432 : _GEN13431;
wire  _GEN13434 = io_x[73] ? _GEN13433 : _GEN13430;
wire  _GEN13435 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13436 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13437 = io_x[25] ? _GEN13436 : _GEN13435;
wire  _GEN13438 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13439 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13440 = io_x[25] ? _GEN13439 : _GEN13438;
wire  _GEN13441 = io_x[73] ? _GEN13440 : _GEN13437;
wire  _GEN13442 = io_x[75] ? _GEN13441 : _GEN13434;
wire  _GEN13443 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13444 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13445 = io_x[25] ? _GEN13444 : _GEN13443;
wire  _GEN13446 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13447 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13448 = io_x[25] ? _GEN13447 : _GEN13446;
wire  _GEN13449 = io_x[73] ? _GEN13448 : _GEN13445;
wire  _GEN13450 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13451 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13452 = io_x[25] ? _GEN13451 : _GEN13450;
wire  _GEN13453 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13454 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13455 = io_x[25] ? _GEN13454 : _GEN13453;
wire  _GEN13456 = io_x[73] ? _GEN13455 : _GEN13452;
wire  _GEN13457 = io_x[75] ? _GEN13456 : _GEN13449;
wire  _GEN13458 = io_x[21] ? _GEN13457 : _GEN13442;
wire  _GEN13459 = io_x[71] ? _GEN13458 : _GEN13427;
wire  _GEN13460 = io_x[29] ? _GEN13459 : _GEN13396;
wire  _GEN13461 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13462 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13463 = io_x[25] ? _GEN13462 : _GEN13461;
wire  _GEN13464 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13465 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13466 = io_x[25] ? _GEN13465 : _GEN13464;
wire  _GEN13467 = io_x[73] ? _GEN13466 : _GEN13463;
wire  _GEN13468 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13469 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13470 = io_x[25] ? _GEN13469 : _GEN13468;
wire  _GEN13471 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13472 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13473 = io_x[25] ? _GEN13472 : _GEN13471;
wire  _GEN13474 = io_x[73] ? _GEN13473 : _GEN13470;
wire  _GEN13475 = io_x[75] ? _GEN13474 : _GEN13467;
wire  _GEN13476 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13477 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13478 = io_x[25] ? _GEN13477 : _GEN13476;
wire  _GEN13479 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13480 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13481 = io_x[25] ? _GEN13480 : _GEN13479;
wire  _GEN13482 = io_x[73] ? _GEN13481 : _GEN13478;
wire  _GEN13483 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13484 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13485 = io_x[25] ? _GEN13484 : _GEN13483;
wire  _GEN13486 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13487 = io_x[25] ? _GEN13486 : _GEN13373;
wire  _GEN13488 = io_x[73] ? _GEN13487 : _GEN13485;
wire  _GEN13489 = io_x[75] ? _GEN13488 : _GEN13482;
wire  _GEN13490 = io_x[21] ? _GEN13489 : _GEN13475;
wire  _GEN13491 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13492 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13493 = io_x[25] ? _GEN13492 : _GEN13491;
wire  _GEN13494 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13495 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13496 = io_x[25] ? _GEN13495 : _GEN13494;
wire  _GEN13497 = io_x[73] ? _GEN13496 : _GEN13493;
wire  _GEN13498 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13499 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13500 = io_x[25] ? _GEN13499 : _GEN13498;
wire  _GEN13501 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13502 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13503 = io_x[25] ? _GEN13502 : _GEN13501;
wire  _GEN13504 = io_x[73] ? _GEN13503 : _GEN13500;
wire  _GEN13505 = io_x[75] ? _GEN13504 : _GEN13497;
wire  _GEN13506 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13507 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13508 = io_x[25] ? _GEN13507 : _GEN13506;
wire  _GEN13509 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13510 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13511 = io_x[25] ? _GEN13510 : _GEN13509;
wire  _GEN13512 = io_x[73] ? _GEN13511 : _GEN13508;
wire  _GEN13513 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13514 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13515 = io_x[25] ? _GEN13514 : _GEN13513;
wire  _GEN13516 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13517 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13518 = io_x[25] ? _GEN13517 : _GEN13516;
wire  _GEN13519 = io_x[73] ? _GEN13518 : _GEN13515;
wire  _GEN13520 = io_x[75] ? _GEN13519 : _GEN13512;
wire  _GEN13521 = io_x[21] ? _GEN13520 : _GEN13505;
wire  _GEN13522 = io_x[71] ? _GEN13521 : _GEN13490;
wire  _GEN13523 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13524 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13525 = io_x[25] ? _GEN13524 : _GEN13523;
wire  _GEN13526 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13527 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13528 = io_x[25] ? _GEN13527 : _GEN13526;
wire  _GEN13529 = io_x[73] ? _GEN13528 : _GEN13525;
wire  _GEN13530 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13531 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13532 = io_x[25] ? _GEN13531 : _GEN13530;
wire  _GEN13533 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13534 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13535 = io_x[25] ? _GEN13534 : _GEN13533;
wire  _GEN13536 = io_x[73] ? _GEN13535 : _GEN13532;
wire  _GEN13537 = io_x[75] ? _GEN13536 : _GEN13529;
wire  _GEN13538 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13539 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13540 = io_x[25] ? _GEN13539 : _GEN13538;
wire  _GEN13541 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13542 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13543 = io_x[25] ? _GEN13542 : _GEN13541;
wire  _GEN13544 = io_x[73] ? _GEN13543 : _GEN13540;
wire  _GEN13545 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13546 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13547 = io_x[25] ? _GEN13546 : _GEN13545;
wire  _GEN13548 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13549 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13550 = io_x[25] ? _GEN13549 : _GEN13548;
wire  _GEN13551 = io_x[73] ? _GEN13550 : _GEN13547;
wire  _GEN13552 = io_x[75] ? _GEN13551 : _GEN13544;
wire  _GEN13553 = io_x[21] ? _GEN13552 : _GEN13537;
wire  _GEN13554 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13555 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13556 = io_x[25] ? _GEN13555 : _GEN13554;
wire  _GEN13557 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13558 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13559 = io_x[25] ? _GEN13558 : _GEN13557;
wire  _GEN13560 = io_x[73] ? _GEN13559 : _GEN13556;
wire  _GEN13561 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13562 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13563 = io_x[25] ? _GEN13562 : _GEN13561;
wire  _GEN13564 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13565 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13566 = io_x[25] ? _GEN13565 : _GEN13564;
wire  _GEN13567 = io_x[73] ? _GEN13566 : _GEN13563;
wire  _GEN13568 = io_x[75] ? _GEN13567 : _GEN13560;
wire  _GEN13569 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13570 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13571 = io_x[25] ? _GEN13570 : _GEN13569;
wire  _GEN13572 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13573 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13574 = io_x[25] ? _GEN13573 : _GEN13572;
wire  _GEN13575 = io_x[73] ? _GEN13574 : _GEN13571;
wire  _GEN13576 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13577 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13578 = io_x[25] ? _GEN13577 : _GEN13576;
wire  _GEN13579 = io_x[17] ? _GEN13332 : _GEN13333;
wire  _GEN13580 = io_x[17] ? _GEN13333 : _GEN13332;
wire  _GEN13581 = io_x[25] ? _GEN13580 : _GEN13579;
wire  _GEN13582 = io_x[73] ? _GEN13581 : _GEN13578;
wire  _GEN13583 = io_x[75] ? _GEN13582 : _GEN13575;
wire  _GEN13584 = io_x[21] ? _GEN13583 : _GEN13568;
wire  _GEN13585 = io_x[71] ? _GEN13584 : _GEN13553;
wire  _GEN13586 = io_x[29] ? _GEN13585 : _GEN13522;
wire  _GEN13587 = io_x[79] ? _GEN13586 : _GEN13460;
assign io_y[7] = _GEN13587;
wire  _GEN13588 = 1'b0;
wire  _GEN13589 = 1'b1;
wire  _GEN13590 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13591 = 1'b0;
wire  _GEN13592 = io_x[24] ? _GEN13591 : _GEN13590;
wire  _GEN13593 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13594 = io_x[24] ? _GEN13593 : _GEN13591;
wire  _GEN13595 = io_x[74] ? _GEN13594 : _GEN13592;
wire  _GEN13596 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13597 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13598 = io_x[24] ? _GEN13597 : _GEN13596;
wire  _GEN13599 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13600 = io_x[24] ? _GEN13599 : _GEN13591;
wire  _GEN13601 = io_x[74] ? _GEN13600 : _GEN13598;
wire  _GEN13602 = io_x[19] ? _GEN13601 : _GEN13595;
wire  _GEN13603 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13604 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13605 = io_x[24] ? _GEN13604 : _GEN13603;
wire  _GEN13606 = 1'b1;
wire  _GEN13607 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13608 = io_x[24] ? _GEN13607 : _GEN13606;
wire  _GEN13609 = io_x[74] ? _GEN13608 : _GEN13605;
wire  _GEN13610 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13611 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13612 = io_x[24] ? _GEN13611 : _GEN13610;
wire  _GEN13613 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13614 = io_x[24] ? _GEN13613 : _GEN13606;
wire  _GEN13615 = io_x[74] ? _GEN13614 : _GEN13612;
wire  _GEN13616 = io_x[19] ? _GEN13615 : _GEN13609;
wire  _GEN13617 = io_x[21] ? _GEN13616 : _GEN13602;
wire  _GEN13618 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13619 = io_x[24] ? _GEN13591 : _GEN13618;
wire  _GEN13620 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13621 = io_x[24] ? _GEN13606 : _GEN13620;
wire  _GEN13622 = io_x[74] ? _GEN13621 : _GEN13619;
wire  _GEN13623 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13624 = io_x[24] ? _GEN13623 : _GEN13591;
wire  _GEN13625 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13626 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13627 = io_x[24] ? _GEN13626 : _GEN13625;
wire  _GEN13628 = io_x[74] ? _GEN13627 : _GEN13624;
wire  _GEN13629 = io_x[19] ? _GEN13628 : _GEN13622;
wire  _GEN13630 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13631 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13632 = io_x[24] ? _GEN13631 : _GEN13630;
wire  _GEN13633 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13634 = io_x[24] ? _GEN13591 : _GEN13633;
wire  _GEN13635 = io_x[74] ? _GEN13634 : _GEN13632;
wire  _GEN13636 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13637 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13638 = io_x[24] ? _GEN13637 : _GEN13636;
wire  _GEN13639 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13640 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13641 = io_x[24] ? _GEN13640 : _GEN13639;
wire  _GEN13642 = io_x[74] ? _GEN13641 : _GEN13638;
wire  _GEN13643 = io_x[19] ? _GEN13642 : _GEN13635;
wire  _GEN13644 = io_x[21] ? _GEN13643 : _GEN13629;
wire  _GEN13645 = io_x[23] ? _GEN13644 : _GEN13617;
wire  _GEN13646 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13647 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13648 = io_x[24] ? _GEN13647 : _GEN13646;
wire  _GEN13649 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13650 = io_x[24] ? _GEN13606 : _GEN13649;
wire  _GEN13651 = io_x[74] ? _GEN13650 : _GEN13648;
wire  _GEN13652 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13653 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13654 = io_x[24] ? _GEN13653 : _GEN13652;
wire  _GEN13655 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13656 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13657 = io_x[24] ? _GEN13656 : _GEN13655;
wire  _GEN13658 = io_x[74] ? _GEN13657 : _GEN13654;
wire  _GEN13659 = io_x[19] ? _GEN13658 : _GEN13651;
wire  _GEN13660 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13661 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13662 = io_x[24] ? _GEN13661 : _GEN13660;
wire  _GEN13663 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13664 = io_x[24] ? _GEN13663 : _GEN13606;
wire  _GEN13665 = io_x[74] ? _GEN13664 : _GEN13662;
wire  _GEN13666 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13667 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13668 = io_x[24] ? _GEN13667 : _GEN13666;
wire  _GEN13669 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13670 = io_x[24] ? _GEN13669 : _GEN13606;
wire  _GEN13671 = io_x[74] ? _GEN13670 : _GEN13668;
wire  _GEN13672 = io_x[19] ? _GEN13671 : _GEN13665;
wire  _GEN13673 = io_x[21] ? _GEN13672 : _GEN13659;
wire  _GEN13674 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13675 = io_x[24] ? _GEN13674 : _GEN13591;
wire  _GEN13676 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13677 = io_x[24] ? _GEN13606 : _GEN13676;
wire  _GEN13678 = io_x[74] ? _GEN13677 : _GEN13675;
wire  _GEN13679 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13680 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13681 = io_x[24] ? _GEN13680 : _GEN13679;
wire  _GEN13682 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13683 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13684 = io_x[24] ? _GEN13683 : _GEN13682;
wire  _GEN13685 = io_x[74] ? _GEN13684 : _GEN13681;
wire  _GEN13686 = io_x[19] ? _GEN13685 : _GEN13678;
wire  _GEN13687 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13688 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13689 = io_x[24] ? _GEN13688 : _GEN13687;
wire  _GEN13690 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13691 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13692 = io_x[24] ? _GEN13691 : _GEN13690;
wire  _GEN13693 = io_x[74] ? _GEN13692 : _GEN13689;
wire  _GEN13694 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13695 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13696 = io_x[24] ? _GEN13695 : _GEN13694;
wire  _GEN13697 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13698 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13699 = io_x[24] ? _GEN13698 : _GEN13697;
wire  _GEN13700 = io_x[74] ? _GEN13699 : _GEN13696;
wire  _GEN13701 = io_x[19] ? _GEN13700 : _GEN13693;
wire  _GEN13702 = io_x[21] ? _GEN13701 : _GEN13686;
wire  _GEN13703 = io_x[23] ? _GEN13702 : _GEN13673;
wire  _GEN13704 = io_x[25] ? _GEN13703 : _GEN13645;
wire  _GEN13705 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13706 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13707 = io_x[24] ? _GEN13706 : _GEN13705;
wire  _GEN13708 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13709 = io_x[24] ? _GEN13591 : _GEN13708;
wire  _GEN13710 = io_x[74] ? _GEN13709 : _GEN13707;
wire  _GEN13711 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13712 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13713 = io_x[24] ? _GEN13712 : _GEN13711;
wire  _GEN13714 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13715 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13716 = io_x[24] ? _GEN13715 : _GEN13714;
wire  _GEN13717 = io_x[74] ? _GEN13716 : _GEN13713;
wire  _GEN13718 = io_x[19] ? _GEN13717 : _GEN13710;
wire  _GEN13719 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13720 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13721 = io_x[24] ? _GEN13720 : _GEN13719;
wire  _GEN13722 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13723 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13724 = io_x[24] ? _GEN13723 : _GEN13722;
wire  _GEN13725 = io_x[74] ? _GEN13724 : _GEN13721;
wire  _GEN13726 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13727 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13728 = io_x[24] ? _GEN13727 : _GEN13726;
wire  _GEN13729 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13730 = io_x[24] ? _GEN13729 : _GEN13606;
wire  _GEN13731 = io_x[74] ? _GEN13730 : _GEN13728;
wire  _GEN13732 = io_x[19] ? _GEN13731 : _GEN13725;
wire  _GEN13733 = io_x[21] ? _GEN13732 : _GEN13718;
wire  _GEN13734 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13735 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13736 = io_x[24] ? _GEN13735 : _GEN13734;
wire  _GEN13737 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13738 = io_x[24] ? _GEN13591 : _GEN13737;
wire  _GEN13739 = io_x[74] ? _GEN13738 : _GEN13736;
wire  _GEN13740 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13741 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13742 = io_x[24] ? _GEN13741 : _GEN13740;
wire  _GEN13743 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13744 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13745 = io_x[24] ? _GEN13744 : _GEN13743;
wire  _GEN13746 = io_x[74] ? _GEN13745 : _GEN13742;
wire  _GEN13747 = io_x[19] ? _GEN13746 : _GEN13739;
wire  _GEN13748 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13749 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13750 = io_x[24] ? _GEN13749 : _GEN13748;
wire  _GEN13751 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13752 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13753 = io_x[24] ? _GEN13752 : _GEN13751;
wire  _GEN13754 = io_x[74] ? _GEN13753 : _GEN13750;
wire  _GEN13755 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13756 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13757 = io_x[24] ? _GEN13756 : _GEN13755;
wire  _GEN13758 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13759 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13760 = io_x[24] ? _GEN13759 : _GEN13758;
wire  _GEN13761 = io_x[74] ? _GEN13760 : _GEN13757;
wire  _GEN13762 = io_x[19] ? _GEN13761 : _GEN13754;
wire  _GEN13763 = io_x[21] ? _GEN13762 : _GEN13747;
wire  _GEN13764 = io_x[23] ? _GEN13763 : _GEN13733;
wire  _GEN13765 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13766 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13767 = io_x[24] ? _GEN13766 : _GEN13765;
wire  _GEN13768 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13769 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13770 = io_x[24] ? _GEN13769 : _GEN13768;
wire  _GEN13771 = io_x[74] ? _GEN13770 : _GEN13767;
wire  _GEN13772 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13773 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13774 = io_x[24] ? _GEN13773 : _GEN13772;
wire  _GEN13775 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13776 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13777 = io_x[24] ? _GEN13776 : _GEN13775;
wire  _GEN13778 = io_x[74] ? _GEN13777 : _GEN13774;
wire  _GEN13779 = io_x[19] ? _GEN13778 : _GEN13771;
wire  _GEN13780 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13781 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13782 = io_x[24] ? _GEN13781 : _GEN13780;
wire  _GEN13783 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13784 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13785 = io_x[24] ? _GEN13784 : _GEN13783;
wire  _GEN13786 = io_x[74] ? _GEN13785 : _GEN13782;
wire  _GEN13787 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13788 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13789 = io_x[24] ? _GEN13788 : _GEN13787;
wire  _GEN13790 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13791 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13792 = io_x[24] ? _GEN13791 : _GEN13790;
wire  _GEN13793 = io_x[74] ? _GEN13792 : _GEN13789;
wire  _GEN13794 = io_x[19] ? _GEN13793 : _GEN13786;
wire  _GEN13795 = io_x[21] ? _GEN13794 : _GEN13779;
wire  _GEN13796 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13797 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13798 = io_x[24] ? _GEN13797 : _GEN13796;
wire  _GEN13799 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13800 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13801 = io_x[24] ? _GEN13800 : _GEN13799;
wire  _GEN13802 = io_x[74] ? _GEN13801 : _GEN13798;
wire  _GEN13803 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13804 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13805 = io_x[24] ? _GEN13804 : _GEN13803;
wire  _GEN13806 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13807 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13808 = io_x[24] ? _GEN13807 : _GEN13806;
wire  _GEN13809 = io_x[74] ? _GEN13808 : _GEN13805;
wire  _GEN13810 = io_x[19] ? _GEN13809 : _GEN13802;
wire  _GEN13811 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13812 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13813 = io_x[24] ? _GEN13812 : _GEN13811;
wire  _GEN13814 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13815 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13816 = io_x[24] ? _GEN13815 : _GEN13814;
wire  _GEN13817 = io_x[74] ? _GEN13816 : _GEN13813;
wire  _GEN13818 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13819 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13820 = io_x[24] ? _GEN13819 : _GEN13818;
wire  _GEN13821 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13822 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13823 = io_x[24] ? _GEN13822 : _GEN13821;
wire  _GEN13824 = io_x[74] ? _GEN13823 : _GEN13820;
wire  _GEN13825 = io_x[19] ? _GEN13824 : _GEN13817;
wire  _GEN13826 = io_x[21] ? _GEN13825 : _GEN13810;
wire  _GEN13827 = io_x[23] ? _GEN13826 : _GEN13795;
wire  _GEN13828 = io_x[25] ? _GEN13827 : _GEN13764;
wire  _GEN13829 = io_x[16] ? _GEN13828 : _GEN13704;
wire  _GEN13830 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13831 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13832 = io_x[24] ? _GEN13831 : _GEN13830;
wire  _GEN13833 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13834 = io_x[24] ? _GEN13833 : _GEN13606;
wire  _GEN13835 = io_x[74] ? _GEN13834 : _GEN13832;
wire  _GEN13836 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13837 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13838 = io_x[24] ? _GEN13837 : _GEN13836;
wire  _GEN13839 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13840 = io_x[24] ? _GEN13839 : _GEN13606;
wire  _GEN13841 = io_x[74] ? _GEN13840 : _GEN13838;
wire  _GEN13842 = io_x[19] ? _GEN13841 : _GEN13835;
wire  _GEN13843 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13844 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13845 = io_x[24] ? _GEN13844 : _GEN13843;
wire  _GEN13846 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13847 = io_x[24] ? _GEN13846 : _GEN13606;
wire  _GEN13848 = io_x[74] ? _GEN13847 : _GEN13845;
wire  _GEN13849 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13850 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13851 = io_x[24] ? _GEN13850 : _GEN13849;
wire  _GEN13852 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13853 = io_x[24] ? _GEN13852 : _GEN13606;
wire  _GEN13854 = io_x[74] ? _GEN13853 : _GEN13851;
wire  _GEN13855 = io_x[19] ? _GEN13854 : _GEN13848;
wire  _GEN13856 = io_x[21] ? _GEN13855 : _GEN13842;
wire  _GEN13857 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13858 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13859 = io_x[24] ? _GEN13858 : _GEN13857;
wire  _GEN13860 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13861 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13862 = io_x[24] ? _GEN13861 : _GEN13860;
wire  _GEN13863 = io_x[74] ? _GEN13862 : _GEN13859;
wire  _GEN13864 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13865 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13866 = io_x[24] ? _GEN13865 : _GEN13864;
wire  _GEN13867 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13868 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13869 = io_x[24] ? _GEN13868 : _GEN13867;
wire  _GEN13870 = io_x[74] ? _GEN13869 : _GEN13866;
wire  _GEN13871 = io_x[19] ? _GEN13870 : _GEN13863;
wire  _GEN13872 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13873 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13874 = io_x[24] ? _GEN13873 : _GEN13872;
wire  _GEN13875 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13876 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13877 = io_x[24] ? _GEN13876 : _GEN13875;
wire  _GEN13878 = io_x[74] ? _GEN13877 : _GEN13874;
wire  _GEN13879 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13880 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13881 = io_x[24] ? _GEN13880 : _GEN13879;
wire  _GEN13882 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13883 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13884 = io_x[24] ? _GEN13883 : _GEN13882;
wire  _GEN13885 = io_x[74] ? _GEN13884 : _GEN13881;
wire  _GEN13886 = io_x[19] ? _GEN13885 : _GEN13878;
wire  _GEN13887 = io_x[21] ? _GEN13886 : _GEN13871;
wire  _GEN13888 = io_x[23] ? _GEN13887 : _GEN13856;
wire  _GEN13889 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13890 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13891 = io_x[24] ? _GEN13890 : _GEN13889;
wire  _GEN13892 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13893 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13894 = io_x[24] ? _GEN13893 : _GEN13892;
wire  _GEN13895 = io_x[74] ? _GEN13894 : _GEN13891;
wire  _GEN13896 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13897 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13898 = io_x[24] ? _GEN13897 : _GEN13896;
wire  _GEN13899 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13900 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13901 = io_x[24] ? _GEN13900 : _GEN13899;
wire  _GEN13902 = io_x[74] ? _GEN13901 : _GEN13898;
wire  _GEN13903 = io_x[19] ? _GEN13902 : _GEN13895;
wire  _GEN13904 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13905 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13906 = io_x[24] ? _GEN13905 : _GEN13904;
wire  _GEN13907 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13908 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13909 = io_x[24] ? _GEN13908 : _GEN13907;
wire  _GEN13910 = io_x[74] ? _GEN13909 : _GEN13906;
wire  _GEN13911 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13912 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13913 = io_x[24] ? _GEN13912 : _GEN13911;
wire  _GEN13914 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13915 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13916 = io_x[24] ? _GEN13915 : _GEN13914;
wire  _GEN13917 = io_x[74] ? _GEN13916 : _GEN13913;
wire  _GEN13918 = io_x[19] ? _GEN13917 : _GEN13910;
wire  _GEN13919 = io_x[21] ? _GEN13918 : _GEN13903;
wire  _GEN13920 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13921 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13922 = io_x[24] ? _GEN13921 : _GEN13920;
wire  _GEN13923 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13924 = io_x[24] ? _GEN13923 : _GEN13606;
wire  _GEN13925 = io_x[74] ? _GEN13924 : _GEN13922;
wire  _GEN13926 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13927 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13928 = io_x[24] ? _GEN13927 : _GEN13926;
wire  _GEN13929 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13930 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13931 = io_x[24] ? _GEN13930 : _GEN13929;
wire  _GEN13932 = io_x[74] ? _GEN13931 : _GEN13928;
wire  _GEN13933 = io_x[19] ? _GEN13932 : _GEN13925;
wire  _GEN13934 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13935 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13936 = io_x[24] ? _GEN13935 : _GEN13934;
wire  _GEN13937 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13938 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13939 = io_x[24] ? _GEN13938 : _GEN13937;
wire  _GEN13940 = io_x[74] ? _GEN13939 : _GEN13936;
wire  _GEN13941 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13942 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13943 = io_x[24] ? _GEN13942 : _GEN13941;
wire  _GEN13944 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13945 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13946 = io_x[24] ? _GEN13945 : _GEN13944;
wire  _GEN13947 = io_x[74] ? _GEN13946 : _GEN13943;
wire  _GEN13948 = io_x[19] ? _GEN13947 : _GEN13940;
wire  _GEN13949 = io_x[21] ? _GEN13948 : _GEN13933;
wire  _GEN13950 = io_x[23] ? _GEN13949 : _GEN13919;
wire  _GEN13951 = io_x[25] ? _GEN13950 : _GEN13888;
wire  _GEN13952 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13953 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13954 = io_x[24] ? _GEN13953 : _GEN13952;
wire  _GEN13955 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13956 = io_x[24] ? _GEN13955 : _GEN13591;
wire  _GEN13957 = io_x[74] ? _GEN13956 : _GEN13954;
wire  _GEN13958 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13959 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13960 = io_x[24] ? _GEN13959 : _GEN13958;
wire  _GEN13961 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13962 = io_x[24] ? _GEN13961 : _GEN13606;
wire  _GEN13963 = io_x[74] ? _GEN13962 : _GEN13960;
wire  _GEN13964 = io_x[19] ? _GEN13963 : _GEN13957;
wire  _GEN13965 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13966 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13967 = io_x[24] ? _GEN13966 : _GEN13965;
wire  _GEN13968 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13969 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13970 = io_x[24] ? _GEN13969 : _GEN13968;
wire  _GEN13971 = io_x[74] ? _GEN13970 : _GEN13967;
wire  _GEN13972 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13973 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13974 = io_x[24] ? _GEN13973 : _GEN13972;
wire  _GEN13975 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13976 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13977 = io_x[24] ? _GEN13976 : _GEN13975;
wire  _GEN13978 = io_x[74] ? _GEN13977 : _GEN13974;
wire  _GEN13979 = io_x[19] ? _GEN13978 : _GEN13971;
wire  _GEN13980 = io_x[21] ? _GEN13979 : _GEN13964;
wire  _GEN13981 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13982 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13983 = io_x[24] ? _GEN13982 : _GEN13981;
wire  _GEN13984 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13985 = io_x[24] ? _GEN13606 : _GEN13984;
wire  _GEN13986 = io_x[74] ? _GEN13985 : _GEN13983;
wire  _GEN13987 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13988 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13989 = io_x[24] ? _GEN13988 : _GEN13987;
wire  _GEN13990 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13991 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13992 = io_x[24] ? _GEN13991 : _GEN13990;
wire  _GEN13993 = io_x[74] ? _GEN13992 : _GEN13989;
wire  _GEN13994 = io_x[19] ? _GEN13993 : _GEN13986;
wire  _GEN13995 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN13996 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13997 = io_x[24] ? _GEN13996 : _GEN13995;
wire  _GEN13998 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN13999 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14000 = io_x[24] ? _GEN13999 : _GEN13998;
wire  _GEN14001 = io_x[74] ? _GEN14000 : _GEN13997;
wire  _GEN14002 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14003 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14004 = io_x[24] ? _GEN14003 : _GEN14002;
wire  _GEN14005 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14006 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14007 = io_x[24] ? _GEN14006 : _GEN14005;
wire  _GEN14008 = io_x[74] ? _GEN14007 : _GEN14004;
wire  _GEN14009 = io_x[19] ? _GEN14008 : _GEN14001;
wire  _GEN14010 = io_x[21] ? _GEN14009 : _GEN13994;
wire  _GEN14011 = io_x[23] ? _GEN14010 : _GEN13980;
wire  _GEN14012 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14013 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14014 = io_x[24] ? _GEN14013 : _GEN14012;
wire  _GEN14015 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14016 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14017 = io_x[24] ? _GEN14016 : _GEN14015;
wire  _GEN14018 = io_x[74] ? _GEN14017 : _GEN14014;
wire  _GEN14019 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14020 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14021 = io_x[24] ? _GEN14020 : _GEN14019;
wire  _GEN14022 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14023 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14024 = io_x[24] ? _GEN14023 : _GEN14022;
wire  _GEN14025 = io_x[74] ? _GEN14024 : _GEN14021;
wire  _GEN14026 = io_x[19] ? _GEN14025 : _GEN14018;
wire  _GEN14027 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14028 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14029 = io_x[24] ? _GEN14028 : _GEN14027;
wire  _GEN14030 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14031 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14032 = io_x[24] ? _GEN14031 : _GEN14030;
wire  _GEN14033 = io_x[74] ? _GEN14032 : _GEN14029;
wire  _GEN14034 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14035 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14036 = io_x[24] ? _GEN14035 : _GEN14034;
wire  _GEN14037 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14038 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14039 = io_x[24] ? _GEN14038 : _GEN14037;
wire  _GEN14040 = io_x[74] ? _GEN14039 : _GEN14036;
wire  _GEN14041 = io_x[19] ? _GEN14040 : _GEN14033;
wire  _GEN14042 = io_x[21] ? _GEN14041 : _GEN14026;
wire  _GEN14043 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14044 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14045 = io_x[24] ? _GEN14044 : _GEN14043;
wire  _GEN14046 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14047 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14048 = io_x[24] ? _GEN14047 : _GEN14046;
wire  _GEN14049 = io_x[74] ? _GEN14048 : _GEN14045;
wire  _GEN14050 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14051 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14052 = io_x[24] ? _GEN14051 : _GEN14050;
wire  _GEN14053 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14054 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14055 = io_x[24] ? _GEN14054 : _GEN14053;
wire  _GEN14056 = io_x[74] ? _GEN14055 : _GEN14052;
wire  _GEN14057 = io_x[19] ? _GEN14056 : _GEN14049;
wire  _GEN14058 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14059 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14060 = io_x[24] ? _GEN14059 : _GEN14058;
wire  _GEN14061 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14062 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14063 = io_x[24] ? _GEN14062 : _GEN14061;
wire  _GEN14064 = io_x[74] ? _GEN14063 : _GEN14060;
wire  _GEN14065 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14066 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14067 = io_x[24] ? _GEN14066 : _GEN14065;
wire  _GEN14068 = io_x[20] ? _GEN13588 : _GEN13589;
wire  _GEN14069 = io_x[20] ? _GEN13589 : _GEN13588;
wire  _GEN14070 = io_x[24] ? _GEN14069 : _GEN14068;
wire  _GEN14071 = io_x[74] ? _GEN14070 : _GEN14067;
wire  _GEN14072 = io_x[19] ? _GEN14071 : _GEN14064;
wire  _GEN14073 = io_x[21] ? _GEN14072 : _GEN14057;
wire  _GEN14074 = io_x[23] ? _GEN14073 : _GEN14042;
wire  _GEN14075 = io_x[25] ? _GEN14074 : _GEN14011;
wire  _GEN14076 = io_x[16] ? _GEN14075 : _GEN13951;
wire  _GEN14077 = io_x[28] ? _GEN14076 : _GEN13829;
assign io_y[6] = _GEN14077;
wire  _GEN14078 = 1'b0;
wire  _GEN14079 = 1'b1;
wire  _GEN14080 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14081 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14082 = io_x[71] ? _GEN14081 : _GEN14080;
wire  _GEN14083 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14084 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14085 = io_x[71] ? _GEN14084 : _GEN14083;
wire  _GEN14086 = io_x[77] ? _GEN14085 : _GEN14082;
wire  _GEN14087 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14088 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14089 = io_x[71] ? _GEN14088 : _GEN14087;
wire  _GEN14090 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14091 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14092 = io_x[71] ? _GEN14091 : _GEN14090;
wire  _GEN14093 = io_x[77] ? _GEN14092 : _GEN14089;
wire  _GEN14094 = io_x[33] ? _GEN14093 : _GEN14086;
wire  _GEN14095 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14096 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14097 = io_x[71] ? _GEN14096 : _GEN14095;
wire  _GEN14098 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14099 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14100 = io_x[71] ? _GEN14099 : _GEN14098;
wire  _GEN14101 = io_x[77] ? _GEN14100 : _GEN14097;
wire  _GEN14102 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14103 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14104 = io_x[71] ? _GEN14103 : _GEN14102;
wire  _GEN14105 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14106 = io_x[73] ? _GEN14079 : _GEN14078;
wire  _GEN14107 = io_x[71] ? _GEN14106 : _GEN14105;
wire  _GEN14108 = io_x[77] ? _GEN14107 : _GEN14104;
wire  _GEN14109 = io_x[33] ? _GEN14108 : _GEN14101;
wire  _GEN14110 = io_x[72] ? _GEN14109 : _GEN14094;
assign io_y[5] = _GEN14110;
wire  _GEN14111 = 1'b0;
wire  _GEN14112 = 1'b1;
wire  _GEN14113 = io_x[72] ? _GEN14112 : _GEN14111;
wire  _GEN14114 = io_x[72] ? _GEN14112 : _GEN14111;
wire  _GEN14115 = io_x[32] ? _GEN14114 : _GEN14113;
assign io_y[4] = _GEN14115;
wire  _GEN14116 = 1'b0;
wire  _GEN14117 = 1'b1;
wire  _GEN14118 = io_x[71] ? _GEN14117 : _GEN14116;
assign io_y[3] = _GEN14118;
wire  _GEN14119 = 1'b0;
wire  _GEN14120 = 1'b1;
wire  _GEN14121 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14122 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14123 = io_x[71] ? _GEN14122 : _GEN14121;
wire  _GEN14124 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14125 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14126 = io_x[71] ? _GEN14125 : _GEN14124;
wire  _GEN14127 = io_x[21] ? _GEN14126 : _GEN14123;
wire  _GEN14128 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14129 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14130 = io_x[71] ? _GEN14129 : _GEN14128;
wire  _GEN14131 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14132 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14133 = io_x[71] ? _GEN14132 : _GEN14131;
wire  _GEN14134 = io_x[21] ? _GEN14133 : _GEN14130;
wire  _GEN14135 = io_x[19] ? _GEN14134 : _GEN14127;
wire  _GEN14136 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14137 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14138 = io_x[71] ? _GEN14137 : _GEN14136;
wire  _GEN14139 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14140 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14141 = io_x[71] ? _GEN14140 : _GEN14139;
wire  _GEN14142 = io_x[21] ? _GEN14141 : _GEN14138;
wire  _GEN14143 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14144 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14145 = io_x[71] ? _GEN14144 : _GEN14143;
wire  _GEN14146 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14147 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14148 = io_x[71] ? _GEN14147 : _GEN14146;
wire  _GEN14149 = io_x[21] ? _GEN14148 : _GEN14145;
wire  _GEN14150 = io_x[19] ? _GEN14149 : _GEN14142;
wire  _GEN14151 = io_x[79] ? _GEN14150 : _GEN14135;
wire  _GEN14152 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14153 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14154 = io_x[71] ? _GEN14153 : _GEN14152;
wire  _GEN14155 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14156 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14157 = io_x[71] ? _GEN14156 : _GEN14155;
wire  _GEN14158 = io_x[21] ? _GEN14157 : _GEN14154;
wire  _GEN14159 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14160 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14161 = io_x[71] ? _GEN14160 : _GEN14159;
wire  _GEN14162 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14163 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14164 = io_x[71] ? _GEN14163 : _GEN14162;
wire  _GEN14165 = io_x[21] ? _GEN14164 : _GEN14161;
wire  _GEN14166 = io_x[19] ? _GEN14165 : _GEN14158;
wire  _GEN14167 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14168 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14169 = io_x[71] ? _GEN14168 : _GEN14167;
wire  _GEN14170 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14171 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14172 = io_x[71] ? _GEN14171 : _GEN14170;
wire  _GEN14173 = io_x[21] ? _GEN14172 : _GEN14169;
wire  _GEN14174 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14175 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14176 = io_x[71] ? _GEN14175 : _GEN14174;
wire  _GEN14177 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14178 = io_x[70] ? _GEN14120 : _GEN14119;
wire  _GEN14179 = io_x[71] ? _GEN14178 : _GEN14177;
wire  _GEN14180 = io_x[21] ? _GEN14179 : _GEN14176;
wire  _GEN14181 = io_x[19] ? _GEN14180 : _GEN14173;
wire  _GEN14182 = io_x[79] ? _GEN14181 : _GEN14166;
wire  _GEN14183 = io_x[33] ? _GEN14182 : _GEN14151;
assign io_y[2] = _GEN14183;
wire  _GEN14184 = 1'b0;
wire  _GEN14185 = 1'b1;
wire  _GEN14186 = io_x[69] ? _GEN14185 : _GEN14184;
wire  _GEN14187 = io_x[69] ? _GEN14185 : _GEN14184;
wire  _GEN14188 = io_x[17] ? _GEN14187 : _GEN14186;
wire  _GEN14189 = io_x[69] ? _GEN14185 : _GEN14184;
wire  _GEN14190 = io_x[69] ? _GEN14185 : _GEN14184;
wire  _GEN14191 = io_x[17] ? _GEN14190 : _GEN14189;
wire  _GEN14192 = io_x[71] ? _GEN14191 : _GEN14188;
wire  _GEN14193 = io_x[69] ? _GEN14185 : _GEN14184;
wire  _GEN14194 = io_x[69] ? _GEN14185 : _GEN14184;
wire  _GEN14195 = io_x[17] ? _GEN14194 : _GEN14193;
wire  _GEN14196 = io_x[69] ? _GEN14185 : _GEN14184;
wire  _GEN14197 = io_x[69] ? _GEN14185 : _GEN14184;
wire  _GEN14198 = io_x[17] ? _GEN14197 : _GEN14196;
wire  _GEN14199 = io_x[71] ? _GEN14198 : _GEN14195;
wire  _GEN14200 = io_x[79] ? _GEN14199 : _GEN14192;
assign io_y[1] = _GEN14200;
wire  _GEN14201 = 1'b0;
wire  _GEN14202 = 1'b1;
wire  _GEN14203 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14204 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14205 = io_x[33] ? _GEN14204 : _GEN14203;
wire  _GEN14206 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14207 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14208 = io_x[33] ? _GEN14207 : _GEN14206;
wire  _GEN14209 = io_x[22] ? _GEN14208 : _GEN14205;
wire  _GEN14210 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14211 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14212 = io_x[33] ? _GEN14211 : _GEN14210;
wire  _GEN14213 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14214 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14215 = io_x[33] ? _GEN14214 : _GEN14213;
wire  _GEN14216 = io_x[22] ? _GEN14215 : _GEN14212;
wire  _GEN14217 = io_x[18] ? _GEN14216 : _GEN14209;
wire  _GEN14218 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14219 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14220 = io_x[33] ? _GEN14219 : _GEN14218;
wire  _GEN14221 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14222 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14223 = io_x[33] ? _GEN14222 : _GEN14221;
wire  _GEN14224 = io_x[22] ? _GEN14223 : _GEN14220;
wire  _GEN14225 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14226 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14227 = io_x[33] ? _GEN14226 : _GEN14225;
wire  _GEN14228 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14229 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14230 = io_x[33] ? _GEN14229 : _GEN14228;
wire  _GEN14231 = io_x[22] ? _GEN14230 : _GEN14227;
wire  _GEN14232 = io_x[18] ? _GEN14231 : _GEN14224;
wire  _GEN14233 = io_x[80] ? _GEN14232 : _GEN14217;
wire  _GEN14234 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14235 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14236 = io_x[33] ? _GEN14235 : _GEN14234;
wire  _GEN14237 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14238 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14239 = io_x[33] ? _GEN14238 : _GEN14237;
wire  _GEN14240 = io_x[22] ? _GEN14239 : _GEN14236;
wire  _GEN14241 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14242 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14243 = io_x[33] ? _GEN14242 : _GEN14241;
wire  _GEN14244 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14245 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14246 = io_x[33] ? _GEN14245 : _GEN14244;
wire  _GEN14247 = io_x[22] ? _GEN14246 : _GEN14243;
wire  _GEN14248 = io_x[18] ? _GEN14247 : _GEN14240;
wire  _GEN14249 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14250 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14251 = io_x[33] ? _GEN14250 : _GEN14249;
wire  _GEN14252 = 1'b1;
wire  _GEN14253 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14254 = io_x[33] ? _GEN14253 : _GEN14252;
wire  _GEN14255 = io_x[22] ? _GEN14254 : _GEN14251;
wire  _GEN14256 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14257 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14258 = io_x[33] ? _GEN14257 : _GEN14256;
wire  _GEN14259 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14260 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14261 = io_x[33] ? _GEN14260 : _GEN14259;
wire  _GEN14262 = io_x[22] ? _GEN14261 : _GEN14258;
wire  _GEN14263 = io_x[18] ? _GEN14262 : _GEN14255;
wire  _GEN14264 = io_x[80] ? _GEN14263 : _GEN14248;
wire  _GEN14265 = io_x[20] ? _GEN14264 : _GEN14233;
wire  _GEN14266 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14267 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14268 = io_x[33] ? _GEN14267 : _GEN14266;
wire  _GEN14269 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14270 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14271 = io_x[33] ? _GEN14270 : _GEN14269;
wire  _GEN14272 = io_x[22] ? _GEN14271 : _GEN14268;
wire  _GEN14273 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14274 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14275 = io_x[33] ? _GEN14274 : _GEN14273;
wire  _GEN14276 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14277 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14278 = io_x[33] ? _GEN14277 : _GEN14276;
wire  _GEN14279 = io_x[22] ? _GEN14278 : _GEN14275;
wire  _GEN14280 = io_x[18] ? _GEN14279 : _GEN14272;
wire  _GEN14281 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14282 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14283 = io_x[33] ? _GEN14282 : _GEN14281;
wire  _GEN14284 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14285 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14286 = io_x[33] ? _GEN14285 : _GEN14284;
wire  _GEN14287 = io_x[22] ? _GEN14286 : _GEN14283;
wire  _GEN14288 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14289 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14290 = io_x[33] ? _GEN14289 : _GEN14288;
wire  _GEN14291 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14292 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14293 = io_x[33] ? _GEN14292 : _GEN14291;
wire  _GEN14294 = io_x[22] ? _GEN14293 : _GEN14290;
wire  _GEN14295 = io_x[18] ? _GEN14294 : _GEN14287;
wire  _GEN14296 = io_x[80] ? _GEN14295 : _GEN14280;
wire  _GEN14297 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14298 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14299 = io_x[33] ? _GEN14298 : _GEN14297;
wire  _GEN14300 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14301 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14302 = io_x[33] ? _GEN14301 : _GEN14300;
wire  _GEN14303 = io_x[22] ? _GEN14302 : _GEN14299;
wire  _GEN14304 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14305 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14306 = io_x[33] ? _GEN14305 : _GEN14304;
wire  _GEN14307 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14308 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14309 = io_x[33] ? _GEN14308 : _GEN14307;
wire  _GEN14310 = io_x[22] ? _GEN14309 : _GEN14306;
wire  _GEN14311 = io_x[18] ? _GEN14310 : _GEN14303;
wire  _GEN14312 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14313 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14314 = io_x[33] ? _GEN14313 : _GEN14312;
wire  _GEN14315 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14316 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14317 = io_x[33] ? _GEN14316 : _GEN14315;
wire  _GEN14318 = io_x[22] ? _GEN14317 : _GEN14314;
wire  _GEN14319 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14320 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14321 = io_x[33] ? _GEN14320 : _GEN14319;
wire  _GEN14322 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14323 = io_x[34] ? _GEN14202 : _GEN14201;
wire  _GEN14324 = io_x[33] ? _GEN14323 : _GEN14322;
wire  _GEN14325 = io_x[22] ? _GEN14324 : _GEN14321;
wire  _GEN14326 = io_x[18] ? _GEN14325 : _GEN14318;
wire  _GEN14327 = io_x[80] ? _GEN14326 : _GEN14311;
wire  _GEN14328 = io_x[20] ? _GEN14327 : _GEN14296;
wire  _GEN14329 = io_x[16] ? _GEN14328 : _GEN14265;
assign io_y[0] = _GEN14329;
endmodule