module BBGSharePredictorImp_BSD_sim_split(
    input [31:0] pc,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    output  taken,
    output [8:0] pht_raddr,
    input [31:0] train_pc,
    input  train_taken,
    input [15:0] train_ghr_rdata,
    output  pht_wdata,
    output [8:0] pht_waddr,
    output  ghr_wdata
);

BBGSharePredictorImp_BSD_sim_pred _pred(
    .pc        (pc),
    .pht_rdata (pht_rdata),
    .ghr_rdata (ghr_rdata),
    .taken     (taken),
    .pht_raddr (pht_raddr)
);

BBGSharePredictorImp_BSD_sim_train _train(
    .train_pc        (train_pc),
    .train_taken     (train_taken),
    .train_ghr_rdata (train_ghr_rdata),
    .pht_wdata       (pht_wdata),
    .pht_waddr       (pht_waddr),
    .ghr_wdata       (ghr_wdata)
);
endmodule
module BBGSharePredictorImp_BSD_sim_pred(
    input [31:0] pc,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    output  taken,
    output [8:0] pht_raddr
);
wire [49:0] io_x;
wire [9:0] io_y;
assign io_x = { pc, pht_rdata, ghr_rdata };
assign { taken, pht_raddr } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[17] ? _GEN1 : _GEN0;
assign io_y[9] = _GEN2;
wire  _GEN3 = 1'b0;
wire  _GEN4 = 1'b1;
wire  _GEN5 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN6 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN7 = io_x[11] ? _GEN6 : _GEN5;
wire  _GEN8 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN9 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN10 = io_x[11] ? _GEN9 : _GEN8;
wire  _GEN11 = io_x[15] ? _GEN10 : _GEN7;
wire  _GEN12 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN13 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN14 = io_x[11] ? _GEN13 : _GEN12;
wire  _GEN15 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN16 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN17 = io_x[11] ? _GEN16 : _GEN15;
wire  _GEN18 = io_x[15] ? _GEN17 : _GEN14;
wire  _GEN19 = io_x[3] ? _GEN18 : _GEN11;
wire  _GEN20 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN21 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN22 = io_x[11] ? _GEN21 : _GEN20;
wire  _GEN23 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN24 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN25 = io_x[11] ? _GEN24 : _GEN23;
wire  _GEN26 = io_x[15] ? _GEN25 : _GEN22;
wire  _GEN27 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN28 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN29 = io_x[11] ? _GEN28 : _GEN27;
wire  _GEN30 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN31 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN32 = io_x[11] ? _GEN31 : _GEN30;
wire  _GEN33 = io_x[15] ? _GEN32 : _GEN29;
wire  _GEN34 = io_x[3] ? _GEN33 : _GEN26;
wire  _GEN35 = io_x[28] ? _GEN34 : _GEN19;
wire  _GEN36 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN37 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN38 = io_x[11] ? _GEN37 : _GEN36;
wire  _GEN39 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN40 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN41 = io_x[11] ? _GEN40 : _GEN39;
wire  _GEN42 = io_x[15] ? _GEN41 : _GEN38;
wire  _GEN43 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN44 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN45 = io_x[11] ? _GEN44 : _GEN43;
wire  _GEN46 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN47 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN48 = io_x[11] ? _GEN47 : _GEN46;
wire  _GEN49 = io_x[15] ? _GEN48 : _GEN45;
wire  _GEN50 = io_x[3] ? _GEN49 : _GEN42;
wire  _GEN51 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN52 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN53 = io_x[11] ? _GEN52 : _GEN51;
wire  _GEN54 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN55 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN56 = io_x[11] ? _GEN55 : _GEN54;
wire  _GEN57 = io_x[15] ? _GEN56 : _GEN53;
wire  _GEN58 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN59 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN60 = io_x[11] ? _GEN59 : _GEN58;
wire  _GEN61 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN62 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN63 = io_x[11] ? _GEN62 : _GEN61;
wire  _GEN64 = io_x[15] ? _GEN63 : _GEN60;
wire  _GEN65 = io_x[3] ? _GEN64 : _GEN57;
wire  _GEN66 = io_x[28] ? _GEN65 : _GEN50;
wire  _GEN67 = io_x[20] ? _GEN66 : _GEN35;
assign io_y[8] = _GEN67;
wire  _GEN68 = 1'b0;
wire  _GEN69 = 1'b1;
wire  _GEN70 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN71 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN72 = io_x[10] ? _GEN71 : _GEN70;
wire  _GEN73 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN74 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN75 = io_x[10] ? _GEN74 : _GEN73;
wire  _GEN76 = io_x[2] ? _GEN75 : _GEN72;
wire  _GEN77 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN78 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN79 = io_x[10] ? _GEN78 : _GEN77;
wire  _GEN80 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN81 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN82 = io_x[10] ? _GEN81 : _GEN80;
wire  _GEN83 = io_x[2] ? _GEN82 : _GEN79;
wire  _GEN84 = io_x[14] ? _GEN83 : _GEN76;
wire  _GEN85 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN86 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN87 = io_x[10] ? _GEN86 : _GEN85;
wire  _GEN88 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN89 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN90 = io_x[10] ? _GEN89 : _GEN88;
wire  _GEN91 = io_x[2] ? _GEN90 : _GEN87;
wire  _GEN92 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN93 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN94 = io_x[10] ? _GEN93 : _GEN92;
wire  _GEN95 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN96 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN97 = io_x[10] ? _GEN96 : _GEN95;
wire  _GEN98 = io_x[2] ? _GEN97 : _GEN94;
wire  _GEN99 = io_x[14] ? _GEN98 : _GEN91;
wire  _GEN100 = io_x[27] ? _GEN99 : _GEN84;
wire  _GEN101 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN102 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN103 = io_x[10] ? _GEN102 : _GEN101;
wire  _GEN104 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN105 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN106 = io_x[10] ? _GEN105 : _GEN104;
wire  _GEN107 = io_x[2] ? _GEN106 : _GEN103;
wire  _GEN108 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN109 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN110 = io_x[10] ? _GEN109 : _GEN108;
wire  _GEN111 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN112 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN113 = io_x[10] ? _GEN112 : _GEN111;
wire  _GEN114 = io_x[2] ? _GEN113 : _GEN110;
wire  _GEN115 = io_x[14] ? _GEN114 : _GEN107;
wire  _GEN116 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN117 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN118 = io_x[10] ? _GEN117 : _GEN116;
wire  _GEN119 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN120 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN121 = io_x[10] ? _GEN120 : _GEN119;
wire  _GEN122 = io_x[2] ? _GEN121 : _GEN118;
wire  _GEN123 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN124 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN125 = io_x[10] ? _GEN124 : _GEN123;
wire  _GEN126 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN127 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN128 = io_x[10] ? _GEN127 : _GEN126;
wire  _GEN129 = io_x[2] ? _GEN128 : _GEN125;
wire  _GEN130 = io_x[14] ? _GEN129 : _GEN122;
wire  _GEN131 = io_x[27] ? _GEN130 : _GEN115;
wire  _GEN132 = io_x[25] ? _GEN131 : _GEN100;
assign io_y[7] = _GEN132;
wire  _GEN133 = 1'b0;
wire  _GEN134 = 1'b1;
wire  _GEN135 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN136 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN137 = io_x[9] ? _GEN136 : _GEN135;
wire  _GEN138 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN139 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN140 = io_x[9] ? _GEN139 : _GEN138;
wire  _GEN141 = io_x[1] ? _GEN140 : _GEN137;
wire  _GEN142 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN143 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN144 = io_x[9] ? _GEN143 : _GEN142;
wire  _GEN145 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN146 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN147 = io_x[9] ? _GEN146 : _GEN145;
wire  _GEN148 = io_x[1] ? _GEN147 : _GEN144;
wire  _GEN149 = io_x[13] ? _GEN148 : _GEN141;
wire  _GEN150 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN151 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN152 = io_x[9] ? _GEN151 : _GEN150;
wire  _GEN153 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN154 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN155 = io_x[9] ? _GEN154 : _GEN153;
wire  _GEN156 = io_x[1] ? _GEN155 : _GEN152;
wire  _GEN157 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN158 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN159 = io_x[9] ? _GEN158 : _GEN157;
wire  _GEN160 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN161 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN162 = io_x[9] ? _GEN161 : _GEN160;
wire  _GEN163 = io_x[1] ? _GEN162 : _GEN159;
wire  _GEN164 = io_x[13] ? _GEN163 : _GEN156;
wire  _GEN165 = io_x[26] ? _GEN164 : _GEN149;
wire  _GEN166 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN167 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN168 = io_x[9] ? _GEN167 : _GEN166;
wire  _GEN169 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN170 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN171 = io_x[9] ? _GEN170 : _GEN169;
wire  _GEN172 = io_x[1] ? _GEN171 : _GEN168;
wire  _GEN173 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN174 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN175 = io_x[9] ? _GEN174 : _GEN173;
wire  _GEN176 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN177 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN178 = io_x[9] ? _GEN177 : _GEN176;
wire  _GEN179 = io_x[1] ? _GEN178 : _GEN175;
wire  _GEN180 = io_x[13] ? _GEN179 : _GEN172;
wire  _GEN181 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN182 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN183 = io_x[9] ? _GEN182 : _GEN181;
wire  _GEN184 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN185 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN186 = io_x[9] ? _GEN185 : _GEN184;
wire  _GEN187 = io_x[1] ? _GEN186 : _GEN183;
wire  _GEN188 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN189 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN190 = io_x[9] ? _GEN189 : _GEN188;
wire  _GEN191 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN192 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN193 = io_x[9] ? _GEN192 : _GEN191;
wire  _GEN194 = io_x[1] ? _GEN193 : _GEN190;
wire  _GEN195 = io_x[13] ? _GEN194 : _GEN187;
wire  _GEN196 = io_x[26] ? _GEN195 : _GEN180;
wire  _GEN197 = io_x[11] ? _GEN196 : _GEN165;
assign io_y[6] = _GEN197;
wire  _GEN198 = 1'b0;
wire  _GEN199 = 1'b1;
wire  _GEN200 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN201 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN202 = io_x[12] ? _GEN201 : _GEN200;
wire  _GEN203 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN204 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN205 = io_x[12] ? _GEN204 : _GEN203;
wire  _GEN206 = io_x[4] ? _GEN205 : _GEN202;
wire  _GEN207 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN208 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN209 = io_x[12] ? _GEN208 : _GEN207;
wire  _GEN210 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN211 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN212 = io_x[12] ? _GEN211 : _GEN210;
wire  _GEN213 = io_x[4] ? _GEN212 : _GEN209;
wire  _GEN214 = io_x[0] ? _GEN213 : _GEN206;
wire  _GEN215 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN216 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN217 = io_x[12] ? _GEN216 : _GEN215;
wire  _GEN218 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN219 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN220 = io_x[12] ? _GEN219 : _GEN218;
wire  _GEN221 = io_x[4] ? _GEN220 : _GEN217;
wire  _GEN222 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN223 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN224 = io_x[12] ? _GEN223 : _GEN222;
wire  _GEN225 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN226 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN227 = io_x[12] ? _GEN226 : _GEN225;
wire  _GEN228 = io_x[4] ? _GEN227 : _GEN224;
wire  _GEN229 = io_x[0] ? _GEN228 : _GEN221;
wire  _GEN230 = io_x[25] ? _GEN229 : _GEN214;
wire  _GEN231 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN232 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN233 = io_x[12] ? _GEN232 : _GEN231;
wire  _GEN234 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN235 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN236 = io_x[12] ? _GEN235 : _GEN234;
wire  _GEN237 = io_x[4] ? _GEN236 : _GEN233;
wire  _GEN238 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN239 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN240 = io_x[12] ? _GEN239 : _GEN238;
wire  _GEN241 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN242 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN243 = io_x[12] ? _GEN242 : _GEN241;
wire  _GEN244 = io_x[4] ? _GEN243 : _GEN240;
wire  _GEN245 = io_x[0] ? _GEN244 : _GEN237;
wire  _GEN246 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN247 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN248 = io_x[12] ? _GEN247 : _GEN246;
wire  _GEN249 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN250 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN251 = io_x[12] ? _GEN250 : _GEN249;
wire  _GEN252 = io_x[4] ? _GEN251 : _GEN248;
wire  _GEN253 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN254 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN255 = io_x[12] ? _GEN254 : _GEN253;
wire  _GEN256 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN257 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN258 = io_x[12] ? _GEN257 : _GEN256;
wire  _GEN259 = io_x[4] ? _GEN258 : _GEN255;
wire  _GEN260 = io_x[0] ? _GEN259 : _GEN252;
wire  _GEN261 = io_x[25] ? _GEN260 : _GEN245;
wire  _GEN262 = io_x[23] ? _GEN261 : _GEN230;
assign io_y[5] = _GEN262;
wire  _GEN263 = 1'b0;
wire  _GEN264 = 1'b1;
wire  _GEN265 = io_x[24] ? _GEN264 : _GEN263;
wire  _GEN266 = io_x[24] ? _GEN264 : _GEN263;
wire  _GEN267 = io_x[20] ? _GEN266 : _GEN265;
assign io_y[4] = _GEN267;
wire  _GEN268 = 1'b0;
wire  _GEN269 = 1'b1;
wire  _GEN270 = io_x[23] ? _GEN269 : _GEN268;
wire  _GEN271 = io_x[23] ? _GEN269 : _GEN268;
wire  _GEN272 = io_x[29] ? _GEN271 : _GEN270;
assign io_y[3] = _GEN272;
wire  _GEN273 = 1'b0;
wire  _GEN274 = 1'b1;
wire  _GEN275 = io_x[22] ? _GEN274 : _GEN273;
assign io_y[2] = _GEN275;
wire  _GEN276 = 1'b0;
wire  _GEN277 = 1'b1;
wire  _GEN278 = io_x[21] ? _GEN277 : _GEN276;
wire  _GEN279 = io_x[21] ? _GEN277 : _GEN276;
wire  _GEN280 = io_x[24] ? _GEN279 : _GEN278;
wire  _GEN281 = io_x[21] ? _GEN277 : _GEN276;
wire  _GEN282 = io_x[21] ? _GEN277 : _GEN276;
wire  _GEN283 = io_x[24] ? _GEN282 : _GEN281;
wire  _GEN284 = io_x[25] ? _GEN283 : _GEN280;
assign io_y[1] = _GEN284;
wire  _GEN285 = 1'b0;
wire  _GEN286 = 1'b1;
wire  _GEN287 = io_x[20] ? _GEN286 : _GEN285;
wire  _GEN288 = io_x[20] ? _GEN286 : _GEN285;
wire  _GEN289 = io_x[24] ? _GEN288 : _GEN287;
wire  _GEN290 = io_x[20] ? _GEN286 : _GEN285;
wire  _GEN291 = io_x[20] ? _GEN286 : _GEN285;
wire  _GEN292 = io_x[24] ? _GEN291 : _GEN290;
wire  _GEN293 = io_x[29] ? _GEN292 : _GEN289;
assign io_y[0] = _GEN293;
endmodule
module BBGSharePredictorImp_BSD_sim_train(
    input [31:0] train_pc,
    input  train_taken,
    input [15:0] train_ghr_rdata,
    output  pht_wdata,
    output [8:0] pht_waddr,
    output  ghr_wdata
);
wire [48:0] io_x;
wire [10:0] io_y;
assign io_x = { train_pc, train_taken, train_ghr_rdata };
assign { pht_wdata, pht_waddr, ghr_wdata } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[16] ? _GEN1 : _GEN0;
assign io_y[10] = _GEN2;
wire  _GEN3 = 1'b0;
wire  _GEN4 = 1'b1;
wire  _GEN5 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN6 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN7 = io_x[11] ? _GEN6 : _GEN5;
wire  _GEN8 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN9 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN10 = io_x[11] ? _GEN9 : _GEN8;
wire  _GEN11 = io_x[15] ? _GEN10 : _GEN7;
wire  _GEN12 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN13 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN14 = io_x[11] ? _GEN13 : _GEN12;
wire  _GEN15 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN16 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN17 = io_x[11] ? _GEN16 : _GEN15;
wire  _GEN18 = io_x[15] ? _GEN17 : _GEN14;
wire  _GEN19 = io_x[3] ? _GEN18 : _GEN11;
wire  _GEN20 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN21 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN22 = io_x[11] ? _GEN21 : _GEN20;
wire  _GEN23 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN24 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN25 = io_x[11] ? _GEN24 : _GEN23;
wire  _GEN26 = io_x[15] ? _GEN25 : _GEN22;
wire  _GEN27 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN28 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN29 = io_x[11] ? _GEN28 : _GEN27;
wire  _GEN30 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN31 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN32 = io_x[11] ? _GEN31 : _GEN30;
wire  _GEN33 = io_x[15] ? _GEN32 : _GEN29;
wire  _GEN34 = io_x[3] ? _GEN33 : _GEN26;
wire  _GEN35 = io_x[27] ? _GEN34 : _GEN19;
wire  _GEN36 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN37 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN38 = io_x[11] ? _GEN37 : _GEN36;
wire  _GEN39 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN40 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN41 = io_x[11] ? _GEN40 : _GEN39;
wire  _GEN42 = io_x[15] ? _GEN41 : _GEN38;
wire  _GEN43 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN44 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN45 = io_x[11] ? _GEN44 : _GEN43;
wire  _GEN46 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN47 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN48 = io_x[11] ? _GEN47 : _GEN46;
wire  _GEN49 = io_x[15] ? _GEN48 : _GEN45;
wire  _GEN50 = io_x[3] ? _GEN49 : _GEN42;
wire  _GEN51 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN52 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN53 = io_x[11] ? _GEN52 : _GEN51;
wire  _GEN54 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN55 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN56 = io_x[11] ? _GEN55 : _GEN54;
wire  _GEN57 = io_x[15] ? _GEN56 : _GEN53;
wire  _GEN58 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN59 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN60 = io_x[11] ? _GEN59 : _GEN58;
wire  _GEN61 = io_x[7] ? _GEN3 : _GEN4;
wire  _GEN62 = io_x[7] ? _GEN4 : _GEN3;
wire  _GEN63 = io_x[11] ? _GEN62 : _GEN61;
wire  _GEN64 = io_x[15] ? _GEN63 : _GEN60;
wire  _GEN65 = io_x[3] ? _GEN64 : _GEN57;
wire  _GEN66 = io_x[27] ? _GEN65 : _GEN50;
wire  _GEN67 = io_x[19] ? _GEN66 : _GEN35;
assign io_y[9] = _GEN67;
wire  _GEN68 = 1'b0;
wire  _GEN69 = 1'b1;
wire  _GEN70 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN71 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN72 = io_x[10] ? _GEN71 : _GEN70;
wire  _GEN73 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN74 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN75 = io_x[10] ? _GEN74 : _GEN73;
wire  _GEN76 = io_x[2] ? _GEN75 : _GEN72;
wire  _GEN77 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN78 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN79 = io_x[10] ? _GEN78 : _GEN77;
wire  _GEN80 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN81 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN82 = io_x[10] ? _GEN81 : _GEN80;
wire  _GEN83 = io_x[2] ? _GEN82 : _GEN79;
wire  _GEN84 = io_x[14] ? _GEN83 : _GEN76;
wire  _GEN85 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN86 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN87 = io_x[10] ? _GEN86 : _GEN85;
wire  _GEN88 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN89 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN90 = io_x[10] ? _GEN89 : _GEN88;
wire  _GEN91 = io_x[2] ? _GEN90 : _GEN87;
wire  _GEN92 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN93 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN94 = io_x[10] ? _GEN93 : _GEN92;
wire  _GEN95 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN96 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN97 = io_x[10] ? _GEN96 : _GEN95;
wire  _GEN98 = io_x[2] ? _GEN97 : _GEN94;
wire  _GEN99 = io_x[14] ? _GEN98 : _GEN91;
wire  _GEN100 = io_x[26] ? _GEN99 : _GEN84;
wire  _GEN101 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN102 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN103 = io_x[10] ? _GEN102 : _GEN101;
wire  _GEN104 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN105 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN106 = io_x[10] ? _GEN105 : _GEN104;
wire  _GEN107 = io_x[2] ? _GEN106 : _GEN103;
wire  _GEN108 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN109 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN110 = io_x[10] ? _GEN109 : _GEN108;
wire  _GEN111 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN112 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN113 = io_x[10] ? _GEN112 : _GEN111;
wire  _GEN114 = io_x[2] ? _GEN113 : _GEN110;
wire  _GEN115 = io_x[14] ? _GEN114 : _GEN107;
wire  _GEN116 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN117 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN118 = io_x[10] ? _GEN117 : _GEN116;
wire  _GEN119 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN120 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN121 = io_x[10] ? _GEN120 : _GEN119;
wire  _GEN122 = io_x[2] ? _GEN121 : _GEN118;
wire  _GEN123 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN124 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN125 = io_x[10] ? _GEN124 : _GEN123;
wire  _GEN126 = io_x[6] ? _GEN68 : _GEN69;
wire  _GEN127 = io_x[6] ? _GEN69 : _GEN68;
wire  _GEN128 = io_x[10] ? _GEN127 : _GEN126;
wire  _GEN129 = io_x[2] ? _GEN128 : _GEN125;
wire  _GEN130 = io_x[14] ? _GEN129 : _GEN122;
wire  _GEN131 = io_x[26] ? _GEN130 : _GEN115;
wire  _GEN132 = io_x[24] ? _GEN131 : _GEN100;
assign io_y[8] = _GEN132;
wire  _GEN133 = 1'b0;
wire  _GEN134 = 1'b1;
wire  _GEN135 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN136 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN137 = io_x[9] ? _GEN136 : _GEN135;
wire  _GEN138 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN139 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN140 = io_x[9] ? _GEN139 : _GEN138;
wire  _GEN141 = io_x[1] ? _GEN140 : _GEN137;
wire  _GEN142 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN143 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN144 = io_x[9] ? _GEN143 : _GEN142;
wire  _GEN145 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN146 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN147 = io_x[9] ? _GEN146 : _GEN145;
wire  _GEN148 = io_x[1] ? _GEN147 : _GEN144;
wire  _GEN149 = io_x[13] ? _GEN148 : _GEN141;
wire  _GEN150 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN151 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN152 = io_x[9] ? _GEN151 : _GEN150;
wire  _GEN153 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN154 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN155 = io_x[9] ? _GEN154 : _GEN153;
wire  _GEN156 = io_x[1] ? _GEN155 : _GEN152;
wire  _GEN157 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN158 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN159 = io_x[9] ? _GEN158 : _GEN157;
wire  _GEN160 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN161 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN162 = io_x[9] ? _GEN161 : _GEN160;
wire  _GEN163 = io_x[1] ? _GEN162 : _GEN159;
wire  _GEN164 = io_x[13] ? _GEN163 : _GEN156;
wire  _GEN165 = io_x[25] ? _GEN164 : _GEN149;
wire  _GEN166 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN167 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN168 = io_x[9] ? _GEN167 : _GEN166;
wire  _GEN169 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN170 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN171 = io_x[9] ? _GEN170 : _GEN169;
wire  _GEN172 = io_x[1] ? _GEN171 : _GEN168;
wire  _GEN173 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN174 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN175 = io_x[9] ? _GEN174 : _GEN173;
wire  _GEN176 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN177 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN178 = io_x[9] ? _GEN177 : _GEN176;
wire  _GEN179 = io_x[1] ? _GEN178 : _GEN175;
wire  _GEN180 = io_x[13] ? _GEN179 : _GEN172;
wire  _GEN181 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN182 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN183 = io_x[9] ? _GEN182 : _GEN181;
wire  _GEN184 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN185 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN186 = io_x[9] ? _GEN185 : _GEN184;
wire  _GEN187 = io_x[1] ? _GEN186 : _GEN183;
wire  _GEN188 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN189 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN190 = io_x[9] ? _GEN189 : _GEN188;
wire  _GEN191 = io_x[5] ? _GEN133 : _GEN134;
wire  _GEN192 = io_x[5] ? _GEN134 : _GEN133;
wire  _GEN193 = io_x[9] ? _GEN192 : _GEN191;
wire  _GEN194 = io_x[1] ? _GEN193 : _GEN190;
wire  _GEN195 = io_x[13] ? _GEN194 : _GEN187;
wire  _GEN196 = io_x[25] ? _GEN195 : _GEN180;
wire  _GEN197 = io_x[11] ? _GEN196 : _GEN165;
assign io_y[7] = _GEN197;
wire  _GEN198 = 1'b0;
wire  _GEN199 = 1'b1;
wire  _GEN200 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN201 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN202 = io_x[12] ? _GEN201 : _GEN200;
wire  _GEN203 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN204 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN205 = io_x[12] ? _GEN204 : _GEN203;
wire  _GEN206 = io_x[4] ? _GEN205 : _GEN202;
wire  _GEN207 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN208 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN209 = io_x[12] ? _GEN208 : _GEN207;
wire  _GEN210 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN211 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN212 = io_x[12] ? _GEN211 : _GEN210;
wire  _GEN213 = io_x[4] ? _GEN212 : _GEN209;
wire  _GEN214 = io_x[0] ? _GEN213 : _GEN206;
wire  _GEN215 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN216 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN217 = io_x[12] ? _GEN216 : _GEN215;
wire  _GEN218 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN219 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN220 = io_x[12] ? _GEN219 : _GEN218;
wire  _GEN221 = io_x[4] ? _GEN220 : _GEN217;
wire  _GEN222 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN223 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN224 = io_x[12] ? _GEN223 : _GEN222;
wire  _GEN225 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN226 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN227 = io_x[12] ? _GEN226 : _GEN225;
wire  _GEN228 = io_x[4] ? _GEN227 : _GEN224;
wire  _GEN229 = io_x[0] ? _GEN228 : _GEN221;
wire  _GEN230 = io_x[24] ? _GEN229 : _GEN214;
wire  _GEN231 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN232 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN233 = io_x[12] ? _GEN232 : _GEN231;
wire  _GEN234 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN235 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN236 = io_x[12] ? _GEN235 : _GEN234;
wire  _GEN237 = io_x[4] ? _GEN236 : _GEN233;
wire  _GEN238 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN239 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN240 = io_x[12] ? _GEN239 : _GEN238;
wire  _GEN241 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN242 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN243 = io_x[12] ? _GEN242 : _GEN241;
wire  _GEN244 = io_x[4] ? _GEN243 : _GEN240;
wire  _GEN245 = io_x[0] ? _GEN244 : _GEN237;
wire  _GEN246 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN247 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN248 = io_x[12] ? _GEN247 : _GEN246;
wire  _GEN249 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN250 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN251 = io_x[12] ? _GEN250 : _GEN249;
wire  _GEN252 = io_x[4] ? _GEN251 : _GEN248;
wire  _GEN253 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN254 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN255 = io_x[12] ? _GEN254 : _GEN253;
wire  _GEN256 = io_x[8] ? _GEN198 : _GEN199;
wire  _GEN257 = io_x[8] ? _GEN199 : _GEN198;
wire  _GEN258 = io_x[12] ? _GEN257 : _GEN256;
wire  _GEN259 = io_x[4] ? _GEN258 : _GEN255;
wire  _GEN260 = io_x[0] ? _GEN259 : _GEN252;
wire  _GEN261 = io_x[24] ? _GEN260 : _GEN245;
wire  _GEN262 = io_x[22] ? _GEN261 : _GEN230;
assign io_y[6] = _GEN262;
wire  _GEN263 = 1'b0;
wire  _GEN264 = 1'b1;
wire  _GEN265 = io_x[23] ? _GEN264 : _GEN263;
wire  _GEN266 = io_x[23] ? _GEN264 : _GEN263;
wire  _GEN267 = io_x[19] ? _GEN266 : _GEN265;
assign io_y[5] = _GEN267;
wire  _GEN268 = 1'b0;
wire  _GEN269 = 1'b1;
wire  _GEN270 = io_x[22] ? _GEN269 : _GEN268;
wire  _GEN271 = io_x[22] ? _GEN269 : _GEN268;
wire  _GEN272 = io_x[28] ? _GEN271 : _GEN270;
assign io_y[4] = _GEN272;
wire  _GEN273 = 1'b0;
wire  _GEN274 = 1'b1;
wire  _GEN275 = io_x[21] ? _GEN274 : _GEN273;
assign io_y[3] = _GEN275;
wire  _GEN276 = 1'b0;
wire  _GEN277 = 1'b1;
wire  _GEN278 = io_x[20] ? _GEN277 : _GEN276;
wire  _GEN279 = io_x[20] ? _GEN277 : _GEN276;
wire  _GEN280 = io_x[23] ? _GEN279 : _GEN278;
wire  _GEN281 = io_x[20] ? _GEN277 : _GEN276;
wire  _GEN282 = io_x[20] ? _GEN277 : _GEN276;
wire  _GEN283 = io_x[23] ? _GEN282 : _GEN281;
wire  _GEN284 = io_x[24] ? _GEN283 : _GEN280;
assign io_y[2] = _GEN284;
wire  _GEN285 = 1'b0;
wire  _GEN286 = 1'b1;
wire  _GEN287 = io_x[19] ? _GEN286 : _GEN285;
wire  _GEN288 = io_x[19] ? _GEN286 : _GEN285;
wire  _GEN289 = io_x[23] ? _GEN288 : _GEN287;
wire  _GEN290 = io_x[19] ? _GEN286 : _GEN285;
wire  _GEN291 = io_x[19] ? _GEN286 : _GEN285;
wire  _GEN292 = io_x[23] ? _GEN291 : _GEN290;
wire  _GEN293 = io_x[28] ? _GEN292 : _GEN289;
assign io_y[1] = _GEN293;
wire  _GEN294 = 1'b0;
wire  _GEN295 = 1'b1;
wire  _GEN296 = io_x[16] ? _GEN295 : _GEN294;
assign io_y[0] = _GEN296;
endmodule
