module BBGSharePredictorImp_BSD_b_NutShell(
    input [31:0] pc,
    input [31:0] train_pc,
    input  train_taken,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    input [15:0] train_ghr_rdata,
    output  taken,
    output  pht_wdata,
    output [8:0] pht_raddr,
    output [8:0] pht_waddr,
    output  ghr_wdata
);
wire [98:0] io_x;
wire [20:0] io_y;
assign io_x = { pc, train_pc, train_taken, pht_rdata, ghr_rdata, train_ghr_rdata };
assign { taken, pht_wdata, pht_raddr, pht_waddr, ghr_wdata } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN3 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN4 = io_x[32] ? _GEN3 : _GEN2;
wire  _GEN5 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN6 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN7 = io_x[32] ? _GEN6 : _GEN5;
wire  _GEN8 = io_x[45] ? _GEN7 : _GEN4;
wire  _GEN9 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN10 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN11 = io_x[32] ? _GEN10 : _GEN9;
wire  _GEN12 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN13 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN14 = io_x[32] ? _GEN13 : _GEN12;
wire  _GEN15 = io_x[45] ? _GEN14 : _GEN11;
wire  _GEN16 = io_x[42] ? _GEN15 : _GEN8;
assign io_y[20] = _GEN16;
wire  _GEN17 = 1'b0;
wire  _GEN18 = 1'b1;
wire  _GEN19 = io_x[34] ? _GEN18 : _GEN17;
wire  _GEN20 = io_x[34] ? _GEN18 : _GEN17;
wire  _GEN21 = io_x[77] ? _GEN20 : _GEN19;
assign io_y[19] = _GEN21;
wire  _GEN22 = 1'b0;
wire  _GEN23 = 1'b1;
wire  _GEN24 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN25 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN26 = io_x[19] ? _GEN25 : _GEN24;
wire  _GEN27 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN28 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN29 = io_x[19] ? _GEN28 : _GEN27;
wire  _GEN30 = io_x[23] ? _GEN29 : _GEN26;
wire  _GEN31 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN32 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN33 = io_x[19] ? _GEN32 : _GEN31;
wire  _GEN34 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN35 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN36 = io_x[19] ? _GEN35 : _GEN34;
wire  _GEN37 = io_x[23] ? _GEN36 : _GEN33;
wire  _GEN38 = io_x[27] ? _GEN37 : _GEN30;
wire  _GEN39 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN40 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN41 = io_x[19] ? _GEN40 : _GEN39;
wire  _GEN42 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN43 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN44 = io_x[19] ? _GEN43 : _GEN42;
wire  _GEN45 = io_x[23] ? _GEN44 : _GEN41;
wire  _GEN46 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN47 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN48 = io_x[19] ? _GEN47 : _GEN46;
wire  _GEN49 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN50 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN51 = io_x[19] ? _GEN50 : _GEN49;
wire  _GEN52 = io_x[23] ? _GEN51 : _GEN48;
wire  _GEN53 = io_x[27] ? _GEN52 : _GEN45;
wire  _GEN54 = io_x[48] ? _GEN53 : _GEN38;
wire  _GEN55 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN56 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN57 = io_x[19] ? _GEN56 : _GEN55;
wire  _GEN58 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN59 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN60 = io_x[19] ? _GEN59 : _GEN58;
wire  _GEN61 = io_x[23] ? _GEN60 : _GEN57;
wire  _GEN62 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN63 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN64 = io_x[19] ? _GEN63 : _GEN62;
wire  _GEN65 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN66 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN67 = io_x[19] ? _GEN66 : _GEN65;
wire  _GEN68 = io_x[23] ? _GEN67 : _GEN64;
wire  _GEN69 = io_x[27] ? _GEN68 : _GEN61;
wire  _GEN70 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN71 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN72 = io_x[19] ? _GEN71 : _GEN70;
wire  _GEN73 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN74 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN75 = io_x[19] ? _GEN74 : _GEN73;
wire  _GEN76 = io_x[23] ? _GEN75 : _GEN72;
wire  _GEN77 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN78 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN79 = io_x[19] ? _GEN78 : _GEN77;
wire  _GEN80 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN81 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN82 = io_x[19] ? _GEN81 : _GEN80;
wire  _GEN83 = io_x[23] ? _GEN82 : _GEN79;
wire  _GEN84 = io_x[27] ? _GEN83 : _GEN76;
wire  _GEN85 = io_x[48] ? _GEN84 : _GEN69;
wire  _GEN86 = io_x[31] ? _GEN85 : _GEN54;
wire  _GEN87 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN88 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN89 = io_x[19] ? _GEN88 : _GEN87;
wire  _GEN90 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN91 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN92 = io_x[19] ? _GEN91 : _GEN90;
wire  _GEN93 = io_x[23] ? _GEN92 : _GEN89;
wire  _GEN94 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN95 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN96 = io_x[19] ? _GEN95 : _GEN94;
wire  _GEN97 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN98 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN99 = io_x[19] ? _GEN98 : _GEN97;
wire  _GEN100 = io_x[23] ? _GEN99 : _GEN96;
wire  _GEN101 = io_x[27] ? _GEN100 : _GEN93;
wire  _GEN102 = 1'b0;
wire  _GEN103 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN104 = io_x[19] ? _GEN103 : _GEN102;
wire  _GEN105 = 1'b1;
wire  _GEN106 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN107 = io_x[19] ? _GEN106 : _GEN105;
wire  _GEN108 = io_x[23] ? _GEN107 : _GEN104;
wire  _GEN109 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN110 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN111 = io_x[19] ? _GEN110 : _GEN109;
wire  _GEN112 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN113 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN114 = io_x[19] ? _GEN113 : _GEN112;
wire  _GEN115 = io_x[23] ? _GEN114 : _GEN111;
wire  _GEN116 = io_x[27] ? _GEN115 : _GEN108;
wire  _GEN117 = io_x[48] ? _GEN116 : _GEN101;
wire  _GEN118 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN119 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN120 = io_x[19] ? _GEN119 : _GEN118;
wire  _GEN121 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN122 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN123 = io_x[19] ? _GEN122 : _GEN121;
wire  _GEN124 = io_x[23] ? _GEN123 : _GEN120;
wire  _GEN125 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN126 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN127 = io_x[19] ? _GEN126 : _GEN125;
wire  _GEN128 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN129 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN130 = io_x[19] ? _GEN129 : _GEN128;
wire  _GEN131 = io_x[23] ? _GEN130 : _GEN127;
wire  _GEN132 = io_x[27] ? _GEN131 : _GEN124;
wire  _GEN133 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN134 = io_x[19] ? _GEN133 : _GEN105;
wire  _GEN135 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN136 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN137 = io_x[19] ? _GEN136 : _GEN135;
wire  _GEN138 = io_x[23] ? _GEN137 : _GEN134;
wire  _GEN139 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN140 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN141 = io_x[19] ? _GEN140 : _GEN139;
wire  _GEN142 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN143 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN144 = io_x[19] ? _GEN143 : _GEN142;
wire  _GEN145 = io_x[23] ? _GEN144 : _GEN141;
wire  _GEN146 = io_x[27] ? _GEN145 : _GEN138;
wire  _GEN147 = io_x[48] ? _GEN146 : _GEN132;
wire  _GEN148 = io_x[31] ? _GEN147 : _GEN117;
wire  _GEN149 = io_x[3] ? _GEN148 : _GEN86;
wire  _GEN150 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN151 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN152 = io_x[19] ? _GEN151 : _GEN150;
wire  _GEN153 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN154 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN155 = io_x[19] ? _GEN154 : _GEN153;
wire  _GEN156 = io_x[23] ? _GEN155 : _GEN152;
wire  _GEN157 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN158 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN159 = io_x[19] ? _GEN158 : _GEN157;
wire  _GEN160 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN161 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN162 = io_x[19] ? _GEN161 : _GEN160;
wire  _GEN163 = io_x[23] ? _GEN162 : _GEN159;
wire  _GEN164 = io_x[27] ? _GEN163 : _GEN156;
wire  _GEN165 = io_x[19] ? _GEN105 : _GEN102;
wire  _GEN166 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN167 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN168 = io_x[19] ? _GEN167 : _GEN166;
wire  _GEN169 = io_x[23] ? _GEN168 : _GEN165;
wire  _GEN170 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN171 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN172 = io_x[19] ? _GEN171 : _GEN170;
wire  _GEN173 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN174 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN175 = io_x[19] ? _GEN174 : _GEN173;
wire  _GEN176 = io_x[23] ? _GEN175 : _GEN172;
wire  _GEN177 = io_x[27] ? _GEN176 : _GEN169;
wire  _GEN178 = io_x[48] ? _GEN177 : _GEN164;
wire  _GEN179 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN180 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN181 = io_x[19] ? _GEN180 : _GEN179;
wire  _GEN182 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN183 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN184 = io_x[19] ? _GEN183 : _GEN182;
wire  _GEN185 = io_x[23] ? _GEN184 : _GEN181;
wire  _GEN186 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN187 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN188 = io_x[19] ? _GEN187 : _GEN186;
wire  _GEN189 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN190 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN191 = io_x[19] ? _GEN190 : _GEN189;
wire  _GEN192 = io_x[23] ? _GEN191 : _GEN188;
wire  _GEN193 = io_x[27] ? _GEN192 : _GEN185;
wire  _GEN194 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN195 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN196 = io_x[19] ? _GEN195 : _GEN194;
wire  _GEN197 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN198 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN199 = io_x[19] ? _GEN198 : _GEN197;
wire  _GEN200 = io_x[23] ? _GEN199 : _GEN196;
wire  _GEN201 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN202 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN203 = io_x[19] ? _GEN202 : _GEN201;
wire  _GEN204 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN205 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN206 = io_x[19] ? _GEN205 : _GEN204;
wire  _GEN207 = io_x[23] ? _GEN206 : _GEN203;
wire  _GEN208 = io_x[27] ? _GEN207 : _GEN200;
wire  _GEN209 = io_x[48] ? _GEN208 : _GEN193;
wire  _GEN210 = io_x[31] ? _GEN209 : _GEN178;
wire  _GEN211 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN212 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN213 = io_x[19] ? _GEN212 : _GEN211;
wire  _GEN214 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN215 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN216 = io_x[19] ? _GEN215 : _GEN214;
wire  _GEN217 = io_x[23] ? _GEN216 : _GEN213;
wire  _GEN218 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN219 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN220 = io_x[19] ? _GEN219 : _GEN218;
wire  _GEN221 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN222 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN223 = io_x[19] ? _GEN222 : _GEN221;
wire  _GEN224 = io_x[23] ? _GEN223 : _GEN220;
wire  _GEN225 = io_x[27] ? _GEN224 : _GEN217;
wire  _GEN226 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN227 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN228 = io_x[19] ? _GEN227 : _GEN226;
wire  _GEN229 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN230 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN231 = io_x[19] ? _GEN230 : _GEN229;
wire  _GEN232 = io_x[23] ? _GEN231 : _GEN228;
wire  _GEN233 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN234 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN235 = io_x[19] ? _GEN234 : _GEN233;
wire  _GEN236 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN237 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN238 = io_x[19] ? _GEN237 : _GEN236;
wire  _GEN239 = io_x[23] ? _GEN238 : _GEN235;
wire  _GEN240 = io_x[27] ? _GEN239 : _GEN232;
wire  _GEN241 = io_x[48] ? _GEN240 : _GEN225;
wire  _GEN242 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN243 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN244 = io_x[19] ? _GEN243 : _GEN242;
wire  _GEN245 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN246 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN247 = io_x[19] ? _GEN246 : _GEN245;
wire  _GEN248 = io_x[23] ? _GEN247 : _GEN244;
wire  _GEN249 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN250 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN251 = io_x[19] ? _GEN250 : _GEN249;
wire  _GEN252 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN253 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN254 = io_x[19] ? _GEN253 : _GEN252;
wire  _GEN255 = io_x[23] ? _GEN254 : _GEN251;
wire  _GEN256 = io_x[27] ? _GEN255 : _GEN248;
wire  _GEN257 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN258 = io_x[19] ? _GEN257 : _GEN105;
wire  _GEN259 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN260 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN261 = io_x[19] ? _GEN260 : _GEN259;
wire  _GEN262 = io_x[23] ? _GEN261 : _GEN258;
wire  _GEN263 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN264 = io_x[19] ? _GEN263 : _GEN102;
wire  _GEN265 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN266 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN267 = io_x[19] ? _GEN266 : _GEN265;
wire  _GEN268 = io_x[23] ? _GEN267 : _GEN264;
wire  _GEN269 = io_x[27] ? _GEN268 : _GEN262;
wire  _GEN270 = io_x[48] ? _GEN269 : _GEN256;
wire  _GEN271 = io_x[31] ? _GEN270 : _GEN241;
wire  _GEN272 = io_x[3] ? _GEN271 : _GEN210;
wire  _GEN273 = io_x[5] ? _GEN272 : _GEN149;
wire  _GEN274 = 1'b1;
wire  _GEN275 = 1'b1;
wire  _GEN276 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN277 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN278 = io_x[19] ? _GEN277 : _GEN276;
wire  _GEN279 = io_x[23] ? _GEN278 : _GEN275;
wire  _GEN280 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN281 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN282 = io_x[19] ? _GEN281 : _GEN280;
wire  _GEN283 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN284 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN285 = io_x[19] ? _GEN284 : _GEN283;
wire  _GEN286 = io_x[23] ? _GEN285 : _GEN282;
wire  _GEN287 = io_x[27] ? _GEN286 : _GEN279;
wire  _GEN288 = io_x[48] ? _GEN287 : _GEN274;
wire  _GEN289 = 1'b0;
wire  _GEN290 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN291 = io_x[19] ? _GEN102 : _GEN290;
wire  _GEN292 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN293 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN294 = io_x[19] ? _GEN293 : _GEN292;
wire  _GEN295 = io_x[23] ? _GEN294 : _GEN291;
wire  _GEN296 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN297 = io_x[19] ? _GEN296 : _GEN105;
wire  _GEN298 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN299 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN300 = io_x[19] ? _GEN299 : _GEN298;
wire  _GEN301 = io_x[23] ? _GEN300 : _GEN297;
wire  _GEN302 = io_x[27] ? _GEN301 : _GEN295;
wire  _GEN303 = io_x[48] ? _GEN302 : _GEN289;
wire  _GEN304 = io_x[31] ? _GEN303 : _GEN288;
wire  _GEN305 = 1'b1;
wire  _GEN306 = 1'b0;
wire  _GEN307 = io_x[19] ? _GEN105 : _GEN102;
wire  _GEN308 = io_x[19] ? _GEN102 : _GEN105;
wire  _GEN309 = io_x[23] ? _GEN308 : _GEN307;
wire  _GEN310 = io_x[27] ? _GEN309 : _GEN306;
wire  _GEN311 = io_x[48] ? _GEN310 : _GEN274;
wire  _GEN312 = io_x[31] ? _GEN311 : _GEN305;
wire  _GEN313 = io_x[3] ? _GEN312 : _GEN304;
wire  _GEN314 = 1'b1;
wire  _GEN315 = io_x[19] ? _GEN105 : _GEN102;
wire  _GEN316 = io_x[23] ? _GEN315 : _GEN275;
wire  _GEN317 = io_x[27] ? _GEN316 : _GEN314;
wire  _GEN318 = io_x[48] ? _GEN317 : _GEN274;
wire  _GEN319 = 1'b0;
wire  _GEN320 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN321 = io_x[19] ? _GEN105 : _GEN320;
wire  _GEN322 = io_x[23] ? _GEN321 : _GEN319;
wire  _GEN323 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN324 = io_x[19] ? _GEN105 : _GEN323;
wire  _GEN325 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN326 = io_x[19] ? _GEN102 : _GEN325;
wire  _GEN327 = io_x[23] ? _GEN326 : _GEN324;
wire  _GEN328 = io_x[27] ? _GEN327 : _GEN322;
wire  _GEN329 = io_x[48] ? _GEN328 : _GEN274;
wire  _GEN330 = io_x[31] ? _GEN329 : _GEN318;
wire  _GEN331 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN332 = io_x[19] ? _GEN331 : _GEN105;
wire  _GEN333 = io_x[23] ? _GEN332 : _GEN275;
wire  _GEN334 = io_x[27] ? _GEN333 : _GEN314;
wire  _GEN335 = io_x[19] ? _GEN105 : _GEN102;
wire  _GEN336 = io_x[23] ? _GEN335 : _GEN275;
wire  _GEN337 = io_x[27] ? _GEN336 : _GEN314;
wire  _GEN338 = io_x[48] ? _GEN337 : _GEN334;
wire  _GEN339 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN340 = io_x[19] ? _GEN339 : _GEN105;
wire  _GEN341 = io_x[23] ? _GEN340 : _GEN275;
wire  _GEN342 = io_x[27] ? _GEN341 : _GEN314;
wire  _GEN343 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN344 = io_x[19] ? _GEN343 : _GEN102;
wire  _GEN345 = io_x[23] ? _GEN344 : _GEN275;
wire  _GEN346 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN347 = io_x[19] ? _GEN346 : _GEN102;
wire  _GEN348 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN349 = io_x[19] ? _GEN348 : _GEN105;
wire  _GEN350 = io_x[23] ? _GEN349 : _GEN347;
wire  _GEN351 = io_x[27] ? _GEN350 : _GEN345;
wire  _GEN352 = io_x[48] ? _GEN351 : _GEN342;
wire  _GEN353 = io_x[31] ? _GEN352 : _GEN338;
wire  _GEN354 = io_x[3] ? _GEN353 : _GEN330;
wire  _GEN355 = io_x[5] ? _GEN354 : _GEN313;
wire  _GEN356 = io_x[81] ? _GEN355 : _GEN273;
wire  _GEN357 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN358 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN359 = io_x[19] ? _GEN358 : _GEN357;
wire  _GEN360 = io_x[19] ? _GEN105 : _GEN102;
wire  _GEN361 = io_x[23] ? _GEN360 : _GEN359;
wire  _GEN362 = io_x[19] ? _GEN105 : _GEN102;
wire  _GEN363 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN364 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN365 = io_x[19] ? _GEN364 : _GEN363;
wire  _GEN366 = io_x[23] ? _GEN365 : _GEN362;
wire  _GEN367 = io_x[27] ? _GEN366 : _GEN361;
wire  _GEN368 = io_x[48] ? _GEN274 : _GEN367;
wire  _GEN369 = io_x[19] ? _GEN105 : _GEN102;
wire  _GEN370 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN371 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN372 = io_x[19] ? _GEN371 : _GEN370;
wire  _GEN373 = io_x[23] ? _GEN372 : _GEN369;
wire  _GEN374 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN375 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN376 = io_x[19] ? _GEN375 : _GEN374;
wire  _GEN377 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN378 = io_x[19] ? _GEN377 : _GEN102;
wire  _GEN379 = io_x[23] ? _GEN378 : _GEN376;
wire  _GEN380 = io_x[27] ? _GEN379 : _GEN373;
wire  _GEN381 = io_x[48] ? _GEN274 : _GEN380;
wire  _GEN382 = io_x[31] ? _GEN381 : _GEN368;
wire  _GEN383 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN384 = io_x[19] ? _GEN383 : _GEN105;
wire  _GEN385 = io_x[23] ? _GEN275 : _GEN384;
wire  _GEN386 = io_x[23] ? _GEN319 : _GEN275;
wire  _GEN387 = io_x[27] ? _GEN386 : _GEN385;
wire  _GEN388 = io_x[48] ? _GEN274 : _GEN387;
wire  _GEN389 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN390 = io_x[19] ? _GEN389 : _GEN105;
wire  _GEN391 = io_x[23] ? _GEN390 : _GEN275;
wire  _GEN392 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN393 = io_x[19] ? _GEN392 : _GEN102;
wire  _GEN394 = io_x[23] ? _GEN393 : _GEN319;
wire  _GEN395 = io_x[27] ? _GEN394 : _GEN391;
wire  _GEN396 = io_x[48] ? _GEN274 : _GEN395;
wire  _GEN397 = io_x[31] ? _GEN396 : _GEN388;
wire  _GEN398 = io_x[3] ? _GEN397 : _GEN382;
wire  _GEN399 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN400 = io_x[19] ? _GEN105 : _GEN399;
wire  _GEN401 = io_x[23] ? _GEN400 : _GEN275;
wire  _GEN402 = io_x[27] ? _GEN401 : _GEN314;
wire  _GEN403 = io_x[48] ? _GEN274 : _GEN402;
wire  _GEN404 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN405 = io_x[19] ? _GEN404 : _GEN102;
wire  _GEN406 = io_x[23] ? _GEN405 : _GEN275;
wire  _GEN407 = io_x[27] ? _GEN406 : _GEN306;
wire  _GEN408 = io_x[48] ? _GEN274 : _GEN407;
wire  _GEN409 = io_x[31] ? _GEN408 : _GEN403;
wire  _GEN410 = io_x[19] ? _GEN105 : _GEN102;
wire  _GEN411 = io_x[23] ? _GEN410 : _GEN275;
wire  _GEN412 = io_x[19] ? _GEN105 : _GEN102;
wire  _GEN413 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN414 = io_x[19] ? _GEN413 : _GEN105;
wire  _GEN415 = io_x[23] ? _GEN414 : _GEN412;
wire  _GEN416 = io_x[27] ? _GEN415 : _GEN411;
wire  _GEN417 = io_x[48] ? _GEN274 : _GEN416;
wire  _GEN418 = io_x[19] ? _GEN105 : _GEN102;
wire  _GEN419 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN420 = io_x[19] ? _GEN419 : _GEN102;
wire  _GEN421 = io_x[23] ? _GEN420 : _GEN418;
wire  _GEN422 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN423 = io_x[19] ? _GEN422 : _GEN105;
wire  _GEN424 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN425 = io_x[19] ? _GEN424 : _GEN102;
wire  _GEN426 = io_x[23] ? _GEN425 : _GEN423;
wire  _GEN427 = io_x[27] ? _GEN426 : _GEN421;
wire  _GEN428 = io_x[48] ? _GEN274 : _GEN427;
wire  _GEN429 = io_x[31] ? _GEN428 : _GEN417;
wire  _GEN430 = io_x[3] ? _GEN429 : _GEN409;
wire  _GEN431 = io_x[5] ? _GEN430 : _GEN398;
wire  _GEN432 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN433 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN434 = io_x[19] ? _GEN433 : _GEN432;
wire  _GEN435 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN436 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN437 = io_x[19] ? _GEN436 : _GEN435;
wire  _GEN438 = io_x[23] ? _GEN437 : _GEN434;
wire  _GEN439 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN440 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN441 = io_x[19] ? _GEN440 : _GEN439;
wire  _GEN442 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN443 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN444 = io_x[19] ? _GEN443 : _GEN442;
wire  _GEN445 = io_x[23] ? _GEN444 : _GEN441;
wire  _GEN446 = io_x[27] ? _GEN445 : _GEN438;
wire  _GEN447 = io_x[48] ? _GEN274 : _GEN446;
wire  _GEN448 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN449 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN450 = io_x[19] ? _GEN449 : _GEN448;
wire  _GEN451 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN452 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN453 = io_x[19] ? _GEN452 : _GEN451;
wire  _GEN454 = io_x[23] ? _GEN453 : _GEN450;
wire  _GEN455 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN456 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN457 = io_x[19] ? _GEN456 : _GEN455;
wire  _GEN458 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN459 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN460 = io_x[19] ? _GEN459 : _GEN458;
wire  _GEN461 = io_x[23] ? _GEN460 : _GEN457;
wire  _GEN462 = io_x[27] ? _GEN461 : _GEN454;
wire  _GEN463 = io_x[48] ? _GEN274 : _GEN462;
wire  _GEN464 = io_x[31] ? _GEN463 : _GEN447;
wire  _GEN465 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN466 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN467 = io_x[19] ? _GEN466 : _GEN465;
wire  _GEN468 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN469 = io_x[19] ? _GEN468 : _GEN102;
wire  _GEN470 = io_x[23] ? _GEN469 : _GEN467;
wire  _GEN471 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN472 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN473 = io_x[19] ? _GEN472 : _GEN471;
wire  _GEN474 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN475 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN476 = io_x[19] ? _GEN475 : _GEN474;
wire  _GEN477 = io_x[23] ? _GEN476 : _GEN473;
wire  _GEN478 = io_x[27] ? _GEN477 : _GEN470;
wire  _GEN479 = io_x[48] ? _GEN274 : _GEN478;
wire  _GEN480 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN481 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN482 = io_x[19] ? _GEN481 : _GEN480;
wire  _GEN483 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN484 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN485 = io_x[19] ? _GEN484 : _GEN483;
wire  _GEN486 = io_x[23] ? _GEN485 : _GEN482;
wire  _GEN487 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN488 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN489 = io_x[19] ? _GEN488 : _GEN487;
wire  _GEN490 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN491 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN492 = io_x[19] ? _GEN491 : _GEN490;
wire  _GEN493 = io_x[23] ? _GEN492 : _GEN489;
wire  _GEN494 = io_x[27] ? _GEN493 : _GEN486;
wire  _GEN495 = io_x[48] ? _GEN274 : _GEN494;
wire  _GEN496 = io_x[31] ? _GEN495 : _GEN479;
wire  _GEN497 = io_x[3] ? _GEN496 : _GEN464;
wire  _GEN498 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN499 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN500 = io_x[19] ? _GEN499 : _GEN498;
wire  _GEN501 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN502 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN503 = io_x[19] ? _GEN502 : _GEN501;
wire  _GEN504 = io_x[23] ? _GEN503 : _GEN500;
wire  _GEN505 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN506 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN507 = io_x[19] ? _GEN506 : _GEN505;
wire  _GEN508 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN509 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN510 = io_x[19] ? _GEN509 : _GEN508;
wire  _GEN511 = io_x[23] ? _GEN510 : _GEN507;
wire  _GEN512 = io_x[27] ? _GEN511 : _GEN504;
wire  _GEN513 = io_x[48] ? _GEN274 : _GEN512;
wire  _GEN514 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN515 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN516 = io_x[19] ? _GEN515 : _GEN514;
wire  _GEN517 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN518 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN519 = io_x[19] ? _GEN518 : _GEN517;
wire  _GEN520 = io_x[23] ? _GEN519 : _GEN516;
wire  _GEN521 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN522 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN523 = io_x[19] ? _GEN522 : _GEN521;
wire  _GEN524 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN525 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN526 = io_x[19] ? _GEN525 : _GEN524;
wire  _GEN527 = io_x[23] ? _GEN526 : _GEN523;
wire  _GEN528 = io_x[27] ? _GEN527 : _GEN520;
wire  _GEN529 = io_x[48] ? _GEN274 : _GEN528;
wire  _GEN530 = io_x[31] ? _GEN529 : _GEN513;
wire  _GEN531 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN532 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN533 = io_x[19] ? _GEN532 : _GEN531;
wire  _GEN534 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN535 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN536 = io_x[19] ? _GEN535 : _GEN534;
wire  _GEN537 = io_x[23] ? _GEN536 : _GEN533;
wire  _GEN538 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN539 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN540 = io_x[19] ? _GEN539 : _GEN538;
wire  _GEN541 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN542 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN543 = io_x[19] ? _GEN542 : _GEN541;
wire  _GEN544 = io_x[23] ? _GEN543 : _GEN540;
wire  _GEN545 = io_x[27] ? _GEN544 : _GEN537;
wire  _GEN546 = io_x[48] ? _GEN274 : _GEN545;
wire  _GEN547 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN548 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN549 = io_x[19] ? _GEN548 : _GEN547;
wire  _GEN550 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN551 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN552 = io_x[19] ? _GEN551 : _GEN550;
wire  _GEN553 = io_x[23] ? _GEN552 : _GEN549;
wire  _GEN554 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN555 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN556 = io_x[19] ? _GEN555 : _GEN554;
wire  _GEN557 = io_x[77] ? _GEN22 : _GEN23;
wire  _GEN558 = io_x[77] ? _GEN23 : _GEN22;
wire  _GEN559 = io_x[19] ? _GEN558 : _GEN557;
wire  _GEN560 = io_x[23] ? _GEN559 : _GEN556;
wire  _GEN561 = io_x[27] ? _GEN560 : _GEN553;
wire  _GEN562 = io_x[48] ? _GEN274 : _GEN561;
wire  _GEN563 = io_x[31] ? _GEN562 : _GEN546;
wire  _GEN564 = io_x[3] ? _GEN563 : _GEN530;
wire  _GEN565 = io_x[5] ? _GEN564 : _GEN497;
wire  _GEN566 = io_x[81] ? _GEN565 : _GEN431;
wire  _GEN567 = io_x[49] ? _GEN566 : _GEN356;
assign io_y[18] = _GEN567;
wire  _GEN568 = 1'b0;
wire  _GEN569 = 1'b1;
wire  _GEN570 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN571 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN572 = io_x[18] ? _GEN571 : _GEN570;
wire  _GEN573 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN574 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN575 = io_x[18] ? _GEN574 : _GEN573;
wire  _GEN576 = io_x[26] ? _GEN575 : _GEN572;
wire  _GEN577 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN578 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN579 = io_x[18] ? _GEN578 : _GEN577;
wire  _GEN580 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN581 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN582 = io_x[18] ? _GEN581 : _GEN580;
wire  _GEN583 = io_x[26] ? _GEN582 : _GEN579;
wire  _GEN584 = io_x[30] ? _GEN583 : _GEN576;
wire  _GEN585 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN586 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN587 = io_x[18] ? _GEN586 : _GEN585;
wire  _GEN588 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN589 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN590 = io_x[18] ? _GEN589 : _GEN588;
wire  _GEN591 = io_x[26] ? _GEN590 : _GEN587;
wire  _GEN592 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN593 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN594 = io_x[18] ? _GEN593 : _GEN592;
wire  _GEN595 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN596 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN597 = io_x[18] ? _GEN596 : _GEN595;
wire  _GEN598 = io_x[26] ? _GEN597 : _GEN594;
wire  _GEN599 = io_x[30] ? _GEN598 : _GEN591;
wire  _GEN600 = io_x[76] ? _GEN599 : _GEN584;
wire  _GEN601 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN602 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN603 = io_x[18] ? _GEN602 : _GEN601;
wire  _GEN604 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN605 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN606 = io_x[18] ? _GEN605 : _GEN604;
wire  _GEN607 = io_x[26] ? _GEN606 : _GEN603;
wire  _GEN608 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN609 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN610 = io_x[18] ? _GEN609 : _GEN608;
wire  _GEN611 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN612 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN613 = io_x[18] ? _GEN612 : _GEN611;
wire  _GEN614 = io_x[26] ? _GEN613 : _GEN610;
wire  _GEN615 = io_x[30] ? _GEN614 : _GEN607;
wire  _GEN616 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN617 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN618 = io_x[18] ? _GEN617 : _GEN616;
wire  _GEN619 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN620 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN621 = io_x[18] ? _GEN620 : _GEN619;
wire  _GEN622 = io_x[26] ? _GEN621 : _GEN618;
wire  _GEN623 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN624 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN625 = io_x[18] ? _GEN624 : _GEN623;
wire  _GEN626 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN627 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN628 = io_x[18] ? _GEN627 : _GEN626;
wire  _GEN629 = io_x[26] ? _GEN628 : _GEN625;
wire  _GEN630 = io_x[30] ? _GEN629 : _GEN622;
wire  _GEN631 = io_x[76] ? _GEN630 : _GEN615;
wire  _GEN632 = io_x[45] ? _GEN631 : _GEN600;
wire  _GEN633 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN634 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN635 = io_x[18] ? _GEN634 : _GEN633;
wire  _GEN636 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN637 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN638 = io_x[18] ? _GEN637 : _GEN636;
wire  _GEN639 = io_x[26] ? _GEN638 : _GEN635;
wire  _GEN640 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN641 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN642 = io_x[18] ? _GEN641 : _GEN640;
wire  _GEN643 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN644 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN645 = io_x[18] ? _GEN644 : _GEN643;
wire  _GEN646 = io_x[26] ? _GEN645 : _GEN642;
wire  _GEN647 = io_x[30] ? _GEN646 : _GEN639;
wire  _GEN648 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN649 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN650 = io_x[18] ? _GEN649 : _GEN648;
wire  _GEN651 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN652 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN653 = io_x[18] ? _GEN652 : _GEN651;
wire  _GEN654 = io_x[26] ? _GEN653 : _GEN650;
wire  _GEN655 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN656 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN657 = io_x[18] ? _GEN656 : _GEN655;
wire  _GEN658 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN659 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN660 = io_x[18] ? _GEN659 : _GEN658;
wire  _GEN661 = io_x[26] ? _GEN660 : _GEN657;
wire  _GEN662 = io_x[30] ? _GEN661 : _GEN654;
wire  _GEN663 = io_x[76] ? _GEN662 : _GEN647;
wire  _GEN664 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN665 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN666 = io_x[18] ? _GEN665 : _GEN664;
wire  _GEN667 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN668 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN669 = io_x[18] ? _GEN668 : _GEN667;
wire  _GEN670 = io_x[26] ? _GEN669 : _GEN666;
wire  _GEN671 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN672 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN673 = io_x[18] ? _GEN672 : _GEN671;
wire  _GEN674 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN675 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN676 = io_x[18] ? _GEN675 : _GEN674;
wire  _GEN677 = io_x[26] ? _GEN676 : _GEN673;
wire  _GEN678 = io_x[30] ? _GEN677 : _GEN670;
wire  _GEN679 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN680 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN681 = io_x[18] ? _GEN680 : _GEN679;
wire  _GEN682 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN683 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN684 = io_x[18] ? _GEN683 : _GEN682;
wire  _GEN685 = io_x[26] ? _GEN684 : _GEN681;
wire  _GEN686 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN687 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN688 = io_x[18] ? _GEN687 : _GEN686;
wire  _GEN689 = io_x[22] ? _GEN568 : _GEN569;
wire  _GEN690 = io_x[22] ? _GEN569 : _GEN568;
wire  _GEN691 = io_x[18] ? _GEN690 : _GEN689;
wire  _GEN692 = io_x[26] ? _GEN691 : _GEN688;
wire  _GEN693 = io_x[30] ? _GEN692 : _GEN685;
wire  _GEN694 = io_x[76] ? _GEN693 : _GEN678;
wire  _GEN695 = io_x[45] ? _GEN694 : _GEN663;
wire  _GEN696 = io_x[75] ? _GEN695 : _GEN632;
assign io_y[17] = _GEN696;
wire  _GEN697 = 1'b0;
wire  _GEN698 = 1'b1;
wire  _GEN699 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN700 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN701 = io_x[17] ? _GEN700 : _GEN699;
wire  _GEN702 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN703 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN704 = io_x[17] ? _GEN703 : _GEN702;
wire  _GEN705 = io_x[25] ? _GEN704 : _GEN701;
wire  _GEN706 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN707 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN708 = io_x[17] ? _GEN707 : _GEN706;
wire  _GEN709 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN710 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN711 = io_x[17] ? _GEN710 : _GEN709;
wire  _GEN712 = io_x[25] ? _GEN711 : _GEN708;
wire  _GEN713 = io_x[21] ? _GEN712 : _GEN705;
wire  _GEN714 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN715 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN716 = io_x[17] ? _GEN715 : _GEN714;
wire  _GEN717 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN718 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN719 = io_x[17] ? _GEN718 : _GEN717;
wire  _GEN720 = io_x[25] ? _GEN719 : _GEN716;
wire  _GEN721 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN722 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN723 = io_x[17] ? _GEN722 : _GEN721;
wire  _GEN724 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN725 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN726 = io_x[17] ? _GEN725 : _GEN724;
wire  _GEN727 = io_x[25] ? _GEN726 : _GEN723;
wire  _GEN728 = io_x[21] ? _GEN727 : _GEN720;
wire  _GEN729 = io_x[0] ? _GEN728 : _GEN713;
wire  _GEN730 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN731 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN732 = io_x[17] ? _GEN731 : _GEN730;
wire  _GEN733 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN734 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN735 = io_x[17] ? _GEN734 : _GEN733;
wire  _GEN736 = io_x[25] ? _GEN735 : _GEN732;
wire  _GEN737 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN738 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN739 = io_x[17] ? _GEN738 : _GEN737;
wire  _GEN740 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN741 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN742 = io_x[17] ? _GEN741 : _GEN740;
wire  _GEN743 = io_x[25] ? _GEN742 : _GEN739;
wire  _GEN744 = io_x[21] ? _GEN743 : _GEN736;
wire  _GEN745 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN746 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN747 = io_x[17] ? _GEN746 : _GEN745;
wire  _GEN748 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN749 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN750 = io_x[17] ? _GEN749 : _GEN748;
wire  _GEN751 = io_x[25] ? _GEN750 : _GEN747;
wire  _GEN752 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN753 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN754 = io_x[17] ? _GEN753 : _GEN752;
wire  _GEN755 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN756 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN757 = io_x[17] ? _GEN756 : _GEN755;
wire  _GEN758 = io_x[25] ? _GEN757 : _GEN754;
wire  _GEN759 = io_x[21] ? _GEN758 : _GEN751;
wire  _GEN760 = io_x[0] ? _GEN759 : _GEN744;
wire  _GEN761 = io_x[12] ? _GEN760 : _GEN729;
wire  _GEN762 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN763 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN764 = io_x[17] ? _GEN763 : _GEN762;
wire  _GEN765 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN766 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN767 = io_x[17] ? _GEN766 : _GEN765;
wire  _GEN768 = io_x[25] ? _GEN767 : _GEN764;
wire  _GEN769 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN770 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN771 = io_x[17] ? _GEN770 : _GEN769;
wire  _GEN772 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN773 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN774 = io_x[17] ? _GEN773 : _GEN772;
wire  _GEN775 = io_x[25] ? _GEN774 : _GEN771;
wire  _GEN776 = io_x[21] ? _GEN775 : _GEN768;
wire  _GEN777 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN778 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN779 = io_x[17] ? _GEN778 : _GEN777;
wire  _GEN780 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN781 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN782 = io_x[17] ? _GEN781 : _GEN780;
wire  _GEN783 = io_x[25] ? _GEN782 : _GEN779;
wire  _GEN784 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN785 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN786 = io_x[17] ? _GEN785 : _GEN784;
wire  _GEN787 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN788 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN789 = io_x[17] ? _GEN788 : _GEN787;
wire  _GEN790 = io_x[25] ? _GEN789 : _GEN786;
wire  _GEN791 = io_x[21] ? _GEN790 : _GEN783;
wire  _GEN792 = io_x[0] ? _GEN791 : _GEN776;
wire  _GEN793 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN794 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN795 = io_x[17] ? _GEN794 : _GEN793;
wire  _GEN796 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN797 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN798 = io_x[17] ? _GEN797 : _GEN796;
wire  _GEN799 = io_x[25] ? _GEN798 : _GEN795;
wire  _GEN800 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN801 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN802 = io_x[17] ? _GEN801 : _GEN800;
wire  _GEN803 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN804 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN805 = io_x[17] ? _GEN804 : _GEN803;
wire  _GEN806 = io_x[25] ? _GEN805 : _GEN802;
wire  _GEN807 = io_x[21] ? _GEN806 : _GEN799;
wire  _GEN808 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN809 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN810 = io_x[17] ? _GEN809 : _GEN808;
wire  _GEN811 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN812 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN813 = io_x[17] ? _GEN812 : _GEN811;
wire  _GEN814 = io_x[25] ? _GEN813 : _GEN810;
wire  _GEN815 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN816 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN817 = io_x[17] ? _GEN816 : _GEN815;
wire  _GEN818 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN819 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN820 = io_x[17] ? _GEN819 : _GEN818;
wire  _GEN821 = io_x[25] ? _GEN820 : _GEN817;
wire  _GEN822 = io_x[21] ? _GEN821 : _GEN814;
wire  _GEN823 = io_x[0] ? _GEN822 : _GEN807;
wire  _GEN824 = io_x[12] ? _GEN823 : _GEN792;
wire  _GEN825 = io_x[75] ? _GEN824 : _GEN761;
wire  _GEN826 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN827 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN828 = io_x[17] ? _GEN827 : _GEN826;
wire  _GEN829 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN830 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN831 = io_x[17] ? _GEN830 : _GEN829;
wire  _GEN832 = io_x[25] ? _GEN831 : _GEN828;
wire  _GEN833 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN834 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN835 = io_x[17] ? _GEN834 : _GEN833;
wire  _GEN836 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN837 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN838 = io_x[17] ? _GEN837 : _GEN836;
wire  _GEN839 = io_x[25] ? _GEN838 : _GEN835;
wire  _GEN840 = io_x[21] ? _GEN839 : _GEN832;
wire  _GEN841 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN842 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN843 = io_x[17] ? _GEN842 : _GEN841;
wire  _GEN844 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN845 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN846 = io_x[17] ? _GEN845 : _GEN844;
wire  _GEN847 = io_x[25] ? _GEN846 : _GEN843;
wire  _GEN848 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN849 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN850 = io_x[17] ? _GEN849 : _GEN848;
wire  _GEN851 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN852 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN853 = io_x[17] ? _GEN852 : _GEN851;
wire  _GEN854 = io_x[25] ? _GEN853 : _GEN850;
wire  _GEN855 = io_x[21] ? _GEN854 : _GEN847;
wire  _GEN856 = io_x[0] ? _GEN855 : _GEN840;
wire  _GEN857 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN858 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN859 = io_x[17] ? _GEN858 : _GEN857;
wire  _GEN860 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN861 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN862 = io_x[17] ? _GEN861 : _GEN860;
wire  _GEN863 = io_x[25] ? _GEN862 : _GEN859;
wire  _GEN864 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN865 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN866 = io_x[17] ? _GEN865 : _GEN864;
wire  _GEN867 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN868 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN869 = io_x[17] ? _GEN868 : _GEN867;
wire  _GEN870 = io_x[25] ? _GEN869 : _GEN866;
wire  _GEN871 = io_x[21] ? _GEN870 : _GEN863;
wire  _GEN872 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN873 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN874 = io_x[17] ? _GEN873 : _GEN872;
wire  _GEN875 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN876 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN877 = io_x[17] ? _GEN876 : _GEN875;
wire  _GEN878 = io_x[25] ? _GEN877 : _GEN874;
wire  _GEN879 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN880 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN881 = io_x[17] ? _GEN880 : _GEN879;
wire  _GEN882 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN883 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN884 = io_x[17] ? _GEN883 : _GEN882;
wire  _GEN885 = io_x[25] ? _GEN884 : _GEN881;
wire  _GEN886 = io_x[21] ? _GEN885 : _GEN878;
wire  _GEN887 = io_x[0] ? _GEN886 : _GEN871;
wire  _GEN888 = io_x[12] ? _GEN887 : _GEN856;
wire  _GEN889 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN890 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN891 = io_x[17] ? _GEN890 : _GEN889;
wire  _GEN892 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN893 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN894 = io_x[17] ? _GEN893 : _GEN892;
wire  _GEN895 = io_x[25] ? _GEN894 : _GEN891;
wire  _GEN896 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN897 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN898 = io_x[17] ? _GEN897 : _GEN896;
wire  _GEN899 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN900 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN901 = io_x[17] ? _GEN900 : _GEN899;
wire  _GEN902 = io_x[25] ? _GEN901 : _GEN898;
wire  _GEN903 = io_x[21] ? _GEN902 : _GEN895;
wire  _GEN904 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN905 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN906 = io_x[17] ? _GEN905 : _GEN904;
wire  _GEN907 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN908 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN909 = io_x[17] ? _GEN908 : _GEN907;
wire  _GEN910 = io_x[25] ? _GEN909 : _GEN906;
wire  _GEN911 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN912 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN913 = io_x[17] ? _GEN912 : _GEN911;
wire  _GEN914 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN915 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN916 = io_x[17] ? _GEN915 : _GEN914;
wire  _GEN917 = io_x[25] ? _GEN916 : _GEN913;
wire  _GEN918 = io_x[21] ? _GEN917 : _GEN910;
wire  _GEN919 = io_x[0] ? _GEN918 : _GEN903;
wire  _GEN920 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN921 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN922 = io_x[17] ? _GEN921 : _GEN920;
wire  _GEN923 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN924 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN925 = io_x[17] ? _GEN924 : _GEN923;
wire  _GEN926 = io_x[25] ? _GEN925 : _GEN922;
wire  _GEN927 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN928 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN929 = io_x[17] ? _GEN928 : _GEN927;
wire  _GEN930 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN931 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN932 = io_x[17] ? _GEN931 : _GEN930;
wire  _GEN933 = io_x[25] ? _GEN932 : _GEN929;
wire  _GEN934 = io_x[21] ? _GEN933 : _GEN926;
wire  _GEN935 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN936 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN937 = io_x[17] ? _GEN936 : _GEN935;
wire  _GEN938 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN939 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN940 = io_x[17] ? _GEN939 : _GEN938;
wire  _GEN941 = io_x[25] ? _GEN940 : _GEN937;
wire  _GEN942 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN943 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN944 = io_x[17] ? _GEN943 : _GEN942;
wire  _GEN945 = io_x[29] ? _GEN697 : _GEN698;
wire  _GEN946 = io_x[29] ? _GEN698 : _GEN697;
wire  _GEN947 = io_x[17] ? _GEN946 : _GEN945;
wire  _GEN948 = io_x[25] ? _GEN947 : _GEN944;
wire  _GEN949 = io_x[21] ? _GEN948 : _GEN941;
wire  _GEN950 = io_x[0] ? _GEN949 : _GEN934;
wire  _GEN951 = io_x[12] ? _GEN950 : _GEN919;
wire  _GEN952 = io_x[75] ? _GEN951 : _GEN888;
wire  _GEN953 = io_x[72] ? _GEN952 : _GEN825;
assign io_y[16] = _GEN953;
wire  _GEN954 = 1'b0;
wire  _GEN955 = 1'b1;
wire  _GEN956 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN957 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN958 = io_x[24] ? _GEN957 : _GEN956;
wire  _GEN959 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN960 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN961 = io_x[24] ? _GEN960 : _GEN959;
wire  _GEN962 = io_x[28] ? _GEN961 : _GEN958;
wire  _GEN963 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN964 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN965 = io_x[24] ? _GEN964 : _GEN963;
wire  _GEN966 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN967 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN968 = io_x[24] ? _GEN967 : _GEN966;
wire  _GEN969 = io_x[28] ? _GEN968 : _GEN965;
wire  _GEN970 = io_x[16] ? _GEN969 : _GEN962;
wire  _GEN971 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN972 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN973 = io_x[24] ? _GEN972 : _GEN971;
wire  _GEN974 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN975 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN976 = io_x[24] ? _GEN975 : _GEN974;
wire  _GEN977 = io_x[28] ? _GEN976 : _GEN973;
wire  _GEN978 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN979 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN980 = io_x[24] ? _GEN979 : _GEN978;
wire  _GEN981 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN982 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN983 = io_x[24] ? _GEN982 : _GEN981;
wire  _GEN984 = io_x[28] ? _GEN983 : _GEN980;
wire  _GEN985 = io_x[16] ? _GEN984 : _GEN977;
wire  _GEN986 = io_x[45] ? _GEN985 : _GEN970;
wire  _GEN987 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN988 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN989 = io_x[24] ? _GEN988 : _GEN987;
wire  _GEN990 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN991 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN992 = io_x[24] ? _GEN991 : _GEN990;
wire  _GEN993 = io_x[28] ? _GEN992 : _GEN989;
wire  _GEN994 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN995 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN996 = io_x[24] ? _GEN995 : _GEN994;
wire  _GEN997 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN998 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN999 = io_x[24] ? _GEN998 : _GEN997;
wire  _GEN1000 = io_x[28] ? _GEN999 : _GEN996;
wire  _GEN1001 = io_x[16] ? _GEN1000 : _GEN993;
wire  _GEN1002 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN1003 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN1004 = io_x[24] ? _GEN1003 : _GEN1002;
wire  _GEN1005 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN1006 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN1007 = io_x[24] ? _GEN1006 : _GEN1005;
wire  _GEN1008 = io_x[28] ? _GEN1007 : _GEN1004;
wire  _GEN1009 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN1010 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN1011 = io_x[24] ? _GEN1010 : _GEN1009;
wire  _GEN1012 = io_x[20] ? _GEN954 : _GEN955;
wire  _GEN1013 = io_x[20] ? _GEN955 : _GEN954;
wire  _GEN1014 = io_x[24] ? _GEN1013 : _GEN1012;
wire  _GEN1015 = io_x[28] ? _GEN1014 : _GEN1011;
wire  _GEN1016 = io_x[16] ? _GEN1015 : _GEN1008;
wire  _GEN1017 = io_x[45] ? _GEN1016 : _GEN1001;
wire  _GEN1018 = io_x[74] ? _GEN1017 : _GEN986;
assign io_y[15] = _GEN1018;
wire  _GEN1019 = 1'b0;
wire  _GEN1020 = 1'b1;
wire  _GEN1021 = io_x[73] ? _GEN1020 : _GEN1019;
wire  _GEN1022 = io_x[73] ? _GEN1020 : _GEN1019;
wire  _GEN1023 = io_x[45] ? _GEN1022 : _GEN1021;
wire  _GEN1024 = io_x[73] ? _GEN1020 : _GEN1019;
wire  _GEN1025 = io_x[73] ? _GEN1020 : _GEN1019;
wire  _GEN1026 = io_x[45] ? _GEN1025 : _GEN1024;
wire  _GEN1027 = io_x[15] ? _GEN1026 : _GEN1023;
assign io_y[14] = _GEN1027;
wire  _GEN1028 = 1'b0;
wire  _GEN1029 = 1'b1;
wire  _GEN1030 = io_x[72] ? _GEN1029 : _GEN1028;
wire  _GEN1031 = io_x[72] ? _GEN1029 : _GEN1028;
wire  _GEN1032 = io_x[17] ? _GEN1031 : _GEN1030;
wire  _GEN1033 = io_x[72] ? _GEN1029 : _GEN1028;
wire  _GEN1034 = io_x[72] ? _GEN1029 : _GEN1028;
wire  _GEN1035 = io_x[17] ? _GEN1034 : _GEN1033;
wire  _GEN1036 = io_x[39] ? _GEN1035 : _GEN1032;
wire  _GEN1037 = io_x[72] ? _GEN1029 : _GEN1028;
wire  _GEN1038 = io_x[72] ? _GEN1029 : _GEN1028;
wire  _GEN1039 = io_x[17] ? _GEN1038 : _GEN1037;
wire  _GEN1040 = io_x[72] ? _GEN1029 : _GEN1028;
wire  _GEN1041 = io_x[72] ? _GEN1029 : _GEN1028;
wire  _GEN1042 = io_x[17] ? _GEN1041 : _GEN1040;
wire  _GEN1043 = io_x[39] ? _GEN1042 : _GEN1039;
wire  _GEN1044 = io_x[19] ? _GEN1043 : _GEN1036;
assign io_y[13] = _GEN1044;
wire  _GEN1045 = 1'b0;
wire  _GEN1046 = 1'b1;
wire  _GEN1047 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1048 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1049 = io_x[39] ? _GEN1048 : _GEN1047;
wire  _GEN1050 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1051 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1052 = io_x[39] ? _GEN1051 : _GEN1050;
wire  _GEN1053 = io_x[74] ? _GEN1052 : _GEN1049;
wire  _GEN1054 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1055 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1056 = io_x[39] ? _GEN1055 : _GEN1054;
wire  _GEN1057 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1058 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1059 = io_x[39] ? _GEN1058 : _GEN1057;
wire  _GEN1060 = io_x[74] ? _GEN1059 : _GEN1056;
wire  _GEN1061 = io_x[81] ? _GEN1060 : _GEN1053;
wire  _GEN1062 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1063 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1064 = io_x[39] ? _GEN1063 : _GEN1062;
wire  _GEN1065 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1066 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1067 = io_x[39] ? _GEN1066 : _GEN1065;
wire  _GEN1068 = io_x[74] ? _GEN1067 : _GEN1064;
wire  _GEN1069 = 1'b0;
wire  _GEN1070 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1071 = io_x[39] ? _GEN1070 : _GEN1069;
wire  _GEN1072 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1073 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1074 = io_x[39] ? _GEN1073 : _GEN1072;
wire  _GEN1075 = io_x[74] ? _GEN1074 : _GEN1071;
wire  _GEN1076 = io_x[81] ? _GEN1075 : _GEN1068;
wire  _GEN1077 = io_x[75] ? _GEN1076 : _GEN1061;
wire  _GEN1078 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1079 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1080 = io_x[39] ? _GEN1079 : _GEN1078;
wire  _GEN1081 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1082 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1083 = io_x[39] ? _GEN1082 : _GEN1081;
wire  _GEN1084 = io_x[74] ? _GEN1083 : _GEN1080;
wire  _GEN1085 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1086 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1087 = io_x[39] ? _GEN1086 : _GEN1085;
wire  _GEN1088 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1089 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1090 = io_x[39] ? _GEN1089 : _GEN1088;
wire  _GEN1091 = io_x[74] ? _GEN1090 : _GEN1087;
wire  _GEN1092 = io_x[81] ? _GEN1091 : _GEN1084;
wire  _GEN1093 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1094 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1095 = io_x[39] ? _GEN1094 : _GEN1093;
wire  _GEN1096 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1097 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1098 = io_x[39] ? _GEN1097 : _GEN1096;
wire  _GEN1099 = io_x[74] ? _GEN1098 : _GEN1095;
wire  _GEN1100 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1101 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1102 = io_x[39] ? _GEN1101 : _GEN1100;
wire  _GEN1103 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1104 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1105 = io_x[39] ? _GEN1104 : _GEN1103;
wire  _GEN1106 = io_x[74] ? _GEN1105 : _GEN1102;
wire  _GEN1107 = io_x[81] ? _GEN1106 : _GEN1099;
wire  _GEN1108 = io_x[75] ? _GEN1107 : _GEN1092;
wire  _GEN1109 = io_x[43] ? _GEN1108 : _GEN1077;
wire  _GEN1110 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1111 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1112 = io_x[39] ? _GEN1111 : _GEN1110;
wire  _GEN1113 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1114 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1115 = io_x[39] ? _GEN1114 : _GEN1113;
wire  _GEN1116 = io_x[74] ? _GEN1115 : _GEN1112;
wire  _GEN1117 = 1'b1;
wire  _GEN1118 = io_x[39] ? _GEN1069 : _GEN1117;
wire  _GEN1119 = io_x[39] ? _GEN1069 : _GEN1117;
wire  _GEN1120 = io_x[74] ? _GEN1119 : _GEN1118;
wire  _GEN1121 = io_x[81] ? _GEN1120 : _GEN1116;
wire  _GEN1122 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1123 = io_x[39] ? _GEN1069 : _GEN1122;
wire  _GEN1124 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1125 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1126 = io_x[39] ? _GEN1125 : _GEN1124;
wire  _GEN1127 = io_x[74] ? _GEN1126 : _GEN1123;
wire  _GEN1128 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1129 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1130 = io_x[39] ? _GEN1129 : _GEN1128;
wire  _GEN1131 = 1'b1;
wire  _GEN1132 = io_x[74] ? _GEN1131 : _GEN1130;
wire  _GEN1133 = io_x[81] ? _GEN1132 : _GEN1127;
wire  _GEN1134 = io_x[75] ? _GEN1133 : _GEN1121;
wire  _GEN1135 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1136 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1137 = io_x[39] ? _GEN1136 : _GEN1135;
wire  _GEN1138 = io_x[39] ? _GEN1069 : _GEN1117;
wire  _GEN1139 = io_x[74] ? _GEN1138 : _GEN1137;
wire  _GEN1140 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1141 = io_x[39] ? _GEN1140 : _GEN1069;
wire  _GEN1142 = io_x[74] ? _GEN1131 : _GEN1141;
wire  _GEN1143 = io_x[81] ? _GEN1142 : _GEN1139;
wire  _GEN1144 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1145 = io_x[39] ? _GEN1144 : _GEN1069;
wire  _GEN1146 = io_x[74] ? _GEN1145 : _GEN1131;
wire  _GEN1147 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1148 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1149 = io_x[39] ? _GEN1148 : _GEN1147;
wire  _GEN1150 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1151 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1152 = io_x[39] ? _GEN1151 : _GEN1150;
wire  _GEN1153 = io_x[74] ? _GEN1152 : _GEN1149;
wire  _GEN1154 = io_x[81] ? _GEN1153 : _GEN1146;
wire  _GEN1155 = io_x[75] ? _GEN1154 : _GEN1143;
wire  _GEN1156 = io_x[43] ? _GEN1155 : _GEN1134;
wire  _GEN1157 = io_x[45] ? _GEN1156 : _GEN1109;
wire  _GEN1158 = 1'b1;
wire  _GEN1159 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1160 = io_x[39] ? _GEN1069 : _GEN1159;
wire  _GEN1161 = io_x[74] ? _GEN1160 : _GEN1131;
wire  _GEN1162 = io_x[81] ? _GEN1161 : _GEN1158;
wire  _GEN1163 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1164 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1165 = io_x[39] ? _GEN1164 : _GEN1163;
wire  _GEN1166 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1167 = io_x[39] ? _GEN1117 : _GEN1166;
wire  _GEN1168 = io_x[74] ? _GEN1167 : _GEN1165;
wire  _GEN1169 = io_x[81] ? _GEN1158 : _GEN1168;
wire  _GEN1170 = io_x[75] ? _GEN1169 : _GEN1162;
wire  _GEN1171 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1172 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1173 = io_x[39] ? _GEN1172 : _GEN1171;
wire  _GEN1174 = io_x[74] ? _GEN1131 : _GEN1173;
wire  _GEN1175 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1176 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1177 = io_x[39] ? _GEN1176 : _GEN1175;
wire  _GEN1178 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1179 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1180 = io_x[39] ? _GEN1179 : _GEN1178;
wire  _GEN1181 = io_x[74] ? _GEN1180 : _GEN1177;
wire  _GEN1182 = io_x[81] ? _GEN1181 : _GEN1174;
wire  _GEN1183 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1184 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1185 = io_x[39] ? _GEN1184 : _GEN1183;
wire  _GEN1186 = io_x[39] ? _GEN1069 : _GEN1117;
wire  _GEN1187 = io_x[74] ? _GEN1186 : _GEN1185;
wire  _GEN1188 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1189 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1190 = io_x[39] ? _GEN1189 : _GEN1188;
wire  _GEN1191 = io_x[74] ? _GEN1190 : _GEN1131;
wire  _GEN1192 = io_x[81] ? _GEN1191 : _GEN1187;
wire  _GEN1193 = io_x[75] ? _GEN1192 : _GEN1182;
wire  _GEN1194 = io_x[43] ? _GEN1193 : _GEN1170;
wire  _GEN1195 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1196 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1197 = io_x[39] ? _GEN1196 : _GEN1195;
wire  _GEN1198 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1199 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1200 = io_x[39] ? _GEN1199 : _GEN1198;
wire  _GEN1201 = io_x[74] ? _GEN1200 : _GEN1197;
wire  _GEN1202 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1203 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1204 = io_x[39] ? _GEN1203 : _GEN1202;
wire  _GEN1205 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1206 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1207 = io_x[39] ? _GEN1206 : _GEN1205;
wire  _GEN1208 = io_x[74] ? _GEN1207 : _GEN1204;
wire  _GEN1209 = io_x[81] ? _GEN1208 : _GEN1201;
wire  _GEN1210 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1211 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1212 = io_x[39] ? _GEN1211 : _GEN1210;
wire  _GEN1213 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1214 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1215 = io_x[39] ? _GEN1214 : _GEN1213;
wire  _GEN1216 = io_x[74] ? _GEN1215 : _GEN1212;
wire  _GEN1217 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1218 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1219 = io_x[39] ? _GEN1218 : _GEN1217;
wire  _GEN1220 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1221 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1222 = io_x[39] ? _GEN1221 : _GEN1220;
wire  _GEN1223 = io_x[74] ? _GEN1222 : _GEN1219;
wire  _GEN1224 = io_x[81] ? _GEN1223 : _GEN1216;
wire  _GEN1225 = io_x[75] ? _GEN1224 : _GEN1209;
wire  _GEN1226 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1227 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1228 = io_x[39] ? _GEN1227 : _GEN1226;
wire  _GEN1229 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1230 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1231 = io_x[39] ? _GEN1230 : _GEN1229;
wire  _GEN1232 = io_x[74] ? _GEN1231 : _GEN1228;
wire  _GEN1233 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1234 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1235 = io_x[39] ? _GEN1234 : _GEN1233;
wire  _GEN1236 = io_x[74] ? _GEN1131 : _GEN1235;
wire  _GEN1237 = io_x[81] ? _GEN1236 : _GEN1232;
wire  _GEN1238 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1239 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1240 = io_x[39] ? _GEN1239 : _GEN1238;
wire  _GEN1241 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1242 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1243 = io_x[39] ? _GEN1242 : _GEN1241;
wire  _GEN1244 = io_x[74] ? _GEN1243 : _GEN1240;
wire  _GEN1245 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1246 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1247 = io_x[39] ? _GEN1246 : _GEN1245;
wire  _GEN1248 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1249 = io_x[71] ? _GEN1046 : _GEN1045;
wire  _GEN1250 = io_x[39] ? _GEN1249 : _GEN1248;
wire  _GEN1251 = io_x[74] ? _GEN1250 : _GEN1247;
wire  _GEN1252 = io_x[81] ? _GEN1251 : _GEN1244;
wire  _GEN1253 = io_x[75] ? _GEN1252 : _GEN1237;
wire  _GEN1254 = io_x[43] ? _GEN1253 : _GEN1225;
wire  _GEN1255 = io_x[45] ? _GEN1254 : _GEN1194;
wire  _GEN1256 = io_x[77] ? _GEN1255 : _GEN1157;
assign io_y[12] = _GEN1256;
wire  _GEN1257 = 1'b0;
wire  _GEN1258 = 1'b1;
wire  _GEN1259 = io_x[70] ? _GEN1258 : _GEN1257;
wire  _GEN1260 = io_x[70] ? _GEN1258 : _GEN1257;
wire  _GEN1261 = io_x[78] ? _GEN1260 : _GEN1259;
wire  _GEN1262 = io_x[70] ? _GEN1258 : _GEN1257;
wire  _GEN1263 = io_x[70] ? _GEN1258 : _GEN1257;
wire  _GEN1264 = io_x[78] ? _GEN1263 : _GEN1262;
wire  _GEN1265 = io_x[41] ? _GEN1264 : _GEN1261;
assign io_y[11] = _GEN1265;
wire  _GEN1266 = 1'b0;
wire  _GEN1267 = 1'b1;
wire  _GEN1268 = io_x[69] ? _GEN1267 : _GEN1266;
wire  _GEN1269 = io_x[69] ? _GEN1267 : _GEN1266;
wire  _GEN1270 = io_x[43] ? _GEN1269 : _GEN1268;
assign io_y[10] = _GEN1270;
wire  _GEN1271 = 1'b0;
wire  _GEN1272 = 1'b1;
wire  _GEN1273 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1274 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1275 = io_x[7] ? _GEN1274 : _GEN1273;
wire  _GEN1276 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1277 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1278 = io_x[7] ? _GEN1277 : _GEN1276;
wire  _GEN1279 = io_x[11] ? _GEN1278 : _GEN1275;
wire  _GEN1280 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1281 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1282 = io_x[7] ? _GEN1281 : _GEN1280;
wire  _GEN1283 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1284 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1285 = io_x[7] ? _GEN1284 : _GEN1283;
wire  _GEN1286 = io_x[11] ? _GEN1285 : _GEN1282;
wire  _GEN1287 = io_x[3] ? _GEN1286 : _GEN1279;
wire  _GEN1288 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1289 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1290 = io_x[7] ? _GEN1289 : _GEN1288;
wire  _GEN1291 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1292 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1293 = io_x[7] ? _GEN1292 : _GEN1291;
wire  _GEN1294 = io_x[11] ? _GEN1293 : _GEN1290;
wire  _GEN1295 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1296 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1297 = io_x[7] ? _GEN1296 : _GEN1295;
wire  _GEN1298 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1299 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1300 = io_x[7] ? _GEN1299 : _GEN1298;
wire  _GEN1301 = io_x[11] ? _GEN1300 : _GEN1297;
wire  _GEN1302 = io_x[3] ? _GEN1301 : _GEN1294;
wire  _GEN1303 = io_x[77] ? _GEN1302 : _GEN1287;
wire  _GEN1304 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1305 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1306 = io_x[7] ? _GEN1305 : _GEN1304;
wire  _GEN1307 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1308 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1309 = io_x[7] ? _GEN1308 : _GEN1307;
wire  _GEN1310 = io_x[11] ? _GEN1309 : _GEN1306;
wire  _GEN1311 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1312 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1313 = io_x[7] ? _GEN1312 : _GEN1311;
wire  _GEN1314 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1315 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1316 = io_x[7] ? _GEN1315 : _GEN1314;
wire  _GEN1317 = io_x[11] ? _GEN1316 : _GEN1313;
wire  _GEN1318 = io_x[3] ? _GEN1317 : _GEN1310;
wire  _GEN1319 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1320 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1321 = io_x[7] ? _GEN1320 : _GEN1319;
wire  _GEN1322 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1323 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1324 = io_x[7] ? _GEN1323 : _GEN1322;
wire  _GEN1325 = io_x[11] ? _GEN1324 : _GEN1321;
wire  _GEN1326 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1327 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1328 = io_x[7] ? _GEN1327 : _GEN1326;
wire  _GEN1329 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1330 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1331 = io_x[7] ? _GEN1330 : _GEN1329;
wire  _GEN1332 = io_x[11] ? _GEN1331 : _GEN1328;
wire  _GEN1333 = io_x[3] ? _GEN1332 : _GEN1325;
wire  _GEN1334 = io_x[77] ? _GEN1333 : _GEN1318;
wire  _GEN1335 = io_x[15] ? _GEN1334 : _GEN1303;
wire  _GEN1336 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1337 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1338 = io_x[7] ? _GEN1337 : _GEN1336;
wire  _GEN1339 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1340 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1341 = io_x[7] ? _GEN1340 : _GEN1339;
wire  _GEN1342 = io_x[11] ? _GEN1341 : _GEN1338;
wire  _GEN1343 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1344 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1345 = io_x[7] ? _GEN1344 : _GEN1343;
wire  _GEN1346 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1347 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1348 = io_x[7] ? _GEN1347 : _GEN1346;
wire  _GEN1349 = io_x[11] ? _GEN1348 : _GEN1345;
wire  _GEN1350 = io_x[3] ? _GEN1349 : _GEN1342;
wire  _GEN1351 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1352 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1353 = io_x[7] ? _GEN1352 : _GEN1351;
wire  _GEN1354 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1355 = 1'b1;
wire  _GEN1356 = io_x[7] ? _GEN1355 : _GEN1354;
wire  _GEN1357 = io_x[11] ? _GEN1356 : _GEN1353;
wire  _GEN1358 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1359 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1360 = io_x[7] ? _GEN1359 : _GEN1358;
wire  _GEN1361 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1362 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1363 = io_x[7] ? _GEN1362 : _GEN1361;
wire  _GEN1364 = io_x[11] ? _GEN1363 : _GEN1360;
wire  _GEN1365 = io_x[3] ? _GEN1364 : _GEN1357;
wire  _GEN1366 = io_x[77] ? _GEN1365 : _GEN1350;
wire  _GEN1367 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1368 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1369 = io_x[7] ? _GEN1368 : _GEN1367;
wire  _GEN1370 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1371 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1372 = io_x[7] ? _GEN1371 : _GEN1370;
wire  _GEN1373 = io_x[11] ? _GEN1372 : _GEN1369;
wire  _GEN1374 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1375 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1376 = io_x[7] ? _GEN1375 : _GEN1374;
wire  _GEN1377 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1378 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1379 = io_x[7] ? _GEN1378 : _GEN1377;
wire  _GEN1380 = io_x[11] ? _GEN1379 : _GEN1376;
wire  _GEN1381 = io_x[3] ? _GEN1380 : _GEN1373;
wire  _GEN1382 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1383 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1384 = io_x[7] ? _GEN1383 : _GEN1382;
wire  _GEN1385 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1386 = io_x[7] ? _GEN1385 : _GEN1355;
wire  _GEN1387 = io_x[11] ? _GEN1386 : _GEN1384;
wire  _GEN1388 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1389 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1390 = io_x[7] ? _GEN1389 : _GEN1388;
wire  _GEN1391 = io_x[45] ? _GEN1271 : _GEN1272;
wire  _GEN1392 = io_x[45] ? _GEN1272 : _GEN1271;
wire  _GEN1393 = io_x[7] ? _GEN1392 : _GEN1391;
wire  _GEN1394 = io_x[11] ? _GEN1393 : _GEN1390;
wire  _GEN1395 = io_x[3] ? _GEN1394 : _GEN1387;
wire  _GEN1396 = io_x[77] ? _GEN1395 : _GEN1381;
wire  _GEN1397 = io_x[15] ? _GEN1396 : _GEN1366;
wire  _GEN1398 = io_x[34] ? _GEN1397 : _GEN1335;
assign io_y[9] = _GEN1398;
wire  _GEN1399 = 1'b0;
wire  _GEN1400 = 1'b1;
wire  _GEN1401 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1402 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1403 = io_x[6] ? _GEN1402 : _GEN1401;
wire  _GEN1404 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1405 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1406 = io_x[6] ? _GEN1405 : _GEN1404;
wire  _GEN1407 = io_x[2] ? _GEN1406 : _GEN1403;
wire  _GEN1408 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1409 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1410 = io_x[6] ? _GEN1409 : _GEN1408;
wire  _GEN1411 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1412 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1413 = io_x[6] ? _GEN1412 : _GEN1411;
wire  _GEN1414 = io_x[2] ? _GEN1413 : _GEN1410;
wire  _GEN1415 = io_x[14] ? _GEN1414 : _GEN1407;
wire  _GEN1416 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1417 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1418 = io_x[6] ? _GEN1417 : _GEN1416;
wire  _GEN1419 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1420 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1421 = io_x[6] ? _GEN1420 : _GEN1419;
wire  _GEN1422 = io_x[2] ? _GEN1421 : _GEN1418;
wire  _GEN1423 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1424 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1425 = io_x[6] ? _GEN1424 : _GEN1423;
wire  _GEN1426 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1427 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1428 = io_x[6] ? _GEN1427 : _GEN1426;
wire  _GEN1429 = io_x[2] ? _GEN1428 : _GEN1425;
wire  _GEN1430 = io_x[14] ? _GEN1429 : _GEN1422;
wire  _GEN1431 = io_x[44] ? _GEN1430 : _GEN1415;
wire  _GEN1432 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1433 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1434 = io_x[6] ? _GEN1433 : _GEN1432;
wire  _GEN1435 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1436 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1437 = io_x[6] ? _GEN1436 : _GEN1435;
wire  _GEN1438 = io_x[2] ? _GEN1437 : _GEN1434;
wire  _GEN1439 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1440 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1441 = io_x[6] ? _GEN1440 : _GEN1439;
wire  _GEN1442 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1443 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1444 = io_x[6] ? _GEN1443 : _GEN1442;
wire  _GEN1445 = io_x[2] ? _GEN1444 : _GEN1441;
wire  _GEN1446 = io_x[14] ? _GEN1445 : _GEN1438;
wire  _GEN1447 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1448 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1449 = io_x[6] ? _GEN1448 : _GEN1447;
wire  _GEN1450 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1451 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1452 = io_x[6] ? _GEN1451 : _GEN1450;
wire  _GEN1453 = io_x[2] ? _GEN1452 : _GEN1449;
wire  _GEN1454 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1455 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1456 = io_x[6] ? _GEN1455 : _GEN1454;
wire  _GEN1457 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1458 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1459 = io_x[6] ? _GEN1458 : _GEN1457;
wire  _GEN1460 = io_x[2] ? _GEN1459 : _GEN1456;
wire  _GEN1461 = io_x[14] ? _GEN1460 : _GEN1453;
wire  _GEN1462 = io_x[44] ? _GEN1461 : _GEN1446;
wire  _GEN1463 = io_x[75] ? _GEN1462 : _GEN1431;
wire  _GEN1464 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1465 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1466 = io_x[6] ? _GEN1465 : _GEN1464;
wire  _GEN1467 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1468 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1469 = io_x[6] ? _GEN1468 : _GEN1467;
wire  _GEN1470 = io_x[2] ? _GEN1469 : _GEN1466;
wire  _GEN1471 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1472 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1473 = io_x[6] ? _GEN1472 : _GEN1471;
wire  _GEN1474 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1475 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1476 = io_x[6] ? _GEN1475 : _GEN1474;
wire  _GEN1477 = io_x[2] ? _GEN1476 : _GEN1473;
wire  _GEN1478 = io_x[14] ? _GEN1477 : _GEN1470;
wire  _GEN1479 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1480 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1481 = io_x[6] ? _GEN1480 : _GEN1479;
wire  _GEN1482 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1483 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1484 = io_x[6] ? _GEN1483 : _GEN1482;
wire  _GEN1485 = io_x[2] ? _GEN1484 : _GEN1481;
wire  _GEN1486 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1487 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1488 = io_x[6] ? _GEN1487 : _GEN1486;
wire  _GEN1489 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1490 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1491 = io_x[6] ? _GEN1490 : _GEN1489;
wire  _GEN1492 = io_x[2] ? _GEN1491 : _GEN1488;
wire  _GEN1493 = io_x[14] ? _GEN1492 : _GEN1485;
wire  _GEN1494 = io_x[44] ? _GEN1493 : _GEN1478;
wire  _GEN1495 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1496 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1497 = io_x[6] ? _GEN1496 : _GEN1495;
wire  _GEN1498 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1499 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1500 = io_x[6] ? _GEN1499 : _GEN1498;
wire  _GEN1501 = io_x[2] ? _GEN1500 : _GEN1497;
wire  _GEN1502 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1503 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1504 = io_x[6] ? _GEN1503 : _GEN1502;
wire  _GEN1505 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1506 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1507 = io_x[6] ? _GEN1506 : _GEN1505;
wire  _GEN1508 = io_x[2] ? _GEN1507 : _GEN1504;
wire  _GEN1509 = io_x[14] ? _GEN1508 : _GEN1501;
wire  _GEN1510 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1511 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1512 = io_x[6] ? _GEN1511 : _GEN1510;
wire  _GEN1513 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1514 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1515 = io_x[6] ? _GEN1514 : _GEN1513;
wire  _GEN1516 = io_x[2] ? _GEN1515 : _GEN1512;
wire  _GEN1517 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1518 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1519 = io_x[6] ? _GEN1518 : _GEN1517;
wire  _GEN1520 = io_x[10] ? _GEN1399 : _GEN1400;
wire  _GEN1521 = io_x[10] ? _GEN1400 : _GEN1399;
wire  _GEN1522 = io_x[6] ? _GEN1521 : _GEN1520;
wire  _GEN1523 = io_x[2] ? _GEN1522 : _GEN1519;
wire  _GEN1524 = io_x[14] ? _GEN1523 : _GEN1516;
wire  _GEN1525 = io_x[44] ? _GEN1524 : _GEN1509;
wire  _GEN1526 = io_x[75] ? _GEN1525 : _GEN1494;
wire  _GEN1527 = io_x[20] ? _GEN1526 : _GEN1463;
assign io_y[8] = _GEN1527;
wire  _GEN1528 = 1'b1;
wire  _GEN1529 = 1'b0;
wire  _GEN1530 = 1'b1;
wire  _GEN1531 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1532 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1533 = io_x[1] ? _GEN1532 : _GEN1531;
wire  _GEN1534 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1535 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1536 = io_x[1] ? _GEN1535 : _GEN1534;
wire  _GEN1537 = io_x[9] ? _GEN1536 : _GEN1533;
wire  _GEN1538 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1539 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1540 = io_x[1] ? _GEN1539 : _GEN1538;
wire  _GEN1541 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1542 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1543 = io_x[1] ? _GEN1542 : _GEN1541;
wire  _GEN1544 = io_x[9] ? _GEN1543 : _GEN1540;
wire  _GEN1545 = io_x[13] ? _GEN1544 : _GEN1537;
wire  _GEN1546 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1547 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1548 = io_x[1] ? _GEN1547 : _GEN1546;
wire  _GEN1549 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1550 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1551 = io_x[1] ? _GEN1550 : _GEN1549;
wire  _GEN1552 = io_x[9] ? _GEN1551 : _GEN1548;
wire  _GEN1553 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1554 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1555 = io_x[1] ? _GEN1554 : _GEN1553;
wire  _GEN1556 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1557 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1558 = io_x[1] ? _GEN1557 : _GEN1556;
wire  _GEN1559 = io_x[9] ? _GEN1558 : _GEN1555;
wire  _GEN1560 = io_x[13] ? _GEN1559 : _GEN1552;
wire  _GEN1561 = io_x[2] ? _GEN1560 : _GEN1545;
wire  _GEN1562 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1563 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1564 = io_x[1] ? _GEN1563 : _GEN1562;
wire  _GEN1565 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1566 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1567 = io_x[1] ? _GEN1566 : _GEN1565;
wire  _GEN1568 = io_x[9] ? _GEN1567 : _GEN1564;
wire  _GEN1569 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1570 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1571 = io_x[1] ? _GEN1570 : _GEN1569;
wire  _GEN1572 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1573 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1574 = io_x[1] ? _GEN1573 : _GEN1572;
wire  _GEN1575 = io_x[9] ? _GEN1574 : _GEN1571;
wire  _GEN1576 = io_x[13] ? _GEN1575 : _GEN1568;
wire  _GEN1577 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1578 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1579 = io_x[1] ? _GEN1578 : _GEN1577;
wire  _GEN1580 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1581 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1582 = io_x[1] ? _GEN1581 : _GEN1580;
wire  _GEN1583 = io_x[9] ? _GEN1582 : _GEN1579;
wire  _GEN1584 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1585 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1586 = io_x[1] ? _GEN1585 : _GEN1584;
wire  _GEN1587 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1588 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1589 = io_x[1] ? _GEN1588 : _GEN1587;
wire  _GEN1590 = io_x[9] ? _GEN1589 : _GEN1586;
wire  _GEN1591 = io_x[13] ? _GEN1590 : _GEN1583;
wire  _GEN1592 = io_x[2] ? _GEN1591 : _GEN1576;
wire  _GEN1593 = io_x[81] ? _GEN1592 : _GEN1561;
wire  _GEN1594 = 1'b1;
wire  _GEN1595 = io_x[82] ? _GEN1594 : _GEN1593;
wire  _GEN1596 = 1'b1;
wire  _GEN1597 = io_x[83] ? _GEN1596 : _GEN1595;
wire  _GEN1598 = 1'b1;
wire  _GEN1599 = io_x[84] ? _GEN1598 : _GEN1597;
wire  _GEN1600 = 1'b1;
wire  _GEN1601 = io_x[85] ? _GEN1600 : _GEN1599;
wire  _GEN1602 = 1'b1;
wire  _GEN1603 = io_x[86] ? _GEN1602 : _GEN1601;
wire  _GEN1604 = 1'b1;
wire  _GEN1605 = io_x[87] ? _GEN1604 : _GEN1603;
wire  _GEN1606 = 1'b1;
wire  _GEN1607 = io_x[88] ? _GEN1606 : _GEN1605;
wire  _GEN1608 = 1'b1;
wire  _GEN1609 = io_x[89] ? _GEN1608 : _GEN1607;
wire  _GEN1610 = 1'b1;
wire  _GEN1611 = io_x[90] ? _GEN1610 : _GEN1609;
wire  _GEN1612 = 1'b1;
wire  _GEN1613 = io_x[91] ? _GEN1612 : _GEN1611;
wire  _GEN1614 = 1'b1;
wire  _GEN1615 = io_x[92] ? _GEN1614 : _GEN1613;
wire  _GEN1616 = 1'b1;
wire  _GEN1617 = io_x[93] ? _GEN1616 : _GEN1615;
wire  _GEN1618 = 1'b1;
wire  _GEN1619 = io_x[94] ? _GEN1618 : _GEN1617;
wire  _GEN1620 = 1'b1;
wire  _GEN1621 = io_x[95] ? _GEN1620 : _GEN1619;
wire  _GEN1622 = 1'b1;
wire  _GEN1623 = io_x[96] ? _GEN1622 : _GEN1621;
wire  _GEN1624 = 1'b1;
wire  _GEN1625 = io_x[97] ? _GEN1624 : _GEN1623;
wire  _GEN1626 = io_x[98] ? _GEN1625 : _GEN1528;
wire  _GEN1627 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1628 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1629 = io_x[1] ? _GEN1628 : _GEN1627;
wire  _GEN1630 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1631 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1632 = io_x[1] ? _GEN1631 : _GEN1630;
wire  _GEN1633 = io_x[9] ? _GEN1632 : _GEN1629;
wire  _GEN1634 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1635 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1636 = io_x[1] ? _GEN1635 : _GEN1634;
wire  _GEN1637 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1638 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1639 = io_x[1] ? _GEN1638 : _GEN1637;
wire  _GEN1640 = io_x[9] ? _GEN1639 : _GEN1636;
wire  _GEN1641 = io_x[13] ? _GEN1640 : _GEN1633;
wire  _GEN1642 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1643 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1644 = io_x[1] ? _GEN1643 : _GEN1642;
wire  _GEN1645 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1646 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1647 = io_x[1] ? _GEN1646 : _GEN1645;
wire  _GEN1648 = io_x[9] ? _GEN1647 : _GEN1644;
wire  _GEN1649 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1650 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1651 = io_x[1] ? _GEN1650 : _GEN1649;
wire  _GEN1652 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1653 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1654 = io_x[1] ? _GEN1653 : _GEN1652;
wire  _GEN1655 = io_x[9] ? _GEN1654 : _GEN1651;
wire  _GEN1656 = io_x[13] ? _GEN1655 : _GEN1648;
wire  _GEN1657 = io_x[2] ? _GEN1656 : _GEN1641;
wire  _GEN1658 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1659 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1660 = io_x[1] ? _GEN1659 : _GEN1658;
wire  _GEN1661 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1662 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1663 = io_x[1] ? _GEN1662 : _GEN1661;
wire  _GEN1664 = io_x[9] ? _GEN1663 : _GEN1660;
wire  _GEN1665 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1666 = 1'b1;
wire  _GEN1667 = io_x[1] ? _GEN1666 : _GEN1665;
wire  _GEN1668 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1669 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1670 = io_x[1] ? _GEN1669 : _GEN1668;
wire  _GEN1671 = io_x[9] ? _GEN1670 : _GEN1667;
wire  _GEN1672 = io_x[13] ? _GEN1671 : _GEN1664;
wire  _GEN1673 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1674 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1675 = io_x[1] ? _GEN1674 : _GEN1673;
wire  _GEN1676 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1677 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1678 = io_x[1] ? _GEN1677 : _GEN1676;
wire  _GEN1679 = io_x[9] ? _GEN1678 : _GEN1675;
wire  _GEN1680 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1681 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1682 = io_x[1] ? _GEN1681 : _GEN1680;
wire  _GEN1683 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1684 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1685 = io_x[1] ? _GEN1684 : _GEN1683;
wire  _GEN1686 = io_x[9] ? _GEN1685 : _GEN1682;
wire  _GEN1687 = io_x[13] ? _GEN1686 : _GEN1679;
wire  _GEN1688 = io_x[2] ? _GEN1687 : _GEN1672;
wire  _GEN1689 = io_x[81] ? _GEN1688 : _GEN1657;
wire  _GEN1690 = io_x[82] ? _GEN1594 : _GEN1689;
wire  _GEN1691 = io_x[83] ? _GEN1596 : _GEN1690;
wire  _GEN1692 = io_x[84] ? _GEN1598 : _GEN1691;
wire  _GEN1693 = io_x[85] ? _GEN1600 : _GEN1692;
wire  _GEN1694 = io_x[86] ? _GEN1602 : _GEN1693;
wire  _GEN1695 = io_x[87] ? _GEN1604 : _GEN1694;
wire  _GEN1696 = io_x[88] ? _GEN1606 : _GEN1695;
wire  _GEN1697 = io_x[89] ? _GEN1608 : _GEN1696;
wire  _GEN1698 = io_x[90] ? _GEN1610 : _GEN1697;
wire  _GEN1699 = io_x[91] ? _GEN1612 : _GEN1698;
wire  _GEN1700 = io_x[92] ? _GEN1614 : _GEN1699;
wire  _GEN1701 = io_x[93] ? _GEN1616 : _GEN1700;
wire  _GEN1702 = io_x[94] ? _GEN1618 : _GEN1701;
wire  _GEN1703 = io_x[95] ? _GEN1620 : _GEN1702;
wire  _GEN1704 = io_x[96] ? _GEN1622 : _GEN1703;
wire  _GEN1705 = io_x[97] ? _GEN1624 : _GEN1704;
wire  _GEN1706 = io_x[98] ? _GEN1705 : _GEN1528;
wire  _GEN1707 = io_x[43] ? _GEN1706 : _GEN1626;
wire  _GEN1708 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1709 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1710 = io_x[1] ? _GEN1709 : _GEN1708;
wire  _GEN1711 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1712 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1713 = io_x[1] ? _GEN1712 : _GEN1711;
wire  _GEN1714 = io_x[9] ? _GEN1713 : _GEN1710;
wire  _GEN1715 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1716 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1717 = io_x[1] ? _GEN1716 : _GEN1715;
wire  _GEN1718 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1719 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1720 = io_x[1] ? _GEN1719 : _GEN1718;
wire  _GEN1721 = io_x[9] ? _GEN1720 : _GEN1717;
wire  _GEN1722 = io_x[13] ? _GEN1721 : _GEN1714;
wire  _GEN1723 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1724 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1725 = io_x[1] ? _GEN1724 : _GEN1723;
wire  _GEN1726 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1727 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1728 = io_x[1] ? _GEN1727 : _GEN1726;
wire  _GEN1729 = io_x[9] ? _GEN1728 : _GEN1725;
wire  _GEN1730 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1731 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1732 = io_x[1] ? _GEN1731 : _GEN1730;
wire  _GEN1733 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1734 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1735 = io_x[1] ? _GEN1734 : _GEN1733;
wire  _GEN1736 = io_x[9] ? _GEN1735 : _GEN1732;
wire  _GEN1737 = io_x[13] ? _GEN1736 : _GEN1729;
wire  _GEN1738 = io_x[2] ? _GEN1737 : _GEN1722;
wire  _GEN1739 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1740 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1741 = io_x[1] ? _GEN1740 : _GEN1739;
wire  _GEN1742 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1743 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1744 = io_x[1] ? _GEN1743 : _GEN1742;
wire  _GEN1745 = io_x[9] ? _GEN1744 : _GEN1741;
wire  _GEN1746 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1747 = io_x[1] ? _GEN1666 : _GEN1746;
wire  _GEN1748 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1749 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1750 = io_x[1] ? _GEN1749 : _GEN1748;
wire  _GEN1751 = io_x[9] ? _GEN1750 : _GEN1747;
wire  _GEN1752 = io_x[13] ? _GEN1751 : _GEN1745;
wire  _GEN1753 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1754 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1755 = io_x[1] ? _GEN1754 : _GEN1753;
wire  _GEN1756 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1757 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1758 = io_x[1] ? _GEN1757 : _GEN1756;
wire  _GEN1759 = io_x[9] ? _GEN1758 : _GEN1755;
wire  _GEN1760 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1761 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1762 = io_x[1] ? _GEN1761 : _GEN1760;
wire  _GEN1763 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1764 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1765 = io_x[1] ? _GEN1764 : _GEN1763;
wire  _GEN1766 = io_x[9] ? _GEN1765 : _GEN1762;
wire  _GEN1767 = io_x[13] ? _GEN1766 : _GEN1759;
wire  _GEN1768 = io_x[2] ? _GEN1767 : _GEN1752;
wire  _GEN1769 = io_x[81] ? _GEN1768 : _GEN1738;
wire  _GEN1770 = io_x[82] ? _GEN1594 : _GEN1769;
wire  _GEN1771 = io_x[83] ? _GEN1596 : _GEN1770;
wire  _GEN1772 = io_x[84] ? _GEN1598 : _GEN1771;
wire  _GEN1773 = io_x[85] ? _GEN1600 : _GEN1772;
wire  _GEN1774 = io_x[86] ? _GEN1602 : _GEN1773;
wire  _GEN1775 = io_x[87] ? _GEN1604 : _GEN1774;
wire  _GEN1776 = io_x[88] ? _GEN1606 : _GEN1775;
wire  _GEN1777 = io_x[89] ? _GEN1608 : _GEN1776;
wire  _GEN1778 = io_x[90] ? _GEN1610 : _GEN1777;
wire  _GEN1779 = io_x[91] ? _GEN1612 : _GEN1778;
wire  _GEN1780 = io_x[92] ? _GEN1614 : _GEN1779;
wire  _GEN1781 = io_x[93] ? _GEN1616 : _GEN1780;
wire  _GEN1782 = io_x[94] ? _GEN1618 : _GEN1781;
wire  _GEN1783 = io_x[95] ? _GEN1620 : _GEN1782;
wire  _GEN1784 = io_x[96] ? _GEN1622 : _GEN1783;
wire  _GEN1785 = io_x[97] ? _GEN1624 : _GEN1784;
wire  _GEN1786 = io_x[98] ? _GEN1785 : _GEN1528;
wire  _GEN1787 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1788 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1789 = io_x[1] ? _GEN1788 : _GEN1787;
wire  _GEN1790 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1791 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1792 = io_x[1] ? _GEN1791 : _GEN1790;
wire  _GEN1793 = io_x[9] ? _GEN1792 : _GEN1789;
wire  _GEN1794 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1795 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1796 = io_x[1] ? _GEN1795 : _GEN1794;
wire  _GEN1797 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1798 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1799 = io_x[1] ? _GEN1798 : _GEN1797;
wire  _GEN1800 = io_x[9] ? _GEN1799 : _GEN1796;
wire  _GEN1801 = io_x[13] ? _GEN1800 : _GEN1793;
wire  _GEN1802 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1803 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1804 = io_x[1] ? _GEN1803 : _GEN1802;
wire  _GEN1805 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1806 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1807 = io_x[1] ? _GEN1806 : _GEN1805;
wire  _GEN1808 = io_x[9] ? _GEN1807 : _GEN1804;
wire  _GEN1809 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1810 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1811 = io_x[1] ? _GEN1810 : _GEN1809;
wire  _GEN1812 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1813 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1814 = io_x[1] ? _GEN1813 : _GEN1812;
wire  _GEN1815 = io_x[9] ? _GEN1814 : _GEN1811;
wire  _GEN1816 = io_x[13] ? _GEN1815 : _GEN1808;
wire  _GEN1817 = io_x[2] ? _GEN1816 : _GEN1801;
wire  _GEN1818 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1819 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1820 = io_x[1] ? _GEN1819 : _GEN1818;
wire  _GEN1821 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1822 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1823 = io_x[1] ? _GEN1822 : _GEN1821;
wire  _GEN1824 = io_x[9] ? _GEN1823 : _GEN1820;
wire  _GEN1825 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1826 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1827 = io_x[1] ? _GEN1826 : _GEN1825;
wire  _GEN1828 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1829 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1830 = io_x[1] ? _GEN1829 : _GEN1828;
wire  _GEN1831 = io_x[9] ? _GEN1830 : _GEN1827;
wire  _GEN1832 = io_x[13] ? _GEN1831 : _GEN1824;
wire  _GEN1833 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1834 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1835 = io_x[1] ? _GEN1834 : _GEN1833;
wire  _GEN1836 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1837 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1838 = io_x[1] ? _GEN1837 : _GEN1836;
wire  _GEN1839 = io_x[9] ? _GEN1838 : _GEN1835;
wire  _GEN1840 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1841 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1842 = io_x[1] ? _GEN1841 : _GEN1840;
wire  _GEN1843 = io_x[5] ? _GEN1529 : _GEN1530;
wire  _GEN1844 = io_x[5] ? _GEN1530 : _GEN1529;
wire  _GEN1845 = io_x[1] ? _GEN1844 : _GEN1843;
wire  _GEN1846 = io_x[9] ? _GEN1845 : _GEN1842;
wire  _GEN1847 = io_x[13] ? _GEN1846 : _GEN1839;
wire  _GEN1848 = io_x[2] ? _GEN1847 : _GEN1832;
wire  _GEN1849 = io_x[81] ? _GEN1848 : _GEN1817;
wire  _GEN1850 = io_x[82] ? _GEN1594 : _GEN1849;
wire  _GEN1851 = io_x[83] ? _GEN1596 : _GEN1850;
wire  _GEN1852 = io_x[84] ? _GEN1598 : _GEN1851;
wire  _GEN1853 = io_x[85] ? _GEN1600 : _GEN1852;
wire  _GEN1854 = io_x[86] ? _GEN1602 : _GEN1853;
wire  _GEN1855 = io_x[87] ? _GEN1604 : _GEN1854;
wire  _GEN1856 = io_x[88] ? _GEN1606 : _GEN1855;
wire  _GEN1857 = io_x[89] ? _GEN1608 : _GEN1856;
wire  _GEN1858 = io_x[90] ? _GEN1610 : _GEN1857;
wire  _GEN1859 = io_x[91] ? _GEN1612 : _GEN1858;
wire  _GEN1860 = io_x[92] ? _GEN1614 : _GEN1859;
wire  _GEN1861 = io_x[93] ? _GEN1616 : _GEN1860;
wire  _GEN1862 = io_x[94] ? _GEN1618 : _GEN1861;
wire  _GEN1863 = io_x[95] ? _GEN1620 : _GEN1862;
wire  _GEN1864 = io_x[96] ? _GEN1622 : _GEN1863;
wire  _GEN1865 = io_x[97] ? _GEN1624 : _GEN1864;
wire  _GEN1866 = io_x[98] ? _GEN1865 : _GEN1528;
wire  _GEN1867 = io_x[43] ? _GEN1866 : _GEN1786;
wire  _GEN1868 = io_x[40] ? _GEN1867 : _GEN1707;
assign io_y[7] = _GEN1868;
wire  _GEN1869 = 1'b0;
wire  _GEN1870 = 1'b1;
wire  _GEN1871 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1872 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1873 = io_x[42] ? _GEN1872 : _GEN1871;
wire  _GEN1874 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1875 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1876 = io_x[42] ? _GEN1875 : _GEN1874;
wire  _GEN1877 = io_x[44] ? _GEN1876 : _GEN1873;
wire  _GEN1878 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1879 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1880 = io_x[42] ? _GEN1879 : _GEN1878;
wire  _GEN1881 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1882 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1883 = io_x[42] ? _GEN1882 : _GEN1881;
wire  _GEN1884 = io_x[44] ? _GEN1883 : _GEN1880;
wire  _GEN1885 = io_x[3] ? _GEN1884 : _GEN1877;
wire  _GEN1886 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1887 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1888 = io_x[42] ? _GEN1887 : _GEN1886;
wire  _GEN1889 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1890 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1891 = io_x[42] ? _GEN1890 : _GEN1889;
wire  _GEN1892 = io_x[44] ? _GEN1891 : _GEN1888;
wire  _GEN1893 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1894 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1895 = io_x[42] ? _GEN1894 : _GEN1893;
wire  _GEN1896 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1897 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1898 = io_x[42] ? _GEN1897 : _GEN1896;
wire  _GEN1899 = io_x[44] ? _GEN1898 : _GEN1895;
wire  _GEN1900 = io_x[3] ? _GEN1899 : _GEN1892;
wire  _GEN1901 = io_x[8] ? _GEN1900 : _GEN1885;
wire  _GEN1902 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1903 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1904 = io_x[42] ? _GEN1903 : _GEN1902;
wire  _GEN1905 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1906 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1907 = io_x[42] ? _GEN1906 : _GEN1905;
wire  _GEN1908 = io_x[44] ? _GEN1907 : _GEN1904;
wire  _GEN1909 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1910 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1911 = io_x[42] ? _GEN1910 : _GEN1909;
wire  _GEN1912 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1913 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1914 = io_x[42] ? _GEN1913 : _GEN1912;
wire  _GEN1915 = io_x[44] ? _GEN1914 : _GEN1911;
wire  _GEN1916 = io_x[3] ? _GEN1915 : _GEN1908;
wire  _GEN1917 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1918 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1919 = io_x[42] ? _GEN1918 : _GEN1917;
wire  _GEN1920 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1921 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1922 = io_x[42] ? _GEN1921 : _GEN1920;
wire  _GEN1923 = io_x[44] ? _GEN1922 : _GEN1919;
wire  _GEN1924 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1925 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1926 = io_x[42] ? _GEN1925 : _GEN1924;
wire  _GEN1927 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1928 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1929 = io_x[42] ? _GEN1928 : _GEN1927;
wire  _GEN1930 = io_x[44] ? _GEN1929 : _GEN1926;
wire  _GEN1931 = io_x[3] ? _GEN1930 : _GEN1923;
wire  _GEN1932 = io_x[8] ? _GEN1931 : _GEN1916;
wire  _GEN1933 = io_x[4] ? _GEN1932 : _GEN1901;
wire  _GEN1934 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1935 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1936 = io_x[42] ? _GEN1935 : _GEN1934;
wire  _GEN1937 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1938 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1939 = io_x[42] ? _GEN1938 : _GEN1937;
wire  _GEN1940 = io_x[44] ? _GEN1939 : _GEN1936;
wire  _GEN1941 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1942 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1943 = io_x[42] ? _GEN1942 : _GEN1941;
wire  _GEN1944 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1945 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1946 = io_x[42] ? _GEN1945 : _GEN1944;
wire  _GEN1947 = io_x[44] ? _GEN1946 : _GEN1943;
wire  _GEN1948 = io_x[3] ? _GEN1947 : _GEN1940;
wire  _GEN1949 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1950 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1951 = io_x[42] ? _GEN1950 : _GEN1949;
wire  _GEN1952 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1953 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1954 = io_x[42] ? _GEN1953 : _GEN1952;
wire  _GEN1955 = io_x[44] ? _GEN1954 : _GEN1951;
wire  _GEN1956 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1957 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1958 = io_x[42] ? _GEN1957 : _GEN1956;
wire  _GEN1959 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1960 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1961 = io_x[42] ? _GEN1960 : _GEN1959;
wire  _GEN1962 = io_x[44] ? _GEN1961 : _GEN1958;
wire  _GEN1963 = io_x[3] ? _GEN1962 : _GEN1955;
wire  _GEN1964 = io_x[8] ? _GEN1963 : _GEN1948;
wire  _GEN1965 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1966 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1967 = io_x[42] ? _GEN1966 : _GEN1965;
wire  _GEN1968 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1969 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1970 = io_x[42] ? _GEN1969 : _GEN1968;
wire  _GEN1971 = io_x[44] ? _GEN1970 : _GEN1967;
wire  _GEN1972 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1973 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1974 = io_x[42] ? _GEN1973 : _GEN1972;
wire  _GEN1975 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1976 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1977 = io_x[42] ? _GEN1976 : _GEN1975;
wire  _GEN1978 = io_x[44] ? _GEN1977 : _GEN1974;
wire  _GEN1979 = io_x[3] ? _GEN1978 : _GEN1971;
wire  _GEN1980 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1981 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1982 = io_x[42] ? _GEN1981 : _GEN1980;
wire  _GEN1983 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1984 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1985 = io_x[42] ? _GEN1984 : _GEN1983;
wire  _GEN1986 = io_x[44] ? _GEN1985 : _GEN1982;
wire  _GEN1987 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1988 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1989 = io_x[42] ? _GEN1988 : _GEN1987;
wire  _GEN1990 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN1991 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1992 = io_x[42] ? _GEN1991 : _GEN1990;
wire  _GEN1993 = io_x[44] ? _GEN1992 : _GEN1989;
wire  _GEN1994 = io_x[3] ? _GEN1993 : _GEN1986;
wire  _GEN1995 = io_x[8] ? _GEN1994 : _GEN1979;
wire  _GEN1996 = io_x[4] ? _GEN1995 : _GEN1964;
wire  _GEN1997 = io_x[12] ? _GEN1996 : _GEN1933;
wire  _GEN1998 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN1999 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2000 = io_x[42] ? _GEN1999 : _GEN1998;
wire  _GEN2001 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2002 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2003 = io_x[42] ? _GEN2002 : _GEN2001;
wire  _GEN2004 = io_x[44] ? _GEN2003 : _GEN2000;
wire  _GEN2005 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2006 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2007 = io_x[42] ? _GEN2006 : _GEN2005;
wire  _GEN2008 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2009 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2010 = io_x[42] ? _GEN2009 : _GEN2008;
wire  _GEN2011 = io_x[44] ? _GEN2010 : _GEN2007;
wire  _GEN2012 = io_x[3] ? _GEN2011 : _GEN2004;
wire  _GEN2013 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2014 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2015 = io_x[42] ? _GEN2014 : _GEN2013;
wire  _GEN2016 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2017 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2018 = io_x[42] ? _GEN2017 : _GEN2016;
wire  _GEN2019 = io_x[44] ? _GEN2018 : _GEN2015;
wire  _GEN2020 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2021 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2022 = io_x[42] ? _GEN2021 : _GEN2020;
wire  _GEN2023 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2024 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2025 = io_x[42] ? _GEN2024 : _GEN2023;
wire  _GEN2026 = io_x[44] ? _GEN2025 : _GEN2022;
wire  _GEN2027 = io_x[3] ? _GEN2026 : _GEN2019;
wire  _GEN2028 = io_x[8] ? _GEN2027 : _GEN2012;
wire  _GEN2029 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2030 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2031 = io_x[42] ? _GEN2030 : _GEN2029;
wire  _GEN2032 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2033 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2034 = io_x[42] ? _GEN2033 : _GEN2032;
wire  _GEN2035 = io_x[44] ? _GEN2034 : _GEN2031;
wire  _GEN2036 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2037 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2038 = io_x[42] ? _GEN2037 : _GEN2036;
wire  _GEN2039 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2040 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2041 = io_x[42] ? _GEN2040 : _GEN2039;
wire  _GEN2042 = io_x[44] ? _GEN2041 : _GEN2038;
wire  _GEN2043 = io_x[3] ? _GEN2042 : _GEN2035;
wire  _GEN2044 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2045 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2046 = io_x[42] ? _GEN2045 : _GEN2044;
wire  _GEN2047 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2048 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2049 = io_x[42] ? _GEN2048 : _GEN2047;
wire  _GEN2050 = io_x[44] ? _GEN2049 : _GEN2046;
wire  _GEN2051 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2052 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2053 = io_x[42] ? _GEN2052 : _GEN2051;
wire  _GEN2054 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2055 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2056 = io_x[42] ? _GEN2055 : _GEN2054;
wire  _GEN2057 = io_x[44] ? _GEN2056 : _GEN2053;
wire  _GEN2058 = io_x[3] ? _GEN2057 : _GEN2050;
wire  _GEN2059 = io_x[8] ? _GEN2058 : _GEN2043;
wire  _GEN2060 = io_x[4] ? _GEN2059 : _GEN2028;
wire  _GEN2061 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2062 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2063 = io_x[42] ? _GEN2062 : _GEN2061;
wire  _GEN2064 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2065 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2066 = io_x[42] ? _GEN2065 : _GEN2064;
wire  _GEN2067 = io_x[44] ? _GEN2066 : _GEN2063;
wire  _GEN2068 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2069 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2070 = io_x[42] ? _GEN2069 : _GEN2068;
wire  _GEN2071 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2072 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2073 = io_x[42] ? _GEN2072 : _GEN2071;
wire  _GEN2074 = io_x[44] ? _GEN2073 : _GEN2070;
wire  _GEN2075 = io_x[3] ? _GEN2074 : _GEN2067;
wire  _GEN2076 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2077 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2078 = io_x[42] ? _GEN2077 : _GEN2076;
wire  _GEN2079 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2080 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2081 = io_x[42] ? _GEN2080 : _GEN2079;
wire  _GEN2082 = io_x[44] ? _GEN2081 : _GEN2078;
wire  _GEN2083 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2084 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2085 = io_x[42] ? _GEN2084 : _GEN2083;
wire  _GEN2086 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2087 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2088 = io_x[42] ? _GEN2087 : _GEN2086;
wire  _GEN2089 = io_x[44] ? _GEN2088 : _GEN2085;
wire  _GEN2090 = io_x[3] ? _GEN2089 : _GEN2082;
wire  _GEN2091 = io_x[8] ? _GEN2090 : _GEN2075;
wire  _GEN2092 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2093 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2094 = io_x[42] ? _GEN2093 : _GEN2092;
wire  _GEN2095 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2096 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2097 = io_x[42] ? _GEN2096 : _GEN2095;
wire  _GEN2098 = io_x[44] ? _GEN2097 : _GEN2094;
wire  _GEN2099 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2100 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2101 = io_x[42] ? _GEN2100 : _GEN2099;
wire  _GEN2102 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2103 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2104 = io_x[42] ? _GEN2103 : _GEN2102;
wire  _GEN2105 = io_x[44] ? _GEN2104 : _GEN2101;
wire  _GEN2106 = io_x[3] ? _GEN2105 : _GEN2098;
wire  _GEN2107 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2108 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2109 = io_x[42] ? _GEN2108 : _GEN2107;
wire  _GEN2110 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2111 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2112 = io_x[42] ? _GEN2111 : _GEN2110;
wire  _GEN2113 = io_x[44] ? _GEN2112 : _GEN2109;
wire  _GEN2114 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2115 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2116 = io_x[42] ? _GEN2115 : _GEN2114;
wire  _GEN2117 = io_x[0] ? _GEN1869 : _GEN1870;
wire  _GEN2118 = io_x[0] ? _GEN1870 : _GEN1869;
wire  _GEN2119 = io_x[42] ? _GEN2118 : _GEN2117;
wire  _GEN2120 = io_x[44] ? _GEN2119 : _GEN2116;
wire  _GEN2121 = io_x[3] ? _GEN2120 : _GEN2113;
wire  _GEN2122 = io_x[8] ? _GEN2121 : _GEN2106;
wire  _GEN2123 = io_x[4] ? _GEN2122 : _GEN2091;
wire  _GEN2124 = io_x[12] ? _GEN2123 : _GEN2060;
wire  _GEN2125 = io_x[34] ? _GEN2124 : _GEN1997;
assign io_y[6] = _GEN2125;
wire  _GEN2126 = 1'b0;
wire  _GEN2127 = 1'b1;
wire  _GEN2128 = io_x[41] ? _GEN2127 : _GEN2126;
wire  _GEN2129 = io_x[41] ? _GEN2127 : _GEN2126;
wire  _GEN2130 = io_x[42] ? _GEN2129 : _GEN2128;
wire  _GEN2131 = io_x[41] ? _GEN2127 : _GEN2126;
wire  _GEN2132 = io_x[41] ? _GEN2127 : _GEN2126;
wire  _GEN2133 = io_x[42] ? _GEN2132 : _GEN2131;
wire  _GEN2134 = io_x[15] ? _GEN2133 : _GEN2130;
assign io_y[5] = _GEN2134;
wire  _GEN2135 = 1'b0;
wire  _GEN2136 = 1'b1;
wire  _GEN2137 = io_x[40] ? _GEN2136 : _GEN2135;
wire  _GEN2138 = io_x[40] ? _GEN2136 : _GEN2135;
wire  _GEN2139 = io_x[78] ? _GEN2138 : _GEN2137;
wire  _GEN2140 = io_x[40] ? _GEN2136 : _GEN2135;
wire  _GEN2141 = io_x[40] ? _GEN2136 : _GEN2135;
wire  _GEN2142 = io_x[78] ? _GEN2141 : _GEN2140;
wire  _GEN2143 = io_x[39] ? _GEN2142 : _GEN2139;
assign io_y[4] = _GEN2143;
wire  _GEN2144 = 1'b0;
wire  _GEN2145 = 1'b1;
wire  _GEN2146 = io_x[39] ? _GEN2145 : _GEN2144;
wire  _GEN2147 = io_x[39] ? _GEN2145 : _GEN2144;
wire  _GEN2148 = io_x[70] ? _GEN2147 : _GEN2146;
assign io_y[3] = _GEN2148;
wire  _GEN2149 = 1'b0;
wire  _GEN2150 = 1'b1;
wire  _GEN2151 = io_x[38] ? _GEN2150 : _GEN2149;
wire  _GEN2152 = io_x[38] ? _GEN2150 : _GEN2149;
wire  _GEN2153 = io_x[1] ? _GEN2152 : _GEN2151;
wire  _GEN2154 = io_x[38] ? _GEN2150 : _GEN2149;
wire  _GEN2155 = io_x[38] ? _GEN2150 : _GEN2149;
wire  _GEN2156 = io_x[1] ? _GEN2155 : _GEN2154;
wire  _GEN2157 = io_x[43] ? _GEN2156 : _GEN2153;
wire  _GEN2158 = io_x[38] ? _GEN2150 : _GEN2149;
wire  _GEN2159 = io_x[38] ? _GEN2150 : _GEN2149;
wire  _GEN2160 = io_x[1] ? _GEN2159 : _GEN2158;
wire  _GEN2161 = io_x[38] ? _GEN2150 : _GEN2149;
wire  _GEN2162 = io_x[38] ? _GEN2150 : _GEN2149;
wire  _GEN2163 = io_x[1] ? _GEN2162 : _GEN2161;
wire  _GEN2164 = io_x[43] ? _GEN2163 : _GEN2160;
wire  _GEN2165 = io_x[45] ? _GEN2164 : _GEN2157;
assign io_y[2] = _GEN2165;
wire  _GEN2166 = 1'b0;
wire  _GEN2167 = 1'b1;
wire  _GEN2168 = io_x[37] ? _GEN2167 : _GEN2166;
wire  _GEN2169 = io_x[37] ? _GEN2167 : _GEN2166;
wire  _GEN2170 = io_x[70] ? _GEN2169 : _GEN2168;
assign io_y[1] = _GEN2170;
wire  _GEN2171 = 1'b0;
wire  _GEN2172 = 1'b1;
wire  _GEN2173 = io_x[34] ? _GEN2172 : _GEN2171;
wire  _GEN2174 = io_x[34] ? _GEN2172 : _GEN2171;
wire  _GEN2175 = io_x[77] ? _GEN2174 : _GEN2173;
assign io_y[0] = _GEN2175;
endmodule
