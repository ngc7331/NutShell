module BBGSharePredictorImp_BSD_c_NutShell_less(
    input [31:0] pc,
    input [31:0] train_pc,
    input  train_taken,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    input [15:0] train_ghr_rdata,
    output  taken,
    output  pht_wdata,
    output [8:0] pht_raddr,
    output [8:0] pht_waddr,
    output  ghr_wdata
);
wire [98:0] io_x;
wire [20:0] io_y;
assign io_x = { pc, train_pc, train_taken, pht_rdata, ghr_rdata, train_ghr_rdata };
assign { taken, pht_wdata, pht_raddr, pht_waddr, ghr_wdata } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[33] ? _GEN1 : _GEN0;
assign io_y[20] = _GEN2;
wire  _GEN3 = 1'b0;
wire  _GEN4 = 1'b1;
wire  _GEN5 = io_x[34] ? _GEN4 : _GEN3;
assign io_y[19] = _GEN5;
wire  _GEN6 = 1'b0;
wire  _GEN7 = 1'b1;
wire  _GEN8 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN9 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN10 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN11 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN12 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN13 = io_x[23] ? _GEN12 : _GEN11;
wire  _GEN14 = io_x[19] ? _GEN13 : _GEN10;
wire  _GEN15 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN16 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN17 = io_x[23] ? _GEN16 : _GEN15;
wire  _GEN18 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN19 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN20 = io_x[23] ? _GEN19 : _GEN18;
wire  _GEN21 = io_x[19] ? _GEN20 : _GEN17;
wire  _GEN22 = io_x[31] ? _GEN21 : _GEN14;
wire  _GEN23 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN24 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN25 = io_x[23] ? _GEN24 : _GEN23;
wire  _GEN26 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN27 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN28 = io_x[23] ? _GEN27 : _GEN26;
wire  _GEN29 = io_x[19] ? _GEN28 : _GEN25;
wire  _GEN30 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN31 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN32 = io_x[23] ? _GEN31 : _GEN30;
wire  _GEN33 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN34 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN35 = io_x[23] ? _GEN34 : _GEN33;
wire  _GEN36 = io_x[19] ? _GEN35 : _GEN32;
wire  _GEN37 = io_x[31] ? _GEN36 : _GEN29;
wire  _GEN38 = io_x[27] ? _GEN37 : _GEN22;
wire  _GEN39 = 1'b0;
wire  _GEN40 = 1'b1;
wire  _GEN41 = io_x[23] ? _GEN40 : _GEN39;
wire  _GEN42 = io_x[23] ? _GEN39 : _GEN40;
wire  _GEN43 = io_x[19] ? _GEN42 : _GEN41;
wire  _GEN44 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN45 = io_x[23] ? _GEN44 : _GEN40;
wire  _GEN46 = io_x[23] ? _GEN40 : _GEN39;
wire  _GEN47 = io_x[19] ? _GEN46 : _GEN45;
wire  _GEN48 = io_x[31] ? _GEN47 : _GEN43;
wire  _GEN49 = io_x[23] ? _GEN39 : _GEN40;
wire  _GEN50 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN51 = io_x[23] ? _GEN40 : _GEN50;
wire  _GEN52 = io_x[19] ? _GEN51 : _GEN49;
wire  _GEN53 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN54 = io_x[23] ? _GEN53 : _GEN39;
wire  _GEN55 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN56 = io_x[23] ? _GEN39 : _GEN55;
wire  _GEN57 = io_x[19] ? _GEN56 : _GEN54;
wire  _GEN58 = io_x[31] ? _GEN57 : _GEN52;
wire  _GEN59 = io_x[27] ? _GEN58 : _GEN48;
wire  _GEN60 = io_x[48] ? _GEN59 : _GEN38;
wire  _GEN61 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN62 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN63 = io_x[23] ? _GEN62 : _GEN61;
wire  _GEN64 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN65 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN66 = io_x[23] ? _GEN65 : _GEN64;
wire  _GEN67 = io_x[19] ? _GEN66 : _GEN63;
wire  _GEN68 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN69 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN70 = io_x[23] ? _GEN69 : _GEN68;
wire  _GEN71 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN72 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN73 = io_x[23] ? _GEN72 : _GEN71;
wire  _GEN74 = io_x[19] ? _GEN73 : _GEN70;
wire  _GEN75 = io_x[31] ? _GEN74 : _GEN67;
wire  _GEN76 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN77 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN78 = io_x[23] ? _GEN77 : _GEN76;
wire  _GEN79 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN80 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN81 = io_x[23] ? _GEN80 : _GEN79;
wire  _GEN82 = io_x[19] ? _GEN81 : _GEN78;
wire  _GEN83 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN84 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN85 = io_x[23] ? _GEN84 : _GEN83;
wire  _GEN86 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN87 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN88 = io_x[23] ? _GEN87 : _GEN86;
wire  _GEN89 = io_x[19] ? _GEN88 : _GEN85;
wire  _GEN90 = io_x[31] ? _GEN89 : _GEN82;
wire  _GEN91 = io_x[27] ? _GEN90 : _GEN75;
wire  _GEN92 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN93 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN94 = io_x[23] ? _GEN93 : _GEN92;
wire  _GEN95 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN96 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN97 = io_x[23] ? _GEN96 : _GEN95;
wire  _GEN98 = io_x[19] ? _GEN97 : _GEN94;
wire  _GEN99 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN100 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN101 = io_x[23] ? _GEN100 : _GEN99;
wire  _GEN102 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN103 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN104 = io_x[23] ? _GEN103 : _GEN102;
wire  _GEN105 = io_x[19] ? _GEN104 : _GEN101;
wire  _GEN106 = io_x[31] ? _GEN105 : _GEN98;
wire  _GEN107 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN108 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN109 = io_x[23] ? _GEN108 : _GEN107;
wire  _GEN110 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN111 = io_x[23] ? _GEN110 : _GEN40;
wire  _GEN112 = io_x[19] ? _GEN111 : _GEN109;
wire  _GEN113 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN114 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN115 = io_x[23] ? _GEN114 : _GEN113;
wire  _GEN116 = io_x[77] ? _GEN6 : _GEN7;
wire  _GEN117 = io_x[77] ? _GEN7 : _GEN6;
wire  _GEN118 = io_x[23] ? _GEN117 : _GEN116;
wire  _GEN119 = io_x[19] ? _GEN118 : _GEN115;
wire  _GEN120 = io_x[31] ? _GEN119 : _GEN112;
wire  _GEN121 = io_x[27] ? _GEN120 : _GEN106;
wire  _GEN122 = io_x[48] ? _GEN121 : _GEN91;
wire  _GEN123 = io_x[45] ? _GEN122 : _GEN60;
assign io_y[18] = _GEN123;
wire  _GEN124 = 1'b0;
wire  _GEN125 = 1'b1;
wire  _GEN126 = io_x[30] ? _GEN125 : _GEN124;
wire  _GEN127 = io_x[30] ? _GEN124 : _GEN125;
wire  _GEN128 = io_x[22] ? _GEN127 : _GEN126;
wire  _GEN129 = io_x[30] ? _GEN124 : _GEN125;
wire  _GEN130 = io_x[30] ? _GEN125 : _GEN124;
wire  _GEN131 = io_x[22] ? _GEN130 : _GEN129;
wire  _GEN132 = io_x[18] ? _GEN131 : _GEN128;
wire  _GEN133 = io_x[30] ? _GEN124 : _GEN125;
wire  _GEN134 = io_x[30] ? _GEN125 : _GEN124;
wire  _GEN135 = io_x[22] ? _GEN134 : _GEN133;
wire  _GEN136 = io_x[30] ? _GEN125 : _GEN124;
wire  _GEN137 = io_x[30] ? _GEN124 : _GEN125;
wire  _GEN138 = io_x[22] ? _GEN137 : _GEN136;
wire  _GEN139 = io_x[18] ? _GEN138 : _GEN135;
wire  _GEN140 = io_x[26] ? _GEN139 : _GEN132;
wire  _GEN141 = io_x[30] ? _GEN124 : _GEN125;
wire  _GEN142 = io_x[30] ? _GEN125 : _GEN124;
wire  _GEN143 = io_x[22] ? _GEN142 : _GEN141;
wire  _GEN144 = io_x[30] ? _GEN125 : _GEN124;
wire  _GEN145 = io_x[30] ? _GEN124 : _GEN125;
wire  _GEN146 = io_x[22] ? _GEN145 : _GEN144;
wire  _GEN147 = io_x[18] ? _GEN146 : _GEN143;
wire  _GEN148 = io_x[30] ? _GEN125 : _GEN124;
wire  _GEN149 = io_x[30] ? _GEN124 : _GEN125;
wire  _GEN150 = io_x[22] ? _GEN149 : _GEN148;
wire  _GEN151 = io_x[30] ? _GEN124 : _GEN125;
wire  _GEN152 = io_x[30] ? _GEN125 : _GEN124;
wire  _GEN153 = io_x[22] ? _GEN152 : _GEN151;
wire  _GEN154 = io_x[18] ? _GEN153 : _GEN150;
wire  _GEN155 = io_x[26] ? _GEN154 : _GEN147;
wire  _GEN156 = io_x[76] ? _GEN155 : _GEN140;
assign io_y[17] = _GEN156;
wire  _GEN157 = 1'b0;
wire  _GEN158 = 1'b1;
wire  _GEN159 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN160 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN161 = io_x[25] ? _GEN160 : _GEN159;
wire  _GEN162 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN163 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN164 = io_x[25] ? _GEN163 : _GEN162;
wire  _GEN165 = io_x[21] ? _GEN164 : _GEN161;
wire  _GEN166 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN167 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN168 = io_x[25] ? _GEN167 : _GEN166;
wire  _GEN169 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN170 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN171 = io_x[25] ? _GEN170 : _GEN169;
wire  _GEN172 = io_x[21] ? _GEN171 : _GEN168;
wire  _GEN173 = io_x[17] ? _GEN172 : _GEN165;
wire  _GEN174 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN175 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN176 = io_x[25] ? _GEN175 : _GEN174;
wire  _GEN177 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN178 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN179 = io_x[25] ? _GEN178 : _GEN177;
wire  _GEN180 = io_x[21] ? _GEN179 : _GEN176;
wire  _GEN181 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN182 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN183 = io_x[25] ? _GEN182 : _GEN181;
wire  _GEN184 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN185 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN186 = io_x[25] ? _GEN185 : _GEN184;
wire  _GEN187 = io_x[21] ? _GEN186 : _GEN183;
wire  _GEN188 = io_x[17] ? _GEN187 : _GEN180;
wire  _GEN189 = io_x[27] ? _GEN188 : _GEN173;
wire  _GEN190 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN191 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN192 = io_x[25] ? _GEN191 : _GEN190;
wire  _GEN193 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN194 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN195 = io_x[25] ? _GEN194 : _GEN193;
wire  _GEN196 = io_x[21] ? _GEN195 : _GEN192;
wire  _GEN197 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN198 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN199 = io_x[25] ? _GEN198 : _GEN197;
wire  _GEN200 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN201 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN202 = io_x[25] ? _GEN201 : _GEN200;
wire  _GEN203 = io_x[21] ? _GEN202 : _GEN199;
wire  _GEN204 = io_x[17] ? _GEN203 : _GEN196;
wire  _GEN205 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN206 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN207 = io_x[25] ? _GEN206 : _GEN205;
wire  _GEN208 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN209 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN210 = io_x[25] ? _GEN209 : _GEN208;
wire  _GEN211 = io_x[21] ? _GEN210 : _GEN207;
wire  _GEN212 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN213 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN214 = io_x[25] ? _GEN213 : _GEN212;
wire  _GEN215 = io_x[29] ? _GEN157 : _GEN158;
wire  _GEN216 = io_x[29] ? _GEN158 : _GEN157;
wire  _GEN217 = io_x[25] ? _GEN216 : _GEN215;
wire  _GEN218 = io_x[21] ? _GEN217 : _GEN214;
wire  _GEN219 = io_x[17] ? _GEN218 : _GEN211;
wire  _GEN220 = io_x[27] ? _GEN219 : _GEN204;
wire  _GEN221 = io_x[75] ? _GEN220 : _GEN189;
assign io_y[16] = _GEN221;
wire  _GEN222 = 1'b0;
wire  _GEN223 = 1'b1;
wire  _GEN224 = io_x[20] ? _GEN223 : _GEN222;
wire  _GEN225 = io_x[20] ? _GEN222 : _GEN223;
wire  _GEN226 = io_x[28] ? _GEN225 : _GEN224;
wire  _GEN227 = io_x[20] ? _GEN222 : _GEN223;
wire  _GEN228 = io_x[20] ? _GEN223 : _GEN222;
wire  _GEN229 = io_x[28] ? _GEN228 : _GEN227;
wire  _GEN230 = io_x[16] ? _GEN229 : _GEN226;
wire  _GEN231 = io_x[20] ? _GEN222 : _GEN223;
wire  _GEN232 = io_x[20] ? _GEN223 : _GEN222;
wire  _GEN233 = io_x[28] ? _GEN232 : _GEN231;
wire  _GEN234 = io_x[20] ? _GEN223 : _GEN222;
wire  _GEN235 = io_x[20] ? _GEN222 : _GEN223;
wire  _GEN236 = io_x[28] ? _GEN235 : _GEN234;
wire  _GEN237 = io_x[16] ? _GEN236 : _GEN233;
wire  _GEN238 = io_x[24] ? _GEN237 : _GEN230;
wire  _GEN239 = io_x[20] ? _GEN222 : _GEN223;
wire  _GEN240 = io_x[20] ? _GEN223 : _GEN222;
wire  _GEN241 = io_x[28] ? _GEN240 : _GEN239;
wire  _GEN242 = io_x[20] ? _GEN223 : _GEN222;
wire  _GEN243 = io_x[20] ? _GEN222 : _GEN223;
wire  _GEN244 = io_x[28] ? _GEN243 : _GEN242;
wire  _GEN245 = io_x[16] ? _GEN244 : _GEN241;
wire  _GEN246 = io_x[20] ? _GEN223 : _GEN222;
wire  _GEN247 = io_x[20] ? _GEN222 : _GEN223;
wire  _GEN248 = io_x[28] ? _GEN247 : _GEN246;
wire  _GEN249 = io_x[20] ? _GEN222 : _GEN223;
wire  _GEN250 = io_x[20] ? _GEN223 : _GEN222;
wire  _GEN251 = io_x[28] ? _GEN250 : _GEN249;
wire  _GEN252 = io_x[16] ? _GEN251 : _GEN248;
wire  _GEN253 = io_x[24] ? _GEN252 : _GEN245;
wire  _GEN254 = io_x[74] ? _GEN253 : _GEN238;
assign io_y[15] = _GEN254;
wire  _GEN255 = 1'b0;
wire  _GEN256 = 1'b1;
wire  _GEN257 = io_x[73] ? _GEN256 : _GEN255;
assign io_y[14] = _GEN257;
wire  _GEN258 = 1'b0;
wire  _GEN259 = 1'b1;
wire  _GEN260 = io_x[72] ? _GEN259 : _GEN258;
assign io_y[13] = _GEN260;
wire  _GEN261 = 1'b0;
wire  _GEN262 = 1'b1;
wire  _GEN263 = io_x[71] ? _GEN262 : _GEN261;
assign io_y[12] = _GEN263;
wire  _GEN264 = 1'b0;
wire  _GEN265 = 1'b1;
wire  _GEN266 = io_x[70] ? _GEN265 : _GEN264;
assign io_y[11] = _GEN266;
wire  _GEN267 = 1'b0;
wire  _GEN268 = 1'b1;
wire  _GEN269 = io_x[69] ? _GEN268 : _GEN267;
assign io_y[10] = _GEN269;
wire  _GEN270 = 1'b0;
wire  _GEN271 = 1'b1;
wire  _GEN272 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN273 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN274 = io_x[15] ? _GEN273 : _GEN272;
wire  _GEN275 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN276 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN277 = io_x[15] ? _GEN276 : _GEN275;
wire  _GEN278 = io_x[7] ? _GEN277 : _GEN274;
wire  _GEN279 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN280 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN281 = io_x[15] ? _GEN280 : _GEN279;
wire  _GEN282 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN283 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN284 = io_x[15] ? _GEN283 : _GEN282;
wire  _GEN285 = io_x[7] ? _GEN284 : _GEN281;
wire  _GEN286 = io_x[3] ? _GEN285 : _GEN278;
wire  _GEN287 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN288 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN289 = io_x[15] ? _GEN288 : _GEN287;
wire  _GEN290 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN291 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN292 = io_x[15] ? _GEN291 : _GEN290;
wire  _GEN293 = io_x[7] ? _GEN292 : _GEN289;
wire  _GEN294 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN295 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN296 = io_x[15] ? _GEN295 : _GEN294;
wire  _GEN297 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN298 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN299 = io_x[15] ? _GEN298 : _GEN297;
wire  _GEN300 = io_x[7] ? _GEN299 : _GEN296;
wire  _GEN301 = io_x[3] ? _GEN300 : _GEN293;
wire  _GEN302 = io_x[0] ? _GEN301 : _GEN286;
wire  _GEN303 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN304 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN305 = io_x[15] ? _GEN304 : _GEN303;
wire  _GEN306 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN307 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN308 = io_x[15] ? _GEN307 : _GEN306;
wire  _GEN309 = io_x[7] ? _GEN308 : _GEN305;
wire  _GEN310 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN311 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN312 = io_x[15] ? _GEN311 : _GEN310;
wire  _GEN313 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN314 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN315 = io_x[15] ? _GEN314 : _GEN313;
wire  _GEN316 = io_x[7] ? _GEN315 : _GEN312;
wire  _GEN317 = io_x[3] ? _GEN316 : _GEN309;
wire  _GEN318 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN319 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN320 = io_x[15] ? _GEN319 : _GEN318;
wire  _GEN321 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN322 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN323 = io_x[15] ? _GEN322 : _GEN321;
wire  _GEN324 = io_x[7] ? _GEN323 : _GEN320;
wire  _GEN325 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN326 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN327 = io_x[15] ? _GEN326 : _GEN325;
wire  _GEN328 = io_x[11] ? _GEN270 : _GEN271;
wire  _GEN329 = io_x[11] ? _GEN271 : _GEN270;
wire  _GEN330 = io_x[15] ? _GEN329 : _GEN328;
wire  _GEN331 = io_x[7] ? _GEN330 : _GEN327;
wire  _GEN332 = io_x[3] ? _GEN331 : _GEN324;
wire  _GEN333 = io_x[0] ? _GEN332 : _GEN317;
wire  _GEN334 = io_x[45] ? _GEN333 : _GEN302;
assign io_y[9] = _GEN334;
wire  _GEN335 = 1'b0;
wire  _GEN336 = 1'b1;
wire  _GEN337 = io_x[10] ? _GEN336 : _GEN335;
wire  _GEN338 = io_x[10] ? _GEN335 : _GEN336;
wire  _GEN339 = io_x[14] ? _GEN338 : _GEN337;
wire  _GEN340 = io_x[10] ? _GEN335 : _GEN336;
wire  _GEN341 = io_x[10] ? _GEN336 : _GEN335;
wire  _GEN342 = io_x[14] ? _GEN341 : _GEN340;
wire  _GEN343 = io_x[6] ? _GEN342 : _GEN339;
wire  _GEN344 = io_x[10] ? _GEN335 : _GEN336;
wire  _GEN345 = io_x[10] ? _GEN336 : _GEN335;
wire  _GEN346 = io_x[14] ? _GEN345 : _GEN344;
wire  _GEN347 = io_x[10] ? _GEN336 : _GEN335;
wire  _GEN348 = io_x[10] ? _GEN335 : _GEN336;
wire  _GEN349 = io_x[14] ? _GEN348 : _GEN347;
wire  _GEN350 = io_x[6] ? _GEN349 : _GEN346;
wire  _GEN351 = io_x[2] ? _GEN350 : _GEN343;
wire  _GEN352 = io_x[10] ? _GEN335 : _GEN336;
wire  _GEN353 = io_x[10] ? _GEN336 : _GEN335;
wire  _GEN354 = io_x[14] ? _GEN353 : _GEN352;
wire  _GEN355 = io_x[10] ? _GEN336 : _GEN335;
wire  _GEN356 = io_x[10] ? _GEN335 : _GEN336;
wire  _GEN357 = io_x[14] ? _GEN356 : _GEN355;
wire  _GEN358 = io_x[6] ? _GEN357 : _GEN354;
wire  _GEN359 = io_x[10] ? _GEN336 : _GEN335;
wire  _GEN360 = io_x[10] ? _GEN335 : _GEN336;
wire  _GEN361 = io_x[14] ? _GEN360 : _GEN359;
wire  _GEN362 = io_x[10] ? _GEN335 : _GEN336;
wire  _GEN363 = io_x[10] ? _GEN336 : _GEN335;
wire  _GEN364 = io_x[14] ? _GEN363 : _GEN362;
wire  _GEN365 = io_x[6] ? _GEN364 : _GEN361;
wire  _GEN366 = io_x[2] ? _GEN365 : _GEN358;
wire  _GEN367 = io_x[44] ? _GEN366 : _GEN351;
assign io_y[8] = _GEN367;
wire  _GEN368 = 1'b0;
wire  _GEN369 = 1'b1;
wire  _GEN370 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN371 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN372 = io_x[1] ? _GEN371 : _GEN370;
wire  _GEN373 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN374 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN375 = io_x[1] ? _GEN374 : _GEN373;
wire  _GEN376 = io_x[9] ? _GEN375 : _GEN372;
wire  _GEN377 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN378 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN379 = io_x[1] ? _GEN378 : _GEN377;
wire  _GEN380 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN381 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN382 = io_x[1] ? _GEN381 : _GEN380;
wire  _GEN383 = io_x[9] ? _GEN382 : _GEN379;
wire  _GEN384 = io_x[13] ? _GEN383 : _GEN376;
wire  _GEN385 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN386 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN387 = io_x[1] ? _GEN386 : _GEN385;
wire  _GEN388 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN389 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN390 = io_x[1] ? _GEN389 : _GEN388;
wire  _GEN391 = io_x[9] ? _GEN390 : _GEN387;
wire  _GEN392 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN393 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN394 = io_x[1] ? _GEN393 : _GEN392;
wire  _GEN395 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN396 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN397 = io_x[1] ? _GEN396 : _GEN395;
wire  _GEN398 = io_x[9] ? _GEN397 : _GEN394;
wire  _GEN399 = io_x[13] ? _GEN398 : _GEN391;
wire  _GEN400 = io_x[0] ? _GEN399 : _GEN384;
wire  _GEN401 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN402 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN403 = io_x[1] ? _GEN402 : _GEN401;
wire  _GEN404 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN405 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN406 = io_x[1] ? _GEN405 : _GEN404;
wire  _GEN407 = io_x[9] ? _GEN406 : _GEN403;
wire  _GEN408 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN409 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN410 = io_x[1] ? _GEN409 : _GEN408;
wire  _GEN411 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN412 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN413 = io_x[1] ? _GEN412 : _GEN411;
wire  _GEN414 = io_x[9] ? _GEN413 : _GEN410;
wire  _GEN415 = io_x[13] ? _GEN414 : _GEN407;
wire  _GEN416 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN417 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN418 = io_x[1] ? _GEN417 : _GEN416;
wire  _GEN419 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN420 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN421 = io_x[1] ? _GEN420 : _GEN419;
wire  _GEN422 = io_x[9] ? _GEN421 : _GEN418;
wire  _GEN423 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN424 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN425 = io_x[1] ? _GEN424 : _GEN423;
wire  _GEN426 = io_x[5] ? _GEN368 : _GEN369;
wire  _GEN427 = io_x[5] ? _GEN369 : _GEN368;
wire  _GEN428 = io_x[1] ? _GEN427 : _GEN426;
wire  _GEN429 = io_x[9] ? _GEN428 : _GEN425;
wire  _GEN430 = io_x[13] ? _GEN429 : _GEN422;
wire  _GEN431 = io_x[0] ? _GEN430 : _GEN415;
wire  _GEN432 = io_x[43] ? _GEN431 : _GEN400;
assign io_y[7] = _GEN432;
wire  _GEN433 = 1'b0;
wire  _GEN434 = 1'b1;
wire  _GEN435 = io_x[8] ? _GEN434 : _GEN433;
wire  _GEN436 = io_x[8] ? _GEN433 : _GEN434;
wire  _GEN437 = io_x[12] ? _GEN436 : _GEN435;
wire  _GEN438 = io_x[8] ? _GEN433 : _GEN434;
wire  _GEN439 = io_x[8] ? _GEN434 : _GEN433;
wire  _GEN440 = io_x[12] ? _GEN439 : _GEN438;
wire  _GEN441 = io_x[4] ? _GEN440 : _GEN437;
wire  _GEN442 = io_x[8] ? _GEN433 : _GEN434;
wire  _GEN443 = io_x[8] ? _GEN434 : _GEN433;
wire  _GEN444 = io_x[12] ? _GEN443 : _GEN442;
wire  _GEN445 = io_x[8] ? _GEN434 : _GEN433;
wire  _GEN446 = io_x[8] ? _GEN433 : _GEN434;
wire  _GEN447 = io_x[12] ? _GEN446 : _GEN445;
wire  _GEN448 = io_x[4] ? _GEN447 : _GEN444;
wire  _GEN449 = io_x[0] ? _GEN448 : _GEN441;
wire  _GEN450 = io_x[8] ? _GEN433 : _GEN434;
wire  _GEN451 = io_x[8] ? _GEN434 : _GEN433;
wire  _GEN452 = io_x[12] ? _GEN451 : _GEN450;
wire  _GEN453 = io_x[8] ? _GEN434 : _GEN433;
wire  _GEN454 = io_x[8] ? _GEN433 : _GEN434;
wire  _GEN455 = io_x[12] ? _GEN454 : _GEN453;
wire  _GEN456 = io_x[4] ? _GEN455 : _GEN452;
wire  _GEN457 = io_x[8] ? _GEN434 : _GEN433;
wire  _GEN458 = io_x[8] ? _GEN433 : _GEN434;
wire  _GEN459 = io_x[12] ? _GEN458 : _GEN457;
wire  _GEN460 = io_x[8] ? _GEN433 : _GEN434;
wire  _GEN461 = io_x[8] ? _GEN434 : _GEN433;
wire  _GEN462 = io_x[12] ? _GEN461 : _GEN460;
wire  _GEN463 = io_x[4] ? _GEN462 : _GEN459;
wire  _GEN464 = io_x[0] ? _GEN463 : _GEN456;
wire  _GEN465 = io_x[42] ? _GEN464 : _GEN449;
assign io_y[6] = _GEN465;
wire  _GEN466 = 1'b0;
wire  _GEN467 = 1'b1;
wire  _GEN468 = io_x[41] ? _GEN467 : _GEN466;
assign io_y[5] = _GEN468;
wire  _GEN469 = 1'b0;
wire  _GEN470 = 1'b1;
wire  _GEN471 = io_x[40] ? _GEN470 : _GEN469;
assign io_y[4] = _GEN471;
wire  _GEN472 = 1'b0;
wire  _GEN473 = 1'b1;
wire  _GEN474 = io_x[39] ? _GEN473 : _GEN472;
assign io_y[3] = _GEN474;
wire  _GEN475 = 1'b0;
wire  _GEN476 = 1'b1;
wire  _GEN477 = io_x[38] ? _GEN476 : _GEN475;
assign io_y[2] = _GEN477;
wire  _GEN478 = 1'b0;
wire  _GEN479 = 1'b1;
wire  _GEN480 = io_x[37] ? _GEN479 : _GEN478;
assign io_y[1] = _GEN480;
wire  _GEN481 = 1'b0;
wire  _GEN482 = 1'b1;
wire  _GEN483 = io_x[34] ? _GEN482 : _GEN481;
assign io_y[0] = _GEN483;
endmodule
