module BBGSharePredictorImp_BSD_NutShell(
    input [31:0] pc,
    input [31:0] train_pc,
    input  train_taken,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    input [15:0] train_ghr_rdata,
    output  taken,
    output  pht_wdata,
    output [8:0] pht_raddr,
    output [8:0] pht_waddr,
    output  ghr_wdata
);
wire [98:0] io_x;
wire [20:0] io_y;
assign io_x = { pc, train_pc, train_taken, pht_rdata, ghr_rdata, train_ghr_rdata };
assign { taken, pht_wdata, pht_raddr, pht_waddr, ghr_wdata } = io_y;
wire  _GEN0 = 1'b1;
wire  _GEN1 = 1'b1;
wire  _GEN2 = 1'b1;
wire  _GEN3 = 1'b0;
wire  _GEN4 = io_x[15] ? _GEN3 : _GEN2;
wire  _GEN5 = 1'b1;
wire  _GEN6 = io_x[42] ? _GEN5 : _GEN4;
wire  _GEN7 = io_x[43] ? _GEN6 : _GEN1;
wire  _GEN8 = 1'b1;
wire  _GEN9 = io_x[38] ? _GEN8 : _GEN7;
wire  _GEN10 = 1'b0;
wire  _GEN11 = 1'b1;
wire  _GEN12 = io_x[2] ? _GEN11 : _GEN10;
wire  _GEN13 = io_x[15] ? _GEN12 : _GEN2;
wire  _GEN14 = io_x[42] ? _GEN5 : _GEN13;
wire  _GEN15 = io_x[43] ? _GEN14 : _GEN1;
wire  _GEN16 = 1'b1;
wire  _GEN17 = 1'b1;
wire  _GEN18 = 1'b0;
wire  _GEN19 = 1'b0;
wire  _GEN20 = 1'b1;
wire  _GEN21 = io_x[30] ? _GEN20 : _GEN19;
wire  _GEN22 = io_x[69] ? _GEN21 : _GEN18;
wire  _GEN23 = io_x[16] ? _GEN22 : _GEN17;
wire  _GEN24 = io_x[40] ? _GEN23 : _GEN16;
wire  _GEN25 = 1'b0;
wire  _GEN26 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN27 = io_x[40] ? _GEN26 : _GEN16;
wire  _GEN28 = io_x[2] ? _GEN27 : _GEN24;
wire  _GEN29 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN30 = io_x[40] ? _GEN29 : _GEN16;
wire  _GEN31 = 1'b0;
wire  _GEN32 = 1'b0;
wire  _GEN33 = 1'b0;
wire  _GEN34 = 1'b1;
wire  _GEN35 = 1'b0;
wire  _GEN36 = io_x[19] ? _GEN35 : _GEN34;
wire  _GEN37 = 1'b1;
wire  _GEN38 = io_x[70] ? _GEN37 : _GEN36;
wire  _GEN39 = io_x[7] ? _GEN38 : _GEN33;
wire  _GEN40 = io_x[18] ? _GEN39 : _GEN32;
wire  _GEN41 = io_x[4] ? _GEN40 : _GEN31;
wire  _GEN42 = io_x[30] ? _GEN41 : _GEN19;
wire  _GEN43 = io_x[69] ? _GEN42 : _GEN18;
wire  _GEN44 = io_x[16] ? _GEN43 : _GEN17;
wire  _GEN45 = io_x[40] ? _GEN44 : _GEN16;
wire  _GEN46 = io_x[2] ? _GEN45 : _GEN30;
wire  _GEN47 = io_x[15] ? _GEN46 : _GEN28;
wire  _GEN48 = io_x[42] ? _GEN47 : _GEN5;
wire  _GEN49 = io_x[43] ? _GEN1 : _GEN48;
wire  _GEN50 = io_x[38] ? _GEN49 : _GEN15;
wire  _GEN51 = io_x[17] ? _GEN50 : _GEN9;
wire  _GEN52 = 1'b1;
wire  _GEN53 = io_x[30] ? _GEN20 : _GEN19;
wire  _GEN54 = io_x[69] ? _GEN53 : _GEN52;
wire  _GEN55 = io_x[16] ? _GEN17 : _GEN54;
wire  _GEN56 = io_x[40] ? _GEN55 : _GEN16;
wire  _GEN57 = io_x[2] ? _GEN11 : _GEN56;
wire  _GEN58 = io_x[15] ? _GEN2 : _GEN57;
wire  _GEN59 = io_x[42] ? _GEN5 : _GEN58;
wire  _GEN60 = io_x[43] ? _GEN1 : _GEN59;
wire  _GEN61 = io_x[38] ? _GEN60 : _GEN8;
wire  _GEN62 = io_x[69] ? _GEN18 : _GEN52;
wire  _GEN63 = io_x[16] ? _GEN17 : _GEN62;
wire  _GEN64 = io_x[40] ? _GEN16 : _GEN63;
wire  _GEN65 = io_x[2] ? _GEN11 : _GEN64;
wire  _GEN66 = io_x[15] ? _GEN65 : _GEN2;
wire  _GEN67 = io_x[42] ? _GEN5 : _GEN66;
wire  _GEN68 = io_x[43] ? _GEN1 : _GEN67;
wire  _GEN69 = io_x[16] ? _GEN17 : _GEN25;
wire  _GEN70 = io_x[40] ? _GEN69 : _GEN16;
wire  _GEN71 = io_x[69] ? _GEN18 : _GEN52;
wire  _GEN72 = io_x[16] ? _GEN71 : _GEN25;
wire  _GEN73 = io_x[40] ? _GEN72 : _GEN16;
wire  _GEN74 = io_x[2] ? _GEN73 : _GEN70;
wire  _GEN75 = io_x[30] ? _GEN20 : _GEN19;
wire  _GEN76 = io_x[69] ? _GEN75 : _GEN52;
wire  _GEN77 = io_x[16] ? _GEN76 : _GEN25;
wire  _GEN78 = io_x[40] ? _GEN77 : _GEN16;
wire  _GEN79 = 1'b1;
wire  _GEN80 = io_x[4] ? _GEN79 : _GEN31;
wire  _GEN81 = io_x[30] ? _GEN80 : _GEN20;
wire  _GEN82 = io_x[69] ? _GEN81 : _GEN52;
wire  _GEN83 = io_x[69] ? _GEN18 : _GEN52;
wire  _GEN84 = io_x[16] ? _GEN83 : _GEN82;
wire  _GEN85 = io_x[40] ? _GEN84 : _GEN16;
wire  _GEN86 = io_x[2] ? _GEN85 : _GEN78;
wire  _GEN87 = io_x[15] ? _GEN86 : _GEN74;
wire  _GEN88 = io_x[42] ? _GEN5 : _GEN87;
wire  _GEN89 = io_x[43] ? _GEN1 : _GEN88;
wire  _GEN90 = io_x[38] ? _GEN89 : _GEN68;
wire  _GEN91 = io_x[17] ? _GEN90 : _GEN61;
wire  _GEN92 = io_x[39] ? _GEN91 : _GEN51;
wire  _GEN93 = 1'b1;
wire  _GEN94 = 1'b1;
wire  _GEN95 = 1'b0;
wire  _GEN96 = io_x[70] ? _GEN95 : _GEN37;
wire  _GEN97 = 1'b1;
wire  _GEN98 = io_x[7] ? _GEN97 : _GEN96;
wire  _GEN99 = io_x[18] ? _GEN98 : _GEN94;
wire  _GEN100 = io_x[4] ? _GEN99 : _GEN79;
wire  _GEN101 = io_x[30] ? _GEN20 : _GEN100;
wire  _GEN102 = io_x[69] ? _GEN52 : _GEN101;
wire  _GEN103 = io_x[16] ? _GEN102 : _GEN17;
wire  _GEN104 = io_x[40] ? _GEN103 : _GEN16;
wire  _GEN105 = io_x[2] ? _GEN104 : _GEN11;
wire  _GEN106 = io_x[15] ? _GEN2 : _GEN105;
wire  _GEN107 = io_x[42] ? _GEN106 : _GEN5;
wire  _GEN108 = io_x[43] ? _GEN1 : _GEN107;
wire  _GEN109 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN110 = io_x[40] ? _GEN16 : _GEN109;
wire  _GEN111 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN112 = io_x[40] ? _GEN16 : _GEN111;
wire  _GEN113 = io_x[2] ? _GEN112 : _GEN110;
wire  _GEN114 = io_x[18] ? _GEN32 : _GEN94;
wire  _GEN115 = io_x[4] ? _GEN114 : _GEN79;
wire  _GEN116 = io_x[30] ? _GEN115 : _GEN20;
wire  _GEN117 = io_x[69] ? _GEN18 : _GEN116;
wire  _GEN118 = io_x[16] ? _GEN117 : _GEN17;
wire  _GEN119 = io_x[40] ? _GEN16 : _GEN118;
wire  _GEN120 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN121 = io_x[40] ? _GEN16 : _GEN120;
wire  _GEN122 = io_x[2] ? _GEN121 : _GEN119;
wire  _GEN123 = io_x[15] ? _GEN122 : _GEN113;
wire  _GEN124 = io_x[42] ? _GEN123 : _GEN5;
wire  _GEN125 = io_x[43] ? _GEN1 : _GEN124;
wire  _GEN126 = io_x[38] ? _GEN125 : _GEN108;
wire  _GEN127 = io_x[17] ? _GEN126 : _GEN93;
wire  _GEN128 = io_x[4] ? _GEN79 : _GEN31;
wire  _GEN129 = io_x[30] ? _GEN19 : _GEN128;
wire  _GEN130 = io_x[69] ? _GEN52 : _GEN129;
wire  _GEN131 = io_x[16] ? _GEN130 : _GEN17;
wire  _GEN132 = io_x[40] ? _GEN16 : _GEN131;
wire  _GEN133 = io_x[19] ? _GEN35 : _GEN34;
wire  _GEN134 = io_x[70] ? _GEN37 : _GEN133;
wire  _GEN135 = io_x[7] ? _GEN97 : _GEN134;
wire  _GEN136 = io_x[18] ? _GEN135 : _GEN94;
wire  _GEN137 = io_x[4] ? _GEN79 : _GEN136;
wire  _GEN138 = io_x[30] ? _GEN20 : _GEN137;
wire  _GEN139 = io_x[69] ? _GEN52 : _GEN138;
wire  _GEN140 = io_x[16] ? _GEN139 : _GEN17;
wire  _GEN141 = io_x[40] ? _GEN16 : _GEN140;
wire  _GEN142 = io_x[2] ? _GEN141 : _GEN132;
wire  _GEN143 = io_x[30] ? _GEN20 : _GEN19;
wire  _GEN144 = io_x[69] ? _GEN52 : _GEN143;
wire  _GEN145 = io_x[16] ? _GEN144 : _GEN17;
wire  _GEN146 = io_x[40] ? _GEN16 : _GEN145;
wire  _GEN147 = io_x[2] ? _GEN11 : _GEN146;
wire  _GEN148 = io_x[15] ? _GEN147 : _GEN142;
wire  _GEN149 = io_x[42] ? _GEN148 : _GEN5;
wire  _GEN150 = io_x[43] ? _GEN1 : _GEN149;
wire  _GEN151 = io_x[38] ? _GEN8 : _GEN150;
wire  _GEN152 = io_x[4] ? _GEN79 : _GEN31;
wire  _GEN153 = io_x[30] ? _GEN152 : _GEN20;
wire  _GEN154 = io_x[69] ? _GEN52 : _GEN153;
wire  _GEN155 = io_x[18] ? _GEN94 : _GEN32;
wire  _GEN156 = io_x[4] ? _GEN155 : _GEN79;
wire  _GEN157 = io_x[30] ? _GEN156 : _GEN20;
wire  _GEN158 = io_x[69] ? _GEN52 : _GEN157;
wire  _GEN159 = io_x[16] ? _GEN158 : _GEN154;
wire  _GEN160 = io_x[40] ? _GEN16 : _GEN159;
wire  _GEN161 = io_x[2] ? _GEN11 : _GEN160;
wire  _GEN162 = io_x[7] ? _GEN33 : _GEN97;
wire  _GEN163 = io_x[18] ? _GEN162 : _GEN94;
wire  _GEN164 = io_x[4] ? _GEN163 : _GEN79;
wire  _GEN165 = io_x[30] ? _GEN164 : _GEN20;
wire  _GEN166 = io_x[69] ? _GEN52 : _GEN165;
wire  _GEN167 = io_x[16] ? _GEN166 : _GEN17;
wire  _GEN168 = io_x[40] ? _GEN16 : _GEN167;
wire  _GEN169 = io_x[2] ? _GEN168 : _GEN11;
wire  _GEN170 = io_x[15] ? _GEN169 : _GEN161;
wire  _GEN171 = io_x[42] ? _GEN170 : _GEN5;
wire  _GEN172 = io_x[43] ? _GEN1 : _GEN171;
wire  _GEN173 = io_x[38] ? _GEN8 : _GEN172;
wire  _GEN174 = io_x[17] ? _GEN173 : _GEN151;
wire  _GEN175 = io_x[39] ? _GEN174 : _GEN127;
wire  _GEN176 = io_x[37] ? _GEN175 : _GEN92;
wire  _GEN177 = 1'b1;
wire  _GEN178 = 1'b0;
wire  _GEN179 = io_x[43] ? _GEN178 : _GEN1;
wire  _GEN180 = io_x[38] ? _GEN8 : _GEN179;
wire  _GEN181 = 1'b0;
wire  _GEN182 = io_x[40] ? _GEN16 : _GEN181;
wire  _GEN183 = io_x[2] ? _GEN182 : _GEN11;
wire  _GEN184 = io_x[40] ? _GEN16 : _GEN181;
wire  _GEN185 = io_x[2] ? _GEN184 : _GEN10;
wire  _GEN186 = io_x[15] ? _GEN185 : _GEN183;
wire  _GEN187 = io_x[42] ? _GEN5 : _GEN186;
wire  _GEN188 = io_x[43] ? _GEN187 : _GEN1;
wire  _GEN189 = io_x[2] ? _GEN10 : _GEN11;
wire  _GEN190 = io_x[40] ? _GEN16 : _GEN181;
wire  _GEN191 = io_x[2] ? _GEN190 : _GEN11;
wire  _GEN192 = io_x[15] ? _GEN191 : _GEN189;
wire  _GEN193 = io_x[42] ? _GEN5 : _GEN192;
wire  _GEN194 = io_x[43] ? _GEN1 : _GEN193;
wire  _GEN195 = io_x[38] ? _GEN194 : _GEN188;
wire  _GEN196 = io_x[17] ? _GEN195 : _GEN180;
wire  _GEN197 = io_x[39] ? _GEN196 : _GEN177;
wire  _GEN198 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN199 = io_x[2] ? _GEN198 : _GEN11;
wire  _GEN200 = io_x[15] ? _GEN3 : _GEN199;
wire  _GEN201 = io_x[42] ? _GEN200 : _GEN5;
wire  _GEN202 = io_x[70] ? _GEN95 : _GEN37;
wire  _GEN203 = io_x[7] ? _GEN202 : _GEN97;
wire  _GEN204 = io_x[18] ? _GEN203 : _GEN94;
wire  _GEN205 = io_x[4] ? _GEN204 : _GEN79;
wire  _GEN206 = 1'b1;
wire  _GEN207 = 1'b1;
wire  _GEN208 = 1'b1;
wire  _GEN209 = 1'b0;
wire  _GEN210 = io_x[74] ? _GEN209 : _GEN208;
wire  _GEN211 = io_x[76] ? _GEN210 : _GEN207;
wire  _GEN212 = io_x[31] ? _GEN211 : _GEN206;
wire  _GEN213 = io_x[19] ? _GEN212 : _GEN34;
wire  _GEN214 = io_x[70] ? _GEN95 : _GEN213;
wire  _GEN215 = io_x[7] ? _GEN214 : _GEN33;
wire  _GEN216 = io_x[18] ? _GEN215 : _GEN94;
wire  _GEN217 = io_x[4] ? _GEN216 : _GEN31;
wire  _GEN218 = io_x[30] ? _GEN217 : _GEN205;
wire  _GEN219 = io_x[69] ? _GEN218 : _GEN18;
wire  _GEN220 = io_x[16] ? _GEN219 : _GEN17;
wire  _GEN221 = io_x[40] ? _GEN16 : _GEN220;
wire  _GEN222 = io_x[2] ? _GEN221 : _GEN10;
wire  _GEN223 = io_x[15] ? _GEN222 : _GEN2;
wire  _GEN224 = io_x[42] ? _GEN5 : _GEN223;
wire  _GEN225 = io_x[43] ? _GEN224 : _GEN201;
wire  _GEN226 = io_x[38] ? _GEN225 : _GEN8;
wire  _GEN227 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN228 = io_x[2] ? _GEN10 : _GEN227;
wire  _GEN229 = io_x[15] ? _GEN3 : _GEN228;
wire  _GEN230 = io_x[42] ? _GEN229 : _GEN5;
wire  _GEN231 = io_x[4] ? _GEN31 : _GEN79;
wire  _GEN232 = io_x[30] ? _GEN20 : _GEN231;
wire  _GEN233 = io_x[69] ? _GEN52 : _GEN232;
wire  _GEN234 = io_x[16] ? _GEN233 : _GEN17;
wire  _GEN235 = io_x[40] ? _GEN16 : _GEN234;
wire  _GEN236 = 1'b0;
wire  _GEN237 = io_x[31] ? _GEN236 : _GEN206;
wire  _GEN238 = io_x[19] ? _GEN237 : _GEN34;
wire  _GEN239 = io_x[70] ? _GEN238 : _GEN37;
wire  _GEN240 = io_x[7] ? _GEN239 : _GEN33;
wire  _GEN241 = io_x[18] ? _GEN240 : _GEN32;
wire  _GEN242 = io_x[4] ? _GEN241 : _GEN79;
wire  _GEN243 = io_x[30] ? _GEN242 : _GEN19;
wire  _GEN244 = io_x[69] ? _GEN243 : _GEN18;
wire  _GEN245 = io_x[16] ? _GEN244 : _GEN17;
wire  _GEN246 = io_x[40] ? _GEN16 : _GEN245;
wire  _GEN247 = io_x[2] ? _GEN246 : _GEN235;
wire  _GEN248 = 1'b0;
wire  _GEN249 = io_x[76] ? _GEN248 : _GEN207;
wire  _GEN250 = io_x[31] ? _GEN249 : _GEN236;
wire  _GEN251 = io_x[19] ? _GEN250 : _GEN34;
wire  _GEN252 = io_x[70] ? _GEN95 : _GEN251;
wire  _GEN253 = io_x[7] ? _GEN252 : _GEN33;
wire  _GEN254 = io_x[18] ? _GEN253 : _GEN32;
wire  _GEN255 = io_x[4] ? _GEN254 : _GEN31;
wire  _GEN256 = io_x[30] ? _GEN255 : _GEN19;
wire  _GEN257 = io_x[76] ? _GEN248 : _GEN207;
wire  _GEN258 = io_x[31] ? _GEN257 : _GEN206;
wire  _GEN259 = io_x[19] ? _GEN258 : _GEN34;
wire  _GEN260 = io_x[70] ? _GEN37 : _GEN259;
wire  _GEN261 = io_x[7] ? _GEN33 : _GEN260;
wire  _GEN262 = io_x[76] ? _GEN248 : _GEN207;
wire  _GEN263 = io_x[31] ? _GEN262 : _GEN236;
wire  _GEN264 = io_x[19] ? _GEN263 : _GEN34;
wire  _GEN265 = io_x[70] ? _GEN95 : _GEN264;
wire  _GEN266 = io_x[7] ? _GEN265 : _GEN33;
wire  _GEN267 = io_x[18] ? _GEN266 : _GEN261;
wire  _GEN268 = io_x[4] ? _GEN267 : _GEN31;
wire  _GEN269 = io_x[30] ? _GEN268 : _GEN19;
wire  _GEN270 = io_x[69] ? _GEN269 : _GEN256;
wire  _GEN271 = io_x[16] ? _GEN270 : _GEN17;
wire  _GEN272 = io_x[40] ? _GEN16 : _GEN271;
wire  _GEN273 = io_x[2] ? _GEN272 : _GEN10;
wire  _GEN274 = io_x[15] ? _GEN273 : _GEN247;
wire  _GEN275 = io_x[42] ? _GEN5 : _GEN274;
wire  _GEN276 = io_x[43] ? _GEN275 : _GEN230;
wire  _GEN277 = io_x[38] ? _GEN276 : _GEN8;
wire  _GEN278 = io_x[17] ? _GEN277 : _GEN226;
wire  _GEN279 = io_x[39] ? _GEN177 : _GEN278;
wire  _GEN280 = io_x[37] ? _GEN279 : _GEN197;
wire  _GEN281 = io_x[77] ? _GEN280 : _GEN176;
wire  _GEN282 = 1'b1;
wire  _GEN283 = io_x[7] ? _GEN33 : _GEN97;
wire  _GEN284 = io_x[18] ? _GEN283 : _GEN94;
wire  _GEN285 = io_x[31] ? _GEN236 : _GEN206;
wire  _GEN286 = io_x[19] ? _GEN285 : _GEN34;
wire  _GEN287 = io_x[70] ? _GEN37 : _GEN286;
wire  _GEN288 = io_x[7] ? _GEN287 : _GEN97;
wire  _GEN289 = io_x[18] ? _GEN288 : _GEN94;
wire  _GEN290 = io_x[4] ? _GEN289 : _GEN284;
wire  _GEN291 = io_x[31] ? _GEN236 : _GEN206;
wire  _GEN292 = io_x[19] ? _GEN291 : _GEN34;
wire  _GEN293 = io_x[70] ? _GEN37 : _GEN292;
wire  _GEN294 = io_x[7] ? _GEN293 : _GEN97;
wire  _GEN295 = io_x[18] ? _GEN294 : _GEN94;
wire  _GEN296 = io_x[4] ? _GEN295 : _GEN79;
wire  _GEN297 = io_x[30] ? _GEN296 : _GEN290;
wire  _GEN298 = io_x[69] ? _GEN297 : _GEN52;
wire  _GEN299 = io_x[16] ? _GEN298 : _GEN17;
wire  _GEN300 = io_x[40] ? _GEN16 : _GEN299;
wire  _GEN301 = io_x[2] ? _GEN300 : _GEN11;
wire  _GEN302 = io_x[18] ? _GEN32 : _GEN94;
wire  _GEN303 = io_x[4] ? _GEN302 : _GEN79;
wire  _GEN304 = io_x[19] ? _GEN35 : _GEN34;
wire  _GEN305 = io_x[70] ? _GEN37 : _GEN304;
wire  _GEN306 = io_x[7] ? _GEN305 : _GEN33;
wire  _GEN307 = io_x[18] ? _GEN306 : _GEN94;
wire  _GEN308 = 1'b0;
wire  _GEN309 = 1'b1;
wire  _GEN310 = io_x[21] ? _GEN309 : _GEN308;
wire  _GEN311 = io_x[74] ? _GEN208 : _GEN310;
wire  _GEN312 = io_x[76] ? _GEN207 : _GEN311;
wire  _GEN313 = io_x[31] ? _GEN312 : _GEN236;
wire  _GEN314 = io_x[19] ? _GEN313 : _GEN34;
wire  _GEN315 = io_x[70] ? _GEN37 : _GEN314;
wire  _GEN316 = io_x[7] ? _GEN315 : _GEN97;
wire  _GEN317 = io_x[18] ? _GEN316 : _GEN94;
wire  _GEN318 = io_x[4] ? _GEN317 : _GEN307;
wire  _GEN319 = io_x[30] ? _GEN318 : _GEN303;
wire  _GEN320 = io_x[69] ? _GEN319 : _GEN52;
wire  _GEN321 = io_x[16] ? _GEN320 : _GEN17;
wire  _GEN322 = io_x[40] ? _GEN16 : _GEN321;
wire  _GEN323 = io_x[2] ? _GEN322 : _GEN11;
wire  _GEN324 = io_x[15] ? _GEN323 : _GEN301;
wire  _GEN325 = io_x[42] ? _GEN5 : _GEN324;
wire  _GEN326 = io_x[43] ? _GEN325 : _GEN1;
wire  _GEN327 = io_x[31] ? _GEN206 : _GEN236;
wire  _GEN328 = io_x[19] ? _GEN327 : _GEN34;
wire  _GEN329 = io_x[70] ? _GEN37 : _GEN328;
wire  _GEN330 = io_x[7] ? _GEN97 : _GEN329;
wire  _GEN331 = io_x[18] ? _GEN330 : _GEN94;
wire  _GEN332 = io_x[4] ? _GEN79 : _GEN331;
wire  _GEN333 = io_x[30] ? _GEN332 : _GEN20;
wire  _GEN334 = io_x[69] ? _GEN333 : _GEN52;
wire  _GEN335 = io_x[16] ? _GEN334 : _GEN17;
wire  _GEN336 = io_x[40] ? _GEN335 : _GEN16;
wire  _GEN337 = io_x[2] ? _GEN11 : _GEN336;
wire  _GEN338 = io_x[15] ? _GEN2 : _GEN337;
wire  _GEN339 = io_x[42] ? _GEN338 : _GEN5;
wire  _GEN340 = io_x[43] ? _GEN1 : _GEN339;
wire  _GEN341 = io_x[38] ? _GEN340 : _GEN326;
wire  _GEN342 = io_x[17] ? _GEN341 : _GEN93;
wire  _GEN343 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN344 = io_x[2] ? _GEN343 : _GEN11;
wire  _GEN345 = io_x[15] ? _GEN344 : _GEN2;
wire  _GEN346 = io_x[42] ? _GEN5 : _GEN345;
wire  _GEN347 = io_x[43] ? _GEN1 : _GEN346;
wire  _GEN348 = io_x[38] ? _GEN8 : _GEN347;
wire  _GEN349 = io_x[17] ? _GEN348 : _GEN93;
wire  _GEN350 = io_x[39] ? _GEN349 : _GEN342;
wire  _GEN351 = 1'b1;
wire  _GEN352 = io_x[37] ? _GEN351 : _GEN350;
wire  _GEN353 = io_x[77] ? _GEN352 : _GEN282;
wire  _GEN354 = io_x[78] ? _GEN353 : _GEN281;
wire  _GEN355 = io_x[70] ? _GEN95 : _GEN37;
wire  _GEN356 = io_x[7] ? _GEN355 : _GEN97;
wire  _GEN357 = io_x[18] ? _GEN356 : _GEN94;
wire  _GEN358 = io_x[4] ? _GEN357 : _GEN79;
wire  _GEN359 = io_x[30] ? _GEN20 : _GEN358;
wire  _GEN360 = io_x[69] ? _GEN52 : _GEN359;
wire  _GEN361 = io_x[16] ? _GEN360 : _GEN17;
wire  _GEN362 = io_x[40] ? _GEN16 : _GEN361;
wire  _GEN363 = io_x[2] ? _GEN362 : _GEN11;
wire  _GEN364 = io_x[70] ? _GEN95 : _GEN37;
wire  _GEN365 = io_x[7] ? _GEN97 : _GEN364;
wire  _GEN366 = io_x[18] ? _GEN365 : _GEN94;
wire  _GEN367 = io_x[4] ? _GEN79 : _GEN366;
wire  _GEN368 = io_x[30] ? _GEN367 : _GEN20;
wire  _GEN369 = io_x[69] ? _GEN52 : _GEN368;
wire  _GEN370 = io_x[16] ? _GEN369 : _GEN17;
wire  _GEN371 = io_x[40] ? _GEN16 : _GEN370;
wire  _GEN372 = io_x[2] ? _GEN371 : _GEN11;
wire  _GEN373 = io_x[15] ? _GEN372 : _GEN363;
wire  _GEN374 = io_x[42] ? _GEN373 : _GEN5;
wire  _GEN375 = io_x[43] ? _GEN1 : _GEN374;
wire  _GEN376 = io_x[38] ? _GEN8 : _GEN375;
wire  _GEN377 = io_x[69] ? _GEN52 : _GEN18;
wire  _GEN378 = io_x[16] ? _GEN377 : _GEN17;
wire  _GEN379 = io_x[40] ? _GEN16 : _GEN378;
wire  _GEN380 = io_x[2] ? _GEN379 : _GEN11;
wire  _GEN381 = io_x[40] ? _GEN16 : _GEN181;
wire  _GEN382 = io_x[2] ? _GEN11 : _GEN381;
wire  _GEN383 = io_x[15] ? _GEN382 : _GEN380;
wire  _GEN384 = io_x[42] ? _GEN383 : _GEN5;
wire  _GEN385 = io_x[43] ? _GEN1 : _GEN384;
wire  _GEN386 = io_x[38] ? _GEN8 : _GEN385;
wire  _GEN387 = io_x[17] ? _GEN386 : _GEN376;
wire  _GEN388 = io_x[7] ? _GEN97 : _GEN33;
wire  _GEN389 = io_x[18] ? _GEN388 : _GEN94;
wire  _GEN390 = io_x[4] ? _GEN79 : _GEN389;
wire  _GEN391 = io_x[30] ? _GEN390 : _GEN20;
wire  _GEN392 = io_x[69] ? _GEN391 : _GEN52;
wire  _GEN393 = io_x[16] ? _GEN392 : _GEN17;
wire  _GEN394 = io_x[40] ? _GEN16 : _GEN393;
wire  _GEN395 = io_x[2] ? _GEN394 : _GEN11;
wire  _GEN396 = io_x[15] ? _GEN395 : _GEN2;
wire  _GEN397 = io_x[42] ? _GEN5 : _GEN396;
wire  _GEN398 = io_x[43] ? _GEN1 : _GEN397;
wire  _GEN399 = io_x[38] ? _GEN398 : _GEN8;
wire  _GEN400 = io_x[17] ? _GEN93 : _GEN399;
wire  _GEN401 = io_x[39] ? _GEN400 : _GEN387;
wire  _GEN402 = io_x[43] ? _GEN1 : _GEN178;
wire  _GEN403 = io_x[38] ? _GEN8 : _GEN402;
wire  _GEN404 = io_x[4] ? _GEN31 : _GEN79;
wire  _GEN405 = io_x[30] ? _GEN20 : _GEN404;
wire  _GEN406 = io_x[69] ? _GEN52 : _GEN405;
wire  _GEN407 = io_x[16] ? _GEN17 : _GEN406;
wire  _GEN408 = io_x[40] ? _GEN407 : _GEN16;
wire  _GEN409 = io_x[18] ? _GEN32 : _GEN94;
wire  _GEN410 = io_x[4] ? _GEN409 : _GEN79;
wire  _GEN411 = io_x[30] ? _GEN20 : _GEN410;
wire  _GEN412 = io_x[69] ? _GEN52 : _GEN411;
wire  _GEN413 = io_x[16] ? _GEN17 : _GEN412;
wire  _GEN414 = io_x[40] ? _GEN413 : _GEN16;
wire  _GEN415 = io_x[2] ? _GEN414 : _GEN408;
wire  _GEN416 = io_x[70] ? _GEN95 : _GEN37;
wire  _GEN417 = io_x[7] ? _GEN97 : _GEN416;
wire  _GEN418 = io_x[18] ? _GEN94 : _GEN417;
wire  _GEN419 = io_x[4] ? _GEN79 : _GEN418;
wire  _GEN420 = io_x[30] ? _GEN419 : _GEN20;
wire  _GEN421 = io_x[69] ? _GEN52 : _GEN420;
wire  _GEN422 = io_x[16] ? _GEN17 : _GEN421;
wire  _GEN423 = io_x[40] ? _GEN422 : _GEN16;
wire  _GEN424 = io_x[2] ? _GEN11 : _GEN423;
wire  _GEN425 = io_x[15] ? _GEN424 : _GEN415;
wire  _GEN426 = io_x[42] ? _GEN5 : _GEN425;
wire  _GEN427 = io_x[43] ? _GEN1 : _GEN426;
wire  _GEN428 = io_x[38] ? _GEN8 : _GEN427;
wire  _GEN429 = io_x[17] ? _GEN428 : _GEN403;
wire  _GEN430 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN431 = io_x[2] ? _GEN430 : _GEN10;
wire  _GEN432 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN433 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN434 = io_x[2] ? _GEN433 : _GEN432;
wire  _GEN435 = io_x[15] ? _GEN434 : _GEN431;
wire  _GEN436 = io_x[42] ? _GEN5 : _GEN435;
wire  _GEN437 = io_x[43] ? _GEN1 : _GEN436;
wire  _GEN438 = io_x[38] ? _GEN437 : _GEN8;
wire  _GEN439 = io_x[17] ? _GEN438 : _GEN93;
wire  _GEN440 = io_x[39] ? _GEN439 : _GEN429;
wire  _GEN441 = io_x[37] ? _GEN440 : _GEN401;
wire  _GEN442 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN443 = io_x[2] ? _GEN10 : _GEN442;
wire  _GEN444 = io_x[2] ? _GEN10 : _GEN11;
wire  _GEN445 = io_x[15] ? _GEN444 : _GEN443;
wire  _GEN446 = io_x[42] ? _GEN5 : _GEN445;
wire  _GEN447 = io_x[43] ? _GEN1 : _GEN446;
wire  _GEN448 = io_x[38] ? _GEN447 : _GEN8;
wire  _GEN449 = io_x[69] ? _GEN52 : _GEN18;
wire  _GEN450 = io_x[16] ? _GEN449 : _GEN17;
wire  _GEN451 = io_x[16] ? _GEN17 : _GEN25;
wire  _GEN452 = io_x[40] ? _GEN451 : _GEN450;
wire  _GEN453 = io_x[2] ? _GEN10 : _GEN452;
wire  _GEN454 = io_x[15] ? _GEN3 : _GEN453;
wire  _GEN455 = io_x[42] ? _GEN5 : _GEN454;
wire  _GEN456 = io_x[16] ? _GEN17 : _GEN25;
wire  _GEN457 = io_x[40] ? _GEN456 : _GEN16;
wire  _GEN458 = io_x[2] ? _GEN457 : _GEN11;
wire  _GEN459 = io_x[15] ? _GEN3 : _GEN458;
wire  _GEN460 = io_x[42] ? _GEN5 : _GEN459;
wire  _GEN461 = io_x[43] ? _GEN460 : _GEN455;
wire  _GEN462 = io_x[38] ? _GEN461 : _GEN8;
wire  _GEN463 = io_x[17] ? _GEN462 : _GEN448;
wire  _GEN464 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN465 = io_x[40] ? _GEN464 : _GEN16;
wire  _GEN466 = io_x[2] ? _GEN11 : _GEN465;
wire  _GEN467 = io_x[15] ? _GEN466 : _GEN2;
wire  _GEN468 = io_x[42] ? _GEN5 : _GEN467;
wire  _GEN469 = io_x[43] ? _GEN1 : _GEN468;
wire  _GEN470 = io_x[38] ? _GEN8 : _GEN469;
wire  _GEN471 = 1'b0;
wire  _GEN472 = io_x[42] ? _GEN471 : _GEN5;
wire  _GEN473 = io_x[43] ? _GEN1 : _GEN472;
wire  _GEN474 = io_x[38] ? _GEN473 : _GEN8;
wire  _GEN475 = io_x[17] ? _GEN474 : _GEN470;
wire  _GEN476 = io_x[39] ? _GEN475 : _GEN463;
wire  _GEN477 = io_x[4] ? _GEN79 : _GEN31;
wire  _GEN478 = io_x[30] ? _GEN19 : _GEN477;
wire  _GEN479 = io_x[69] ? _GEN52 : _GEN478;
wire  _GEN480 = io_x[16] ? _GEN479 : _GEN17;
wire  _GEN481 = io_x[40] ? _GEN480 : _GEN16;
wire  _GEN482 = io_x[2] ? _GEN11 : _GEN481;
wire  _GEN483 = io_x[4] ? _GEN79 : _GEN31;
wire  _GEN484 = io_x[30] ? _GEN483 : _GEN20;
wire  _GEN485 = io_x[69] ? _GEN52 : _GEN484;
wire  _GEN486 = io_x[16] ? _GEN485 : _GEN17;
wire  _GEN487 = io_x[40] ? _GEN486 : _GEN16;
wire  _GEN488 = io_x[2] ? _GEN487 : _GEN10;
wire  _GEN489 = io_x[15] ? _GEN488 : _GEN482;
wire  _GEN490 = io_x[42] ? _GEN5 : _GEN489;
wire  _GEN491 = io_x[43] ? _GEN1 : _GEN490;
wire  _GEN492 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN493 = io_x[40] ? _GEN492 : _GEN16;
wire  _GEN494 = io_x[2] ? _GEN493 : _GEN11;
wire  _GEN495 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN496 = io_x[40] ? _GEN495 : _GEN16;
wire  _GEN497 = io_x[2] ? _GEN496 : _GEN11;
wire  _GEN498 = io_x[15] ? _GEN497 : _GEN494;
wire  _GEN499 = io_x[42] ? _GEN5 : _GEN498;
wire  _GEN500 = io_x[4] ? _GEN31 : _GEN79;
wire  _GEN501 = io_x[30] ? _GEN500 : _GEN20;
wire  _GEN502 = io_x[69] ? _GEN52 : _GEN501;
wire  _GEN503 = io_x[16] ? _GEN17 : _GEN502;
wire  _GEN504 = io_x[40] ? _GEN16 : _GEN503;
wire  _GEN505 = io_x[2] ? _GEN504 : _GEN11;
wire  _GEN506 = io_x[15] ? _GEN2 : _GEN505;
wire  _GEN507 = io_x[42] ? _GEN506 : _GEN5;
wire  _GEN508 = io_x[43] ? _GEN507 : _GEN499;
wire  _GEN509 = io_x[38] ? _GEN508 : _GEN491;
wire  _GEN510 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN511 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN512 = io_x[2] ? _GEN511 : _GEN510;
wire  _GEN513 = io_x[15] ? _GEN2 : _GEN512;
wire  _GEN514 = io_x[42] ? _GEN5 : _GEN513;
wire  _GEN515 = io_x[43] ? _GEN1 : _GEN514;
wire  _GEN516 = io_x[2] ? _GEN11 : _GEN10;
wire  _GEN517 = io_x[15] ? _GEN2 : _GEN516;
wire  _GEN518 = io_x[42] ? _GEN5 : _GEN517;
wire  _GEN519 = io_x[69] ? _GEN18 : _GEN52;
wire  _GEN520 = io_x[16] ? _GEN17 : _GEN519;
wire  _GEN521 = io_x[40] ? _GEN520 : _GEN16;
wire  _GEN522 = io_x[2] ? _GEN11 : _GEN521;
wire  _GEN523 = io_x[15] ? _GEN2 : _GEN522;
wire  _GEN524 = io_x[42] ? _GEN5 : _GEN523;
wire  _GEN525 = io_x[43] ? _GEN524 : _GEN518;
wire  _GEN526 = io_x[38] ? _GEN525 : _GEN515;
wire  _GEN527 = io_x[17] ? _GEN526 : _GEN509;
wire  _GEN528 = io_x[42] ? _GEN5 : _GEN471;
wire  _GEN529 = io_x[43] ? _GEN528 : _GEN1;
wire  _GEN530 = io_x[30] ? _GEN20 : _GEN19;
wire  _GEN531 = io_x[69] ? _GEN18 : _GEN530;
wire  _GEN532 = io_x[16] ? _GEN531 : _GEN17;
wire  _GEN533 = io_x[40] ? _GEN532 : _GEN16;
wire  _GEN534 = io_x[70] ? _GEN95 : _GEN37;
wire  _GEN535 = io_x[70] ? _GEN95 : _GEN37;
wire  _GEN536 = io_x[7] ? _GEN535 : _GEN534;
wire  _GEN537 = io_x[18] ? _GEN536 : _GEN94;
wire  _GEN538 = io_x[4] ? _GEN537 : _GEN79;
wire  _GEN539 = io_x[30] ? _GEN20 : _GEN538;
wire  _GEN540 = io_x[69] ? _GEN52 : _GEN539;
wire  _GEN541 = io_x[16] ? _GEN540 : _GEN17;
wire  _GEN542 = io_x[40] ? _GEN541 : _GEN16;
wire  _GEN543 = io_x[2] ? _GEN542 : _GEN533;
wire  _GEN544 = io_x[30] ? _GEN20 : _GEN19;
wire  _GEN545 = io_x[4] ? _GEN79 : _GEN31;
wire  _GEN546 = io_x[30] ? _GEN545 : _GEN20;
wire  _GEN547 = io_x[69] ? _GEN546 : _GEN544;
wire  _GEN548 = io_x[16] ? _GEN547 : _GEN17;
wire  _GEN549 = io_x[40] ? _GEN548 : _GEN16;
wire  _GEN550 = io_x[69] ? _GEN18 : _GEN52;
wire  _GEN551 = io_x[16] ? _GEN550 : _GEN17;
wire  _GEN552 = io_x[40] ? _GEN551 : _GEN16;
wire  _GEN553 = io_x[2] ? _GEN552 : _GEN549;
wire  _GEN554 = io_x[15] ? _GEN553 : _GEN543;
wire  _GEN555 = io_x[42] ? _GEN5 : _GEN554;
wire  _GEN556 = io_x[43] ? _GEN1 : _GEN555;
wire  _GEN557 = io_x[38] ? _GEN556 : _GEN529;
wire  _GEN558 = io_x[17] ? _GEN557 : _GEN93;
wire  _GEN559 = io_x[39] ? _GEN558 : _GEN527;
wire  _GEN560 = io_x[37] ? _GEN559 : _GEN476;
wire  _GEN561 = io_x[77] ? _GEN560 : _GEN441;
wire  _GEN562 = io_x[69] ? _GEN18 : _GEN52;
wire  _GEN563 = io_x[16] ? _GEN562 : _GEN17;
wire  _GEN564 = io_x[40] ? _GEN563 : _GEN16;
wire  _GEN565 = io_x[2] ? _GEN11 : _GEN564;
wire  _GEN566 = io_x[15] ? _GEN2 : _GEN565;
wire  _GEN567 = io_x[42] ? _GEN5 : _GEN566;
wire  _GEN568 = io_x[43] ? _GEN567 : _GEN1;
wire  _GEN569 = io_x[76] ? _GEN207 : _GEN248;
wire  _GEN570 = io_x[31] ? _GEN236 : _GEN569;
wire  _GEN571 = io_x[19] ? _GEN570 : _GEN34;
wire  _GEN572 = io_x[70] ? _GEN37 : _GEN571;
wire  _GEN573 = io_x[7] ? _GEN97 : _GEN572;
wire  _GEN574 = io_x[18] ? _GEN573 : _GEN94;
wire  _GEN575 = io_x[4] ? _GEN79 : _GEN574;
wire  _GEN576 = io_x[76] ? _GEN207 : _GEN248;
wire  _GEN577 = io_x[31] ? _GEN576 : _GEN236;
wire  _GEN578 = io_x[19] ? _GEN577 : _GEN35;
wire  _GEN579 = io_x[70] ? _GEN37 : _GEN578;
wire  _GEN580 = io_x[7] ? _GEN97 : _GEN579;
wire  _GEN581 = io_x[18] ? _GEN580 : _GEN94;
wire  _GEN582 = io_x[4] ? _GEN79 : _GEN581;
wire  _GEN583 = io_x[30] ? _GEN582 : _GEN575;
wire  _GEN584 = io_x[69] ? _GEN583 : _GEN52;
wire  _GEN585 = io_x[16] ? _GEN584 : _GEN17;
wire  _GEN586 = io_x[40] ? _GEN16 : _GEN585;
wire  _GEN587 = io_x[2] ? _GEN11 : _GEN586;
wire  _GEN588 = io_x[15] ? _GEN2 : _GEN587;
wire  _GEN589 = io_x[42] ? _GEN588 : _GEN5;
wire  _GEN590 = io_x[43] ? _GEN589 : _GEN1;
wire  _GEN591 = io_x[38] ? _GEN590 : _GEN568;
wire  _GEN592 = io_x[17] ? _GEN591 : _GEN93;
wire  _GEN593 = io_x[2] ? _GEN11 : _GEN10;
wire  _GEN594 = io_x[15] ? _GEN2 : _GEN593;
wire  _GEN595 = io_x[42] ? _GEN594 : _GEN5;
wire  _GEN596 = io_x[43] ? _GEN595 : _GEN1;
wire  _GEN597 = io_x[38] ? _GEN8 : _GEN596;
wire  _GEN598 = io_x[17] ? _GEN597 : _GEN93;
wire  _GEN599 = io_x[39] ? _GEN598 : _GEN592;
wire  _GEN600 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN601 = io_x[40] ? _GEN16 : _GEN600;
wire  _GEN602 = io_x[2] ? _GEN601 : _GEN11;
wire  _GEN603 = io_x[15] ? _GEN602 : _GEN2;
wire  _GEN604 = io_x[2] ? _GEN10 : _GEN11;
wire  _GEN605 = io_x[15] ? _GEN604 : _GEN2;
wire  _GEN606 = io_x[42] ? _GEN605 : _GEN603;
wire  _GEN607 = io_x[43] ? _GEN606 : _GEN1;
wire  _GEN608 = io_x[38] ? _GEN607 : _GEN8;
wire  _GEN609 = io_x[17] ? _GEN608 : _GEN93;
wire  _GEN610 = io_x[4] ? _GEN31 : _GEN79;
wire  _GEN611 = io_x[30] ? _GEN610 : _GEN19;
wire  _GEN612 = io_x[69] ? _GEN611 : _GEN52;
wire  _GEN613 = io_x[16] ? _GEN612 : _GEN17;
wire  _GEN614 = io_x[40] ? _GEN613 : _GEN16;
wire  _GEN615 = io_x[2] ? _GEN11 : _GEN614;
wire  _GEN616 = io_x[15] ? _GEN615 : _GEN2;
wire  _GEN617 = io_x[42] ? _GEN616 : _GEN5;
wire  _GEN618 = io_x[43] ? _GEN617 : _GEN1;
wire  _GEN619 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN620 = io_x[40] ? _GEN16 : _GEN619;
wire  _GEN621 = io_x[2] ? _GEN11 : _GEN620;
wire  _GEN622 = io_x[15] ? _GEN2 : _GEN621;
wire  _GEN623 = io_x[42] ? _GEN5 : _GEN622;
wire  _GEN624 = io_x[43] ? _GEN623 : _GEN1;
wire  _GEN625 = io_x[38] ? _GEN624 : _GEN618;
wire  _GEN626 = io_x[17] ? _GEN625 : _GEN93;
wire  _GEN627 = io_x[39] ? _GEN626 : _GEN609;
wire  _GEN628 = io_x[37] ? _GEN627 : _GEN599;
wire  _GEN629 = io_x[77] ? _GEN282 : _GEN628;
wire  _GEN630 = io_x[78] ? _GEN629 : _GEN561;
wire  _GEN631 = io_x[79] ? _GEN630 : _GEN354;
wire  _GEN632 = io_x[69] ? _GEN52 : _GEN18;
wire  _GEN633 = io_x[16] ? _GEN17 : _GEN632;
wire  _GEN634 = io_x[40] ? _GEN633 : _GEN16;
wire  _GEN635 = io_x[2] ? _GEN11 : _GEN634;
wire  _GEN636 = io_x[15] ? _GEN2 : _GEN635;
wire  _GEN637 = io_x[42] ? _GEN636 : _GEN5;
wire  _GEN638 = io_x[43] ? _GEN1 : _GEN637;
wire  _GEN639 = io_x[38] ? _GEN8 : _GEN638;
wire  _GEN640 = io_x[18] ? _GEN32 : _GEN94;
wire  _GEN641 = io_x[4] ? _GEN79 : _GEN640;
wire  _GEN642 = io_x[30] ? _GEN20 : _GEN641;
wire  _GEN643 = io_x[69] ? _GEN642 : _GEN52;
wire  _GEN644 = io_x[16] ? _GEN17 : _GEN643;
wire  _GEN645 = io_x[40] ? _GEN644 : _GEN16;
wire  _GEN646 = io_x[2] ? _GEN645 : _GEN11;
wire  _GEN647 = io_x[7] ? _GEN97 : _GEN33;
wire  _GEN648 = io_x[18] ? _GEN94 : _GEN647;
wire  _GEN649 = io_x[4] ? _GEN79 : _GEN648;
wire  _GEN650 = io_x[30] ? _GEN20 : _GEN649;
wire  _GEN651 = io_x[69] ? _GEN650 : _GEN52;
wire  _GEN652 = io_x[16] ? _GEN17 : _GEN651;
wire  _GEN653 = io_x[40] ? _GEN652 : _GEN16;
wire  _GEN654 = io_x[18] ? _GEN32 : _GEN94;
wire  _GEN655 = io_x[4] ? _GEN79 : _GEN654;
wire  _GEN656 = io_x[30] ? _GEN19 : _GEN655;
wire  _GEN657 = io_x[69] ? _GEN656 : _GEN52;
wire  _GEN658 = io_x[16] ? _GEN17 : _GEN657;
wire  _GEN659 = io_x[40] ? _GEN658 : _GEN16;
wire  _GEN660 = io_x[2] ? _GEN659 : _GEN653;
wire  _GEN661 = io_x[15] ? _GEN660 : _GEN646;
wire  _GEN662 = io_x[42] ? _GEN661 : _GEN5;
wire  _GEN663 = io_x[43] ? _GEN662 : _GEN1;
wire  _GEN664 = io_x[38] ? _GEN8 : _GEN663;
wire  _GEN665 = io_x[17] ? _GEN664 : _GEN639;
wire  _GEN666 = io_x[18] ? _GEN32 : _GEN94;
wire  _GEN667 = io_x[4] ? _GEN79 : _GEN666;
wire  _GEN668 = io_x[30] ? _GEN667 : _GEN20;
wire  _GEN669 = io_x[69] ? _GEN668 : _GEN52;
wire  _GEN670 = io_x[16] ? _GEN17 : _GEN669;
wire  _GEN671 = io_x[40] ? _GEN670 : _GEN16;
wire  _GEN672 = io_x[2] ? _GEN671 : _GEN11;
wire  _GEN673 = io_x[31] ? _GEN236 : _GEN206;
wire  _GEN674 = io_x[19] ? _GEN34 : _GEN673;
wire  _GEN675 = io_x[70] ? _GEN674 : _GEN37;
wire  _GEN676 = io_x[7] ? _GEN97 : _GEN675;
wire  _GEN677 = io_x[18] ? _GEN94 : _GEN676;
wire  _GEN678 = io_x[4] ? _GEN79 : _GEN677;
wire  _GEN679 = io_x[30] ? _GEN678 : _GEN20;
wire  _GEN680 = io_x[69] ? _GEN679 : _GEN52;
wire  _GEN681 = io_x[16] ? _GEN17 : _GEN680;
wire  _GEN682 = io_x[40] ? _GEN681 : _GEN16;
wire  _GEN683 = io_x[18] ? _GEN32 : _GEN94;
wire  _GEN684 = io_x[4] ? _GEN79 : _GEN683;
wire  _GEN685 = io_x[18] ? _GEN32 : _GEN94;
wire  _GEN686 = io_x[4] ? _GEN79 : _GEN685;
wire  _GEN687 = io_x[30] ? _GEN686 : _GEN684;
wire  _GEN688 = io_x[69] ? _GEN687 : _GEN52;
wire  _GEN689 = io_x[16] ? _GEN17 : _GEN688;
wire  _GEN690 = io_x[40] ? _GEN689 : _GEN16;
wire  _GEN691 = io_x[2] ? _GEN690 : _GEN682;
wire  _GEN692 = io_x[15] ? _GEN691 : _GEN672;
wire  _GEN693 = io_x[42] ? _GEN692 : _GEN5;
wire  _GEN694 = io_x[43] ? _GEN1 : _GEN693;
wire  _GEN695 = io_x[38] ? _GEN694 : _GEN8;
wire  _GEN696 = io_x[17] ? _GEN695 : _GEN93;
wire  _GEN697 = io_x[39] ? _GEN696 : _GEN665;
wire  _GEN698 = io_x[7] ? _GEN97 : _GEN33;
wire  _GEN699 = io_x[18] ? _GEN94 : _GEN698;
wire  _GEN700 = io_x[4] ? _GEN699 : _GEN79;
wire  _GEN701 = io_x[30] ? _GEN700 : _GEN20;
wire  _GEN702 = io_x[69] ? _GEN52 : _GEN701;
wire  _GEN703 = io_x[16] ? _GEN702 : _GEN17;
wire  _GEN704 = io_x[40] ? _GEN703 : _GEN16;
wire  _GEN705 = io_x[2] ? _GEN11 : _GEN704;
wire  _GEN706 = io_x[15] ? _GEN2 : _GEN705;
wire  _GEN707 = io_x[42] ? _GEN5 : _GEN706;
wire  _GEN708 = io_x[43] ? _GEN1 : _GEN707;
wire  _GEN709 = io_x[38] ? _GEN708 : _GEN8;
wire  _GEN710 = io_x[17] ? _GEN709 : _GEN93;
wire  _GEN711 = io_x[39] ? _GEN710 : _GEN177;
wire  _GEN712 = io_x[37] ? _GEN711 : _GEN697;
wire  _GEN713 = io_x[43] ? _GEN178 : _GEN1;
wire  _GEN714 = io_x[38] ? _GEN8 : _GEN713;
wire  _GEN715 = io_x[17] ? _GEN714 : _GEN93;
wire  _GEN716 = io_x[43] ? _GEN178 : _GEN1;
wire  _GEN717 = io_x[38] ? _GEN8 : _GEN716;
wire  _GEN718 = io_x[17] ? _GEN717 : _GEN93;
wire  _GEN719 = io_x[39] ? _GEN718 : _GEN715;
wire  _GEN720 = io_x[37] ? _GEN719 : _GEN351;
wire  _GEN721 = io_x[77] ? _GEN720 : _GEN712;
wire  _GEN722 = 1'b0;
wire  _GEN723 = io_x[38] ? _GEN8 : _GEN722;
wire  _GEN724 = io_x[17] ? _GEN723 : _GEN93;
wire  _GEN725 = io_x[39] ? _GEN177 : _GEN724;
wire  _GEN726 = io_x[37] ? _GEN725 : _GEN351;
wire  _GEN727 = io_x[38] ? _GEN8 : _GEN722;
wire  _GEN728 = io_x[17] ? _GEN93 : _GEN727;
wire  _GEN729 = io_x[39] ? _GEN728 : _GEN177;
wire  _GEN730 = io_x[43] ? _GEN1 : _GEN178;
wire  _GEN731 = io_x[38] ? _GEN730 : _GEN8;
wire  _GEN732 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN733 = io_x[2] ? _GEN732 : _GEN11;
wire  _GEN734 = io_x[15] ? _GEN2 : _GEN733;
wire  _GEN735 = io_x[42] ? _GEN5 : _GEN734;
wire  _GEN736 = io_x[43] ? _GEN735 : _GEN1;
wire  _GEN737 = io_x[16] ? _GEN17 : _GEN25;
wire  _GEN738 = io_x[40] ? _GEN16 : _GEN737;
wire  _GEN739 = io_x[2] ? _GEN11 : _GEN738;
wire  _GEN740 = io_x[16] ? _GEN17 : _GEN25;
wire  _GEN741 = io_x[40] ? _GEN16 : _GEN740;
wire  _GEN742 = io_x[2] ? _GEN11 : _GEN741;
wire  _GEN743 = io_x[15] ? _GEN742 : _GEN739;
wire  _GEN744 = io_x[42] ? _GEN5 : _GEN743;
wire  _GEN745 = io_x[43] ? _GEN1 : _GEN744;
wire  _GEN746 = io_x[38] ? _GEN745 : _GEN736;
wire  _GEN747 = io_x[17] ? _GEN746 : _GEN731;
wire  _GEN748 = io_x[42] ? _GEN5 : _GEN471;
wire  _GEN749 = io_x[43] ? _GEN748 : _GEN1;
wire  _GEN750 = io_x[38] ? _GEN749 : _GEN8;
wire  _GEN751 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN752 = io_x[2] ? _GEN751 : _GEN11;
wire  _GEN753 = io_x[15] ? _GEN752 : _GEN3;
wire  _GEN754 = io_x[42] ? _GEN5 : _GEN753;
wire  _GEN755 = io_x[43] ? _GEN754 : _GEN1;
wire  _GEN756 = io_x[38] ? _GEN755 : _GEN8;
wire  _GEN757 = io_x[17] ? _GEN756 : _GEN750;
wire  _GEN758 = io_x[39] ? _GEN757 : _GEN747;
wire  _GEN759 = io_x[37] ? _GEN758 : _GEN729;
wire  _GEN760 = io_x[77] ? _GEN759 : _GEN726;
wire  _GEN761 = io_x[78] ? _GEN760 : _GEN721;
wire  _GEN762 = io_x[40] ? _GEN16 : _GEN181;
wire  _GEN763 = io_x[2] ? _GEN762 : _GEN11;
wire  _GEN764 = io_x[76] ? _GEN248 : _GEN207;
wire  _GEN765 = io_x[31] ? _GEN764 : _GEN206;
wire  _GEN766 = io_x[19] ? _GEN765 : _GEN34;
wire  _GEN767 = io_x[70] ? _GEN37 : _GEN766;
wire  _GEN768 = io_x[7] ? _GEN767 : _GEN97;
wire  _GEN769 = io_x[18] ? _GEN768 : _GEN94;
wire  _GEN770 = io_x[4] ? _GEN769 : _GEN79;
wire  _GEN771 = io_x[30] ? _GEN770 : _GEN20;
wire  _GEN772 = io_x[69] ? _GEN771 : _GEN52;
wire  _GEN773 = io_x[16] ? _GEN17 : _GEN772;
wire  _GEN774 = io_x[40] ? _GEN16 : _GEN773;
wire  _GEN775 = io_x[2] ? _GEN774 : _GEN11;
wire  _GEN776 = io_x[15] ? _GEN775 : _GEN763;
wire  _GEN777 = io_x[42] ? _GEN5 : _GEN776;
wire  _GEN778 = io_x[43] ? _GEN1 : _GEN777;
wire  _GEN779 = io_x[38] ? _GEN778 : _GEN8;
wire  _GEN780 = io_x[17] ? _GEN779 : _GEN93;
wire  _GEN781 = io_x[42] ? _GEN5 : _GEN471;
wire  _GEN782 = io_x[43] ? _GEN1 : _GEN781;
wire  _GEN783 = io_x[38] ? _GEN8 : _GEN782;
wire  _GEN784 = io_x[4] ? _GEN79 : _GEN31;
wire  _GEN785 = io_x[30] ? _GEN784 : _GEN20;
wire  _GEN786 = io_x[69] ? _GEN52 : _GEN785;
wire  _GEN787 = io_x[16] ? _GEN786 : _GEN17;
wire  _GEN788 = io_x[40] ? _GEN787 : _GEN16;
wire  _GEN789 = io_x[2] ? _GEN788 : _GEN11;
wire  _GEN790 = io_x[15] ? _GEN2 : _GEN789;
wire  _GEN791 = io_x[42] ? _GEN5 : _GEN790;
wire  _GEN792 = io_x[43] ? _GEN1 : _GEN791;
wire  _GEN793 = io_x[38] ? _GEN792 : _GEN8;
wire  _GEN794 = io_x[17] ? _GEN793 : _GEN783;
wire  _GEN795 = io_x[39] ? _GEN794 : _GEN780;
wire  _GEN796 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN797 = io_x[40] ? _GEN796 : _GEN16;
wire  _GEN798 = io_x[2] ? _GEN797 : _GEN10;
wire  _GEN799 = io_x[15] ? _GEN2 : _GEN798;
wire  _GEN800 = io_x[42] ? _GEN799 : _GEN5;
wire  _GEN801 = io_x[43] ? _GEN1 : _GEN800;
wire  _GEN802 = io_x[38] ? _GEN801 : _GEN8;
wire  _GEN803 = io_x[17] ? _GEN93 : _GEN802;
wire  _GEN804 = io_x[2] ? _GEN10 : _GEN11;
wire  _GEN805 = io_x[15] ? _GEN2 : _GEN804;
wire  _GEN806 = io_x[30] ? _GEN20 : _GEN19;
wire  _GEN807 = io_x[69] ? _GEN52 : _GEN806;
wire  _GEN808 = io_x[16] ? _GEN17 : _GEN807;
wire  _GEN809 = io_x[40] ? _GEN808 : _GEN16;
wire  _GEN810 = io_x[2] ? _GEN809 : _GEN11;
wire  _GEN811 = io_x[15] ? _GEN2 : _GEN810;
wire  _GEN812 = io_x[42] ? _GEN811 : _GEN805;
wire  _GEN813 = io_x[43] ? _GEN1 : _GEN812;
wire  _GEN814 = io_x[38] ? _GEN813 : _GEN8;
wire  _GEN815 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN816 = io_x[40] ? _GEN815 : _GEN16;
wire  _GEN817 = io_x[70] ? _GEN37 : _GEN95;
wire  _GEN818 = io_x[7] ? _GEN817 : _GEN97;
wire  _GEN819 = io_x[18] ? _GEN818 : _GEN94;
wire  _GEN820 = io_x[4] ? _GEN819 : _GEN79;
wire  _GEN821 = io_x[30] ? _GEN820 : _GEN20;
wire  _GEN822 = io_x[69] ? _GEN18 : _GEN821;
wire  _GEN823 = io_x[16] ? _GEN822 : _GEN17;
wire  _GEN824 = io_x[40] ? _GEN823 : _GEN16;
wire  _GEN825 = io_x[2] ? _GEN824 : _GEN816;
wire  _GEN826 = io_x[15] ? _GEN825 : _GEN2;
wire  _GEN827 = io_x[42] ? _GEN826 : _GEN5;
wire  _GEN828 = io_x[43] ? _GEN1 : _GEN827;
wire  _GEN829 = io_x[38] ? _GEN828 : _GEN8;
wire  _GEN830 = io_x[17] ? _GEN829 : _GEN814;
wire  _GEN831 = io_x[39] ? _GEN830 : _GEN803;
wire  _GEN832 = io_x[37] ? _GEN831 : _GEN795;
wire  _GEN833 = io_x[16] ? _GEN17 : _GEN25;
wire  _GEN834 = io_x[40] ? _GEN833 : _GEN16;
wire  _GEN835 = io_x[2] ? _GEN11 : _GEN834;
wire  _GEN836 = io_x[15] ? _GEN835 : _GEN2;
wire  _GEN837 = io_x[42] ? _GEN5 : _GEN836;
wire  _GEN838 = io_x[43] ? _GEN1 : _GEN837;
wire  _GEN839 = io_x[38] ? _GEN8 : _GEN838;
wire  _GEN840 = io_x[17] ? _GEN839 : _GEN93;
wire  _GEN841 = io_x[39] ? _GEN840 : _GEN177;
wire  _GEN842 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN843 = io_x[40] ? _GEN842 : _GEN16;
wire  _GEN844 = io_x[2] ? _GEN11 : _GEN843;
wire  _GEN845 = io_x[15] ? _GEN844 : _GEN2;
wire  _GEN846 = io_x[42] ? _GEN5 : _GEN845;
wire  _GEN847 = io_x[43] ? _GEN1 : _GEN846;
wire  _GEN848 = io_x[38] ? _GEN847 : _GEN8;
wire  _GEN849 = io_x[17] ? _GEN93 : _GEN848;
wire  _GEN850 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN851 = io_x[40] ? _GEN850 : _GEN16;
wire  _GEN852 = io_x[2] ? _GEN851 : _GEN11;
wire  _GEN853 = io_x[15] ? _GEN852 : _GEN2;
wire  _GEN854 = io_x[42] ? _GEN5 : _GEN853;
wire  _GEN855 = io_x[43] ? _GEN854 : _GEN1;
wire  _GEN856 = io_x[30] ? _GEN19 : _GEN20;
wire  _GEN857 = io_x[69] ? _GEN856 : _GEN52;
wire  _GEN858 = io_x[16] ? _GEN857 : _GEN17;
wire  _GEN859 = io_x[40] ? _GEN858 : _GEN16;
wire  _GEN860 = io_x[2] ? _GEN859 : _GEN11;
wire  _GEN861 = io_x[31] ? _GEN206 : _GEN236;
wire  _GEN862 = io_x[19] ? _GEN861 : _GEN34;
wire  _GEN863 = io_x[70] ? _GEN37 : _GEN862;
wire  _GEN864 = io_x[7] ? _GEN863 : _GEN97;
wire  _GEN865 = io_x[18] ? _GEN864 : _GEN94;
wire  _GEN866 = io_x[4] ? _GEN865 : _GEN79;
wire  _GEN867 = io_x[30] ? _GEN866 : _GEN20;
wire  _GEN868 = io_x[69] ? _GEN867 : _GEN52;
wire  _GEN869 = io_x[16] ? _GEN868 : _GEN17;
wire  _GEN870 = io_x[40] ? _GEN869 : _GEN16;
wire  _GEN871 = io_x[2] ? _GEN870 : _GEN11;
wire  _GEN872 = io_x[15] ? _GEN871 : _GEN860;
wire  _GEN873 = io_x[42] ? _GEN5 : _GEN872;
wire  _GEN874 = io_x[43] ? _GEN873 : _GEN1;
wire  _GEN875 = io_x[38] ? _GEN874 : _GEN855;
wire  _GEN876 = io_x[17] ? _GEN93 : _GEN875;
wire  _GEN877 = io_x[39] ? _GEN876 : _GEN849;
wire  _GEN878 = io_x[37] ? _GEN877 : _GEN841;
wire  _GEN879 = io_x[77] ? _GEN878 : _GEN832;
wire  _GEN880 = io_x[69] ? _GEN52 : _GEN18;
wire  _GEN881 = io_x[16] ? _GEN880 : _GEN17;
wire  _GEN882 = io_x[40] ? _GEN881 : _GEN16;
wire  _GEN883 = io_x[2] ? _GEN11 : _GEN882;
wire  _GEN884 = io_x[15] ? _GEN2 : _GEN883;
wire  _GEN885 = io_x[42] ? _GEN884 : _GEN5;
wire  _GEN886 = io_x[43] ? _GEN1 : _GEN885;
wire  _GEN887 = io_x[38] ? _GEN886 : _GEN8;
wire  _GEN888 = io_x[40] ? _GEN16 : _GEN181;
wire  _GEN889 = io_x[2] ? _GEN11 : _GEN888;
wire  _GEN890 = io_x[15] ? _GEN2 : _GEN889;
wire  _GEN891 = io_x[42] ? _GEN5 : _GEN890;
wire  _GEN892 = io_x[43] ? _GEN1 : _GEN891;
wire  _GEN893 = io_x[38] ? _GEN8 : _GEN892;
wire  _GEN894 = io_x[17] ? _GEN893 : _GEN887;
wire  _GEN895 = io_x[39] ? _GEN894 : _GEN177;
wire  _GEN896 = io_x[4] ? _GEN79 : _GEN31;
wire  _GEN897 = io_x[30] ? _GEN20 : _GEN896;
wire  _GEN898 = io_x[69] ? _GEN897 : _GEN52;
wire  _GEN899 = io_x[16] ? _GEN898 : _GEN17;
wire  _GEN900 = io_x[40] ? _GEN899 : _GEN16;
wire  _GEN901 = io_x[69] ? _GEN52 : _GEN18;
wire  _GEN902 = io_x[16] ? _GEN17 : _GEN901;
wire  _GEN903 = io_x[40] ? _GEN902 : _GEN16;
wire  _GEN904 = io_x[2] ? _GEN903 : _GEN900;
wire  _GEN905 = io_x[15] ? _GEN2 : _GEN904;
wire  _GEN906 = io_x[42] ? _GEN5 : _GEN905;
wire  _GEN907 = io_x[43] ? _GEN1 : _GEN906;
wire  _GEN908 = io_x[2] ? _GEN10 : _GEN11;
wire  _GEN909 = io_x[15] ? _GEN2 : _GEN908;
wire  _GEN910 = io_x[42] ? _GEN5 : _GEN909;
wire  _GEN911 = io_x[43] ? _GEN1 : _GEN910;
wire  _GEN912 = io_x[38] ? _GEN911 : _GEN907;
wire  _GEN913 = io_x[17] ? _GEN912 : _GEN93;
wire  _GEN914 = io_x[42] ? _GEN471 : _GEN5;
wire  _GEN915 = io_x[43] ? _GEN914 : _GEN1;
wire  _GEN916 = io_x[2] ? _GEN10 : _GEN11;
wire  _GEN917 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN918 = io_x[40] ? _GEN16 : _GEN917;
wire  _GEN919 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN920 = io_x[40] ? _GEN16 : _GEN919;
wire  _GEN921 = io_x[2] ? _GEN920 : _GEN918;
wire  _GEN922 = io_x[15] ? _GEN921 : _GEN916;
wire  _GEN923 = io_x[42] ? _GEN5 : _GEN922;
wire  _GEN924 = io_x[43] ? _GEN1 : _GEN923;
wire  _GEN925 = io_x[38] ? _GEN924 : _GEN915;
wire  _GEN926 = io_x[31] ? _GEN236 : _GEN206;
wire  _GEN927 = io_x[19] ? _GEN926 : _GEN34;
wire  _GEN928 = io_x[70] ? _GEN927 : _GEN37;
wire  _GEN929 = io_x[7] ? _GEN928 : _GEN97;
wire  _GEN930 = io_x[18] ? _GEN929 : _GEN94;
wire  _GEN931 = io_x[4] ? _GEN79 : _GEN930;
wire  _GEN932 = io_x[30] ? _GEN931 : _GEN20;
wire  _GEN933 = io_x[69] ? _GEN932 : _GEN52;
wire  _GEN934 = io_x[16] ? _GEN933 : _GEN17;
wire  _GEN935 = io_x[40] ? _GEN16 : _GEN934;
wire  _GEN936 = io_x[2] ? _GEN935 : _GEN11;
wire  _GEN937 = io_x[15] ? _GEN936 : _GEN2;
wire  _GEN938 = io_x[42] ? _GEN5 : _GEN937;
wire  _GEN939 = io_x[43] ? _GEN1 : _GEN938;
wire  _GEN940 = io_x[38] ? _GEN939 : _GEN8;
wire  _GEN941 = io_x[17] ? _GEN940 : _GEN925;
wire  _GEN942 = io_x[39] ? _GEN941 : _GEN913;
wire  _GEN943 = io_x[37] ? _GEN942 : _GEN895;
wire  _GEN944 = io_x[69] ? _GEN52 : _GEN18;
wire  _GEN945 = io_x[16] ? _GEN944 : _GEN17;
wire  _GEN946 = io_x[40] ? _GEN945 : _GEN16;
wire  _GEN947 = io_x[2] ? _GEN946 : _GEN11;
wire  _GEN948 = io_x[15] ? _GEN3 : _GEN947;
wire  _GEN949 = io_x[42] ? _GEN5 : _GEN948;
wire  _GEN950 = io_x[43] ? _GEN949 : _GEN1;
wire  _GEN951 = io_x[38] ? _GEN8 : _GEN950;
wire  _GEN952 = io_x[17] ? _GEN951 : _GEN93;
wire  _GEN953 = io_x[39] ? _GEN952 : _GEN177;
wire  _GEN954 = io_x[37] ? _GEN953 : _GEN351;
wire  _GEN955 = io_x[77] ? _GEN954 : _GEN943;
wire  _GEN956 = io_x[78] ? _GEN955 : _GEN879;
wire  _GEN957 = io_x[79] ? _GEN956 : _GEN761;
wire  _GEN958 = io_x[80] ? _GEN957 : _GEN631;
wire  _GEN959 = io_x[69] ? _GEN52 : _GEN18;
wire  _GEN960 = io_x[16] ? _GEN959 : _GEN17;
wire  _GEN961 = io_x[40] ? _GEN960 : _GEN16;
wire  _GEN962 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN963 = io_x[40] ? _GEN962 : _GEN16;
wire  _GEN964 = io_x[2] ? _GEN963 : _GEN961;
wire  _GEN965 = io_x[15] ? _GEN964 : _GEN2;
wire  _GEN966 = io_x[42] ? _GEN5 : _GEN965;
wire  _GEN967 = io_x[43] ? _GEN966 : _GEN1;
wire  _GEN968 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN969 = io_x[2] ? _GEN968 : _GEN11;
wire  _GEN970 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN971 = io_x[40] ? _GEN970 : _GEN16;
wire  _GEN972 = io_x[2] ? _GEN971 : _GEN11;
wire  _GEN973 = io_x[15] ? _GEN972 : _GEN969;
wire  _GEN974 = io_x[42] ? _GEN5 : _GEN973;
wire  _GEN975 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN976 = io_x[40] ? _GEN975 : _GEN16;
wire  _GEN977 = io_x[2] ? _GEN976 : _GEN11;
wire  _GEN978 = io_x[31] ? _GEN206 : _GEN236;
wire  _GEN979 = io_x[19] ? _GEN978 : _GEN34;
wire  _GEN980 = io_x[70] ? _GEN37 : _GEN979;
wire  _GEN981 = io_x[7] ? _GEN980 : _GEN97;
wire  _GEN982 = io_x[18] ? _GEN981 : _GEN94;
wire  _GEN983 = io_x[4] ? _GEN982 : _GEN31;
wire  _GEN984 = io_x[30] ? _GEN983 : _GEN20;
wire  _GEN985 = io_x[69] ? _GEN52 : _GEN984;
wire  _GEN986 = io_x[16] ? _GEN985 : _GEN17;
wire  _GEN987 = io_x[40] ? _GEN986 : _GEN16;
wire  _GEN988 = io_x[2] ? _GEN987 : _GEN11;
wire  _GEN989 = io_x[15] ? _GEN988 : _GEN977;
wire  _GEN990 = io_x[42] ? _GEN5 : _GEN989;
wire  _GEN991 = io_x[43] ? _GEN990 : _GEN974;
wire  _GEN992 = io_x[38] ? _GEN991 : _GEN967;
wire  _GEN993 = io_x[30] ? _GEN20 : _GEN19;
wire  _GEN994 = io_x[69] ? _GEN993 : _GEN52;
wire  _GEN995 = io_x[16] ? _GEN994 : _GEN17;
wire  _GEN996 = io_x[40] ? _GEN995 : _GEN16;
wire  _GEN997 = io_x[2] ? _GEN996 : _GEN11;
wire  _GEN998 = io_x[15] ? _GEN997 : _GEN2;
wire  _GEN999 = io_x[42] ? _GEN5 : _GEN998;
wire  _GEN1000 = io_x[69] ? _GEN18 : _GEN52;
wire  _GEN1001 = io_x[16] ? _GEN17 : _GEN1000;
wire  _GEN1002 = io_x[40] ? _GEN1001 : _GEN16;
wire  _GEN1003 = io_x[2] ? _GEN1002 : _GEN11;
wire  _GEN1004 = io_x[15] ? _GEN2 : _GEN1003;
wire  _GEN1005 = io_x[42] ? _GEN5 : _GEN1004;
wire  _GEN1006 = io_x[43] ? _GEN1005 : _GEN999;
wire  _GEN1007 = io_x[38] ? _GEN1006 : _GEN8;
wire  _GEN1008 = io_x[17] ? _GEN1007 : _GEN992;
wire  _GEN1009 = io_x[30] ? _GEN19 : _GEN20;
wire  _GEN1010 = io_x[69] ? _GEN52 : _GEN1009;
wire  _GEN1011 = io_x[16] ? _GEN1010 : _GEN17;
wire  _GEN1012 = io_x[40] ? _GEN1011 : _GEN181;
wire  _GEN1013 = io_x[2] ? _GEN1012 : _GEN10;
wire  _GEN1014 = io_x[15] ? _GEN1013 : _GEN2;
wire  _GEN1015 = io_x[42] ? _GEN5 : _GEN1014;
wire  _GEN1016 = io_x[30] ? _GEN20 : _GEN19;
wire  _GEN1017 = io_x[69] ? _GEN1016 : _GEN52;
wire  _GEN1018 = io_x[16] ? _GEN17 : _GEN1017;
wire  _GEN1019 = io_x[40] ? _GEN1018 : _GEN16;
wire  _GEN1020 = io_x[2] ? _GEN11 : _GEN1019;
wire  _GEN1021 = io_x[15] ? _GEN1020 : _GEN2;
wire  _GEN1022 = io_x[30] ? _GEN20 : _GEN19;
wire  _GEN1023 = io_x[69] ? _GEN1022 : _GEN52;
wire  _GEN1024 = io_x[16] ? _GEN1023 : _GEN17;
wire  _GEN1025 = io_x[40] ? _GEN1024 : _GEN16;
wire  _GEN1026 = io_x[2] ? _GEN1025 : _GEN11;
wire  _GEN1027 = io_x[15] ? _GEN1026 : _GEN2;
wire  _GEN1028 = io_x[42] ? _GEN1027 : _GEN1021;
wire  _GEN1029 = io_x[43] ? _GEN1028 : _GEN1015;
wire  _GEN1030 = io_x[38] ? _GEN8 : _GEN1029;
wire  _GEN1031 = io_x[30] ? _GEN20 : _GEN19;
wire  _GEN1032 = io_x[69] ? _GEN52 : _GEN1031;
wire  _GEN1033 = io_x[16] ? _GEN1032 : _GEN17;
wire  _GEN1034 = io_x[40] ? _GEN16 : _GEN1033;
wire  _GEN1035 = io_x[2] ? _GEN11 : _GEN1034;
wire  _GEN1036 = io_x[15] ? _GEN1035 : _GEN2;
wire  _GEN1037 = io_x[42] ? _GEN5 : _GEN1036;
wire  _GEN1038 = io_x[43] ? _GEN1037 : _GEN1;
wire  _GEN1039 = io_x[18] ? _GEN32 : _GEN94;
wire  _GEN1040 = io_x[4] ? _GEN1039 : _GEN79;
wire  _GEN1041 = io_x[30] ? _GEN1040 : _GEN20;
wire  _GEN1042 = io_x[69] ? _GEN52 : _GEN1041;
wire  _GEN1043 = io_x[16] ? _GEN1042 : _GEN17;
wire  _GEN1044 = io_x[40] ? _GEN16 : _GEN1043;
wire  _GEN1045 = io_x[2] ? _GEN1044 : _GEN11;
wire  _GEN1046 = io_x[15] ? _GEN1045 : _GEN2;
wire  _GEN1047 = io_x[42] ? _GEN5 : _GEN1046;
wire  _GEN1048 = io_x[43] ? _GEN1 : _GEN1047;
wire  _GEN1049 = io_x[38] ? _GEN1048 : _GEN1038;
wire  _GEN1050 = io_x[17] ? _GEN1049 : _GEN1030;
wire  _GEN1051 = io_x[39] ? _GEN1050 : _GEN1008;
wire  _GEN1052 = io_x[16] ? _GEN17 : _GEN25;
wire  _GEN1053 = io_x[40] ? _GEN1052 : _GEN16;
wire  _GEN1054 = io_x[2] ? _GEN11 : _GEN1053;
wire  _GEN1055 = io_x[15] ? _GEN2 : _GEN1054;
wire  _GEN1056 = io_x[42] ? _GEN5 : _GEN1055;
wire  _GEN1057 = io_x[43] ? _GEN1056 : _GEN1;
wire  _GEN1058 = io_x[40] ? _GEN16 : _GEN181;
wire  _GEN1059 = io_x[2] ? _GEN1058 : _GEN10;
wire  _GEN1060 = io_x[15] ? _GEN3 : _GEN1059;
wire  _GEN1061 = io_x[42] ? _GEN5 : _GEN1060;
wire  _GEN1062 = io_x[40] ? _GEN16 : _GEN181;
wire  _GEN1063 = io_x[2] ? _GEN11 : _GEN1062;
wire  _GEN1064 = io_x[15] ? _GEN2 : _GEN1063;
wire  _GEN1065 = io_x[42] ? _GEN5 : _GEN1064;
wire  _GEN1066 = io_x[43] ? _GEN1065 : _GEN1061;
wire  _GEN1067 = io_x[38] ? _GEN1066 : _GEN1057;
wire  _GEN1068 = io_x[42] ? _GEN5 : _GEN471;
wire  _GEN1069 = io_x[4] ? _GEN79 : _GEN31;
wire  _GEN1070 = io_x[30] ? _GEN1069 : _GEN20;
wire  _GEN1071 = io_x[69] ? _GEN52 : _GEN1070;
wire  _GEN1072 = io_x[16] ? _GEN17 : _GEN1071;
wire  _GEN1073 = io_x[40] ? _GEN16 : _GEN1072;
wire  _GEN1074 = io_x[2] ? _GEN1073 : _GEN11;
wire  _GEN1075 = io_x[15] ? _GEN1074 : _GEN2;
wire  _GEN1076 = io_x[42] ? _GEN5 : _GEN1075;
wire  _GEN1077 = io_x[43] ? _GEN1076 : _GEN1068;
wire  _GEN1078 = io_x[38] ? _GEN1077 : _GEN8;
wire  _GEN1079 = io_x[17] ? _GEN1078 : _GEN1067;
wire  _GEN1080 = io_x[2] ? _GEN10 : _GEN11;
wire  _GEN1081 = io_x[15] ? _GEN2 : _GEN1080;
wire  _GEN1082 = io_x[42] ? _GEN5 : _GEN1081;
wire  _GEN1083 = io_x[43] ? _GEN1082 : _GEN1;
wire  _GEN1084 = io_x[38] ? _GEN1083 : _GEN8;
wire  _GEN1085 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN1086 = io_x[40] ? _GEN1085 : _GEN16;
wire  _GEN1087 = io_x[2] ? _GEN11 : _GEN1086;
wire  _GEN1088 = io_x[69] ? _GEN52 : _GEN18;
wire  _GEN1089 = io_x[16] ? _GEN1088 : _GEN17;
wire  _GEN1090 = io_x[40] ? _GEN1089 : _GEN16;
wire  _GEN1091 = io_x[2] ? _GEN1090 : _GEN11;
wire  _GEN1092 = io_x[15] ? _GEN1091 : _GEN1087;
wire  _GEN1093 = io_x[42] ? _GEN5 : _GEN1092;
wire  _GEN1094 = io_x[43] ? _GEN1093 : _GEN1;
wire  _GEN1095 = io_x[16] ? _GEN17 : _GEN25;
wire  _GEN1096 = io_x[40] ? _GEN1095 : _GEN16;
wire  _GEN1097 = io_x[2] ? _GEN1096 : _GEN11;
wire  _GEN1098 = io_x[15] ? _GEN2 : _GEN1097;
wire  _GEN1099 = io_x[42] ? _GEN5 : _GEN1098;
wire  _GEN1100 = io_x[43] ? _GEN1099 : _GEN1;
wire  _GEN1101 = io_x[38] ? _GEN1100 : _GEN1094;
wire  _GEN1102 = io_x[17] ? _GEN1101 : _GEN1084;
wire  _GEN1103 = io_x[39] ? _GEN1102 : _GEN1079;
wire  _GEN1104 = io_x[37] ? _GEN1103 : _GEN1051;
wire  _GEN1105 = io_x[40] ? _GEN16 : _GEN181;
wire  _GEN1106 = io_x[2] ? _GEN11 : _GEN1105;
wire  _GEN1107 = io_x[15] ? _GEN2 : _GEN1106;
wire  _GEN1108 = io_x[42] ? _GEN1107 : _GEN5;
wire  _GEN1109 = io_x[43] ? _GEN1 : _GEN1108;
wire  _GEN1110 = io_x[38] ? _GEN8 : _GEN1109;
wire  _GEN1111 = io_x[17] ? _GEN93 : _GEN1110;
wire  _GEN1112 = io_x[39] ? _GEN1111 : _GEN177;
wire  _GEN1113 = io_x[15] ? _GEN2 : _GEN3;
wire  _GEN1114 = io_x[42] ? _GEN5 : _GEN1113;
wire  _GEN1115 = io_x[43] ? _GEN1 : _GEN1114;
wire  _GEN1116 = io_x[16] ? _GEN25 : _GEN17;
wire  _GEN1117 = io_x[40] ? _GEN16 : _GEN1116;
wire  _GEN1118 = io_x[2] ? _GEN11 : _GEN1117;
wire  _GEN1119 = io_x[15] ? _GEN2 : _GEN1118;
wire  _GEN1120 = io_x[42] ? _GEN1119 : _GEN5;
wire  _GEN1121 = io_x[43] ? _GEN1 : _GEN1120;
wire  _GEN1122 = io_x[38] ? _GEN1121 : _GEN1115;
wire  _GEN1123 = io_x[30] ? _GEN19 : _GEN20;
wire  _GEN1124 = io_x[69] ? _GEN52 : _GEN1123;
wire  _GEN1125 = io_x[16] ? _GEN1124 : _GEN25;
wire  _GEN1126 = io_x[40] ? _GEN1125 : _GEN16;
wire  _GEN1127 = io_x[2] ? _GEN11 : _GEN1126;
wire  _GEN1128 = io_x[15] ? _GEN2 : _GEN1127;
wire  _GEN1129 = io_x[42] ? _GEN5 : _GEN1128;
wire  _GEN1130 = io_x[43] ? _GEN1 : _GEN1129;
wire  _GEN1131 = io_x[18] ? _GEN94 : _GEN32;
wire  _GEN1132 = io_x[4] ? _GEN1131 : _GEN79;
wire  _GEN1133 = io_x[30] ? _GEN1132 : _GEN20;
wire  _GEN1134 = io_x[69] ? _GEN52 : _GEN1133;
wire  _GEN1135 = io_x[16] ? _GEN1134 : _GEN17;
wire  _GEN1136 = io_x[40] ? _GEN16 : _GEN1135;
wire  _GEN1137 = io_x[2] ? _GEN1136 : _GEN11;
wire  _GEN1138 = io_x[15] ? _GEN2 : _GEN1137;
wire  _GEN1139 = io_x[42] ? _GEN1138 : _GEN5;
wire  _GEN1140 = io_x[43] ? _GEN1 : _GEN1139;
wire  _GEN1141 = io_x[38] ? _GEN1140 : _GEN1130;
wire  _GEN1142 = io_x[17] ? _GEN1141 : _GEN1122;
wire  _GEN1143 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN1144 = io_x[2] ? _GEN11 : _GEN1143;
wire  _GEN1145 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN1146 = io_x[2] ? _GEN11 : _GEN1145;
wire  _GEN1147 = io_x[15] ? _GEN1146 : _GEN1144;
wire  _GEN1148 = io_x[42] ? _GEN1147 : _GEN5;
wire  _GEN1149 = io_x[43] ? _GEN1 : _GEN1148;
wire  _GEN1150 = io_x[38] ? _GEN1149 : _GEN8;
wire  _GEN1151 = io_x[17] ? _GEN1150 : _GEN93;
wire  _GEN1152 = io_x[39] ? _GEN1151 : _GEN1142;
wire  _GEN1153 = io_x[37] ? _GEN1152 : _GEN1112;
wire  _GEN1154 = io_x[77] ? _GEN1153 : _GEN1104;
wire  _GEN1155 = io_x[43] ? _GEN178 : _GEN1;
wire  _GEN1156 = io_x[38] ? _GEN1155 : _GEN8;
wire  _GEN1157 = io_x[2] ? _GEN10 : _GEN11;
wire  _GEN1158 = io_x[2] ? _GEN10 : _GEN11;
wire  _GEN1159 = io_x[15] ? _GEN1158 : _GEN1157;
wire  _GEN1160 = io_x[42] ? _GEN5 : _GEN1159;
wire  _GEN1161 = io_x[43] ? _GEN1160 : _GEN1;
wire  _GEN1162 = io_x[16] ? _GEN17 : _GEN25;
wire  _GEN1163 = io_x[40] ? _GEN16 : _GEN1162;
wire  _GEN1164 = io_x[19] ? _GEN34 : _GEN35;
wire  _GEN1165 = io_x[70] ? _GEN37 : _GEN1164;
wire  _GEN1166 = io_x[7] ? _GEN1165 : _GEN97;
wire  _GEN1167 = io_x[18] ? _GEN1166 : _GEN94;
wire  _GEN1168 = io_x[4] ? _GEN1167 : _GEN79;
wire  _GEN1169 = io_x[30] ? _GEN20 : _GEN1168;
wire  _GEN1170 = io_x[69] ? _GEN1169 : _GEN52;
wire  _GEN1171 = io_x[16] ? _GEN1170 : _GEN25;
wire  _GEN1172 = io_x[40] ? _GEN16 : _GEN1171;
wire  _GEN1173 = io_x[2] ? _GEN1172 : _GEN1163;
wire  _GEN1174 = io_x[15] ? _GEN3 : _GEN1173;
wire  _GEN1175 = io_x[42] ? _GEN5 : _GEN1174;
wire  _GEN1176 = io_x[43] ? _GEN1175 : _GEN1;
wire  _GEN1177 = io_x[38] ? _GEN1176 : _GEN1161;
wire  _GEN1178 = io_x[17] ? _GEN1177 : _GEN1156;
wire  _GEN1179 = io_x[39] ? _GEN177 : _GEN1178;
wire  _GEN1180 = io_x[38] ? _GEN8 : _GEN722;
wire  _GEN1181 = io_x[40] ? _GEN16 : _GEN181;
wire  _GEN1182 = io_x[2] ? _GEN1181 : _GEN10;
wire  _GEN1183 = io_x[40] ? _GEN16 : _GEN181;
wire  _GEN1184 = io_x[2] ? _GEN1183 : _GEN10;
wire  _GEN1185 = io_x[15] ? _GEN1184 : _GEN1182;
wire  _GEN1186 = io_x[42] ? _GEN5 : _GEN1185;
wire  _GEN1187 = io_x[43] ? _GEN1186 : _GEN1;
wire  _GEN1188 = io_x[38] ? _GEN8 : _GEN1187;
wire  _GEN1189 = io_x[17] ? _GEN1188 : _GEN1180;
wire  _GEN1190 = io_x[16] ? _GEN17 : _GEN25;
wire  _GEN1191 = io_x[40] ? _GEN16 : _GEN1190;
wire  _GEN1192 = io_x[2] ? _GEN11 : _GEN1191;
wire  _GEN1193 = io_x[15] ? _GEN3 : _GEN1192;
wire  _GEN1194 = io_x[42] ? _GEN1193 : _GEN5;
wire  _GEN1195 = io_x[43] ? _GEN1194 : _GEN1;
wire  _GEN1196 = io_x[15] ? _GEN3 : _GEN2;
wire  _GEN1197 = io_x[42] ? _GEN1196 : _GEN5;
wire  _GEN1198 = io_x[43] ? _GEN1197 : _GEN1;
wire  _GEN1199 = io_x[38] ? _GEN1198 : _GEN1195;
wire  _GEN1200 = io_x[17] ? _GEN93 : _GEN1199;
wire  _GEN1201 = io_x[39] ? _GEN1200 : _GEN1189;
wire  _GEN1202 = io_x[37] ? _GEN1201 : _GEN1179;
wire  _GEN1203 = io_x[2] ? _GEN10 : _GEN11;
wire  _GEN1204 = io_x[15] ? _GEN2 : _GEN1203;
wire  _GEN1205 = io_x[42] ? _GEN5 : _GEN1204;
wire  _GEN1206 = io_x[4] ? _GEN79 : _GEN31;
wire  _GEN1207 = io_x[30] ? _GEN19 : _GEN1206;
wire  _GEN1208 = io_x[69] ? _GEN1207 : _GEN52;
wire  _GEN1209 = io_x[16] ? _GEN17 : _GEN1208;
wire  _GEN1210 = io_x[40] ? _GEN16 : _GEN1209;
wire  _GEN1211 = io_x[2] ? _GEN1210 : _GEN11;
wire  _GEN1212 = io_x[15] ? _GEN2 : _GEN1211;
wire  _GEN1213 = io_x[42] ? _GEN1212 : _GEN5;
wire  _GEN1214 = io_x[43] ? _GEN1213 : _GEN1205;
wire  _GEN1215 = io_x[15] ? _GEN2 : _GEN3;
wire  _GEN1216 = io_x[42] ? _GEN5 : _GEN1215;
wire  _GEN1217 = io_x[43] ? _GEN1216 : _GEN1;
wire  _GEN1218 = io_x[38] ? _GEN1217 : _GEN1214;
wire  _GEN1219 = io_x[17] ? _GEN1218 : _GEN93;
wire  _GEN1220 = io_x[39] ? _GEN177 : _GEN1219;
wire  _GEN1221 = io_x[18] ? _GEN94 : _GEN32;
wire  _GEN1222 = io_x[4] ? _GEN79 : _GEN1221;
wire  _GEN1223 = io_x[30] ? _GEN20 : _GEN1222;
wire  _GEN1224 = io_x[69] ? _GEN1223 : _GEN52;
wire  _GEN1225 = io_x[16] ? _GEN1224 : _GEN17;
wire  _GEN1226 = io_x[40] ? _GEN1225 : _GEN16;
wire  _GEN1227 = io_x[2] ? _GEN11 : _GEN1226;
wire  _GEN1228 = io_x[15] ? _GEN2 : _GEN1227;
wire  _GEN1229 = io_x[7] ? _GEN33 : _GEN97;
wire  _GEN1230 = io_x[18] ? _GEN94 : _GEN1229;
wire  _GEN1231 = io_x[4] ? _GEN1230 : _GEN79;
wire  _GEN1232 = io_x[4] ? _GEN31 : _GEN79;
wire  _GEN1233 = io_x[30] ? _GEN1232 : _GEN1231;
wire  _GEN1234 = io_x[69] ? _GEN1233 : _GEN52;
wire  _GEN1235 = io_x[16] ? _GEN17 : _GEN1234;
wire  _GEN1236 = io_x[40] ? _GEN16 : _GEN1235;
wire  _GEN1237 = io_x[7] ? _GEN97 : _GEN33;
wire  _GEN1238 = io_x[18] ? _GEN32 : _GEN1237;
wire  _GEN1239 = io_x[4] ? _GEN79 : _GEN1238;
wire  _GEN1240 = io_x[30] ? _GEN20 : _GEN1239;
wire  _GEN1241 = io_x[69] ? _GEN1240 : _GEN52;
wire  _GEN1242 = io_x[16] ? _GEN17 : _GEN1241;
wire  _GEN1243 = io_x[40] ? _GEN16 : _GEN1242;
wire  _GEN1244 = io_x[2] ? _GEN1243 : _GEN1236;
wire  _GEN1245 = io_x[4] ? _GEN31 : _GEN79;
wire  _GEN1246 = io_x[30] ? _GEN1245 : _GEN20;
wire  _GEN1247 = io_x[69] ? _GEN1246 : _GEN52;
wire  _GEN1248 = io_x[16] ? _GEN17 : _GEN1247;
wire  _GEN1249 = io_x[40] ? _GEN16 : _GEN1248;
wire  _GEN1250 = io_x[4] ? _GEN79 : _GEN31;
wire  _GEN1251 = io_x[70] ? _GEN95 : _GEN37;
wire  _GEN1252 = io_x[7] ? _GEN1251 : _GEN97;
wire  _GEN1253 = io_x[18] ? _GEN94 : _GEN1252;
wire  _GEN1254 = io_x[4] ? _GEN1253 : _GEN31;
wire  _GEN1255 = io_x[30] ? _GEN1254 : _GEN1250;
wire  _GEN1256 = io_x[69] ? _GEN1255 : _GEN52;
wire  _GEN1257 = io_x[16] ? _GEN17 : _GEN1256;
wire  _GEN1258 = io_x[40] ? _GEN16 : _GEN1257;
wire  _GEN1259 = io_x[2] ? _GEN1258 : _GEN1249;
wire  _GEN1260 = io_x[15] ? _GEN1259 : _GEN1244;
wire  _GEN1261 = io_x[42] ? _GEN1260 : _GEN1228;
wire  _GEN1262 = io_x[43] ? _GEN1261 : _GEN1;
wire  _GEN1263 = io_x[38] ? _GEN8 : _GEN1262;
wire  _GEN1264 = io_x[17] ? _GEN93 : _GEN1263;
wire  _GEN1265 = io_x[43] ? _GEN178 : _GEN1;
wire  _GEN1266 = io_x[38] ? _GEN8 : _GEN1265;
wire  _GEN1267 = io_x[43] ? _GEN178 : _GEN1;
wire  _GEN1268 = io_x[38] ? _GEN8 : _GEN1267;
wire  _GEN1269 = io_x[17] ? _GEN1268 : _GEN1266;
wire  _GEN1270 = io_x[39] ? _GEN1269 : _GEN1264;
wire  _GEN1271 = io_x[37] ? _GEN1270 : _GEN1220;
wire  _GEN1272 = io_x[77] ? _GEN1271 : _GEN1202;
wire  _GEN1273 = io_x[78] ? _GEN1272 : _GEN1154;
wire  _GEN1274 = io_x[69] ? _GEN18 : _GEN52;
wire  _GEN1275 = io_x[16] ? _GEN1274 : _GEN17;
wire  _GEN1276 = io_x[40] ? _GEN16 : _GEN1275;
wire  _GEN1277 = io_x[2] ? _GEN11 : _GEN1276;
wire  _GEN1278 = io_x[15] ? _GEN2 : _GEN1277;
wire  _GEN1279 = io_x[42] ? _GEN5 : _GEN1278;
wire  _GEN1280 = io_x[43] ? _GEN1 : _GEN1279;
wire  _GEN1281 = io_x[38] ? _GEN8 : _GEN1280;
wire  _GEN1282 = io_x[42] ? _GEN471 : _GEN5;
wire  _GEN1283 = io_x[43] ? _GEN1 : _GEN1282;
wire  _GEN1284 = io_x[2] ? _GEN10 : _GEN11;
wire  _GEN1285 = io_x[15] ? _GEN3 : _GEN1284;
wire  _GEN1286 = io_x[42] ? _GEN5 : _GEN1285;
wire  _GEN1287 = io_x[43] ? _GEN1286 : _GEN1;
wire  _GEN1288 = io_x[38] ? _GEN1287 : _GEN1283;
wire  _GEN1289 = io_x[17] ? _GEN1288 : _GEN1281;
wire  _GEN1290 = io_x[39] ? _GEN177 : _GEN1289;
wire  _GEN1291 = io_x[40] ? _GEN181 : _GEN16;
wire  _GEN1292 = io_x[2] ? _GEN11 : _GEN1291;
wire  _GEN1293 = io_x[15] ? _GEN2 : _GEN1292;
wire  _GEN1294 = io_x[42] ? _GEN5 : _GEN1293;
wire  _GEN1295 = io_x[43] ? _GEN1294 : _GEN1;
wire  _GEN1296 = io_x[38] ? _GEN8 : _GEN1295;
wire  _GEN1297 = io_x[19] ? _GEN34 : _GEN35;
wire  _GEN1298 = io_x[70] ? _GEN37 : _GEN1297;
wire  _GEN1299 = io_x[7] ? _GEN97 : _GEN1298;
wire  _GEN1300 = io_x[18] ? _GEN1299 : _GEN94;
wire  _GEN1301 = io_x[4] ? _GEN79 : _GEN1300;
wire  _GEN1302 = io_x[30] ? _GEN20 : _GEN1301;
wire  _GEN1303 = io_x[69] ? _GEN1302 : _GEN52;
wire  _GEN1304 = io_x[16] ? _GEN1303 : _GEN17;
wire  _GEN1305 = io_x[40] ? _GEN1304 : _GEN16;
wire  _GEN1306 = io_x[2] ? _GEN11 : _GEN1305;
wire  _GEN1307 = io_x[15] ? _GEN2 : _GEN1306;
wire  _GEN1308 = io_x[42] ? _GEN1307 : _GEN5;
wire  _GEN1309 = io_x[43] ? _GEN1308 : _GEN1;
wire  _GEN1310 = io_x[38] ? _GEN1309 : _GEN8;
wire  _GEN1311 = io_x[17] ? _GEN1310 : _GEN1296;
wire  _GEN1312 = io_x[39] ? _GEN177 : _GEN1311;
wire  _GEN1313 = io_x[37] ? _GEN1312 : _GEN1290;
wire  _GEN1314 = io_x[77] ? _GEN1313 : _GEN282;
wire  _GEN1315 = 1'b1;
wire  _GEN1316 = io_x[78] ? _GEN1315 : _GEN1314;
wire  _GEN1317 = io_x[79] ? _GEN1316 : _GEN1273;
wire  _GEN1318 = 1'b1;
wire  _GEN1319 = io_x[80] ? _GEN1318 : _GEN1317;
wire  _GEN1320 = io_x[81] ? _GEN1319 : _GEN958;
wire  _GEN1321 = 1'b1;
wire  _GEN1322 = io_x[82] ? _GEN1321 : _GEN1320;
wire  _GEN1323 = 1'b1;
wire  _GEN1324 = io_x[83] ? _GEN1323 : _GEN1322;
wire  _GEN1325 = 1'b1;
wire  _GEN1326 = io_x[84] ? _GEN1325 : _GEN1324;
wire  _GEN1327 = 1'b1;
wire  _GEN1328 = io_x[85] ? _GEN1327 : _GEN1326;
wire  _GEN1329 = 1'b1;
wire  _GEN1330 = io_x[86] ? _GEN1329 : _GEN1328;
wire  _GEN1331 = 1'b1;
wire  _GEN1332 = io_x[87] ? _GEN1331 : _GEN1330;
wire  _GEN1333 = 1'b1;
wire  _GEN1334 = io_x[88] ? _GEN1333 : _GEN1332;
wire  _GEN1335 = 1'b1;
wire  _GEN1336 = io_x[89] ? _GEN1335 : _GEN1334;
wire  _GEN1337 = 1'b1;
wire  _GEN1338 = io_x[90] ? _GEN1337 : _GEN1336;
wire  _GEN1339 = 1'b1;
wire  _GEN1340 = io_x[91] ? _GEN1339 : _GEN1338;
wire  _GEN1341 = 1'b1;
wire  _GEN1342 = io_x[92] ? _GEN1341 : _GEN1340;
wire  _GEN1343 = 1'b1;
wire  _GEN1344 = io_x[93] ? _GEN1343 : _GEN1342;
wire  _GEN1345 = 1'b1;
wire  _GEN1346 = io_x[94] ? _GEN1345 : _GEN1344;
wire  _GEN1347 = 1'b1;
wire  _GEN1348 = io_x[95] ? _GEN1347 : _GEN1346;
wire  _GEN1349 = 1'b1;
wire  _GEN1350 = io_x[96] ? _GEN1349 : _GEN1348;
wire  _GEN1351 = 1'b1;
wire  _GEN1352 = io_x[97] ? _GEN1351 : _GEN1350;
wire  _GEN1353 = io_x[98] ? _GEN1352 : _GEN0;
wire  _GEN1354 = 1'b1;
wire  _GEN1355 = io_x[33] ? _GEN1354 : _GEN1353;
wire  _GEN1356 = 1'b0;
wire  _GEN1357 = io_x[33] ? _GEN1354 : _GEN1356;
wire  _GEN1358 = io_x[32] ? _GEN1357 : _GEN1355;
assign io_y[20] = _GEN1358;
wire  _GEN1359 = 1'b0;
wire  _GEN1360 = 1'b1;
wire  _GEN1361 = io_x[34] ? _GEN1360 : _GEN1359;
wire  _GEN1362 = io_x[34] ? _GEN1360 : _GEN1359;
wire  _GEN1363 = io_x[38] ? _GEN1362 : _GEN1361;
wire  _GEN1364 = io_x[34] ? _GEN1360 : _GEN1359;
wire  _GEN1365 = io_x[34] ? _GEN1360 : _GEN1359;
wire  _GEN1366 = io_x[38] ? _GEN1365 : _GEN1364;
wire  _GEN1367 = io_x[44] ? _GEN1366 : _GEN1363;
wire  _GEN1368 = io_x[34] ? _GEN1360 : _GEN1359;
wire  _GEN1369 = io_x[34] ? _GEN1360 : _GEN1359;
wire  _GEN1370 = io_x[38] ? _GEN1369 : _GEN1368;
wire  _GEN1371 = io_x[34] ? _GEN1360 : _GEN1359;
wire  _GEN1372 = io_x[34] ? _GEN1360 : _GEN1359;
wire  _GEN1373 = io_x[38] ? _GEN1372 : _GEN1371;
wire  _GEN1374 = io_x[44] ? _GEN1373 : _GEN1370;
wire  _GEN1375 = io_x[4] ? _GEN1374 : _GEN1367;
assign io_y[19] = _GEN1375;
wire  _GEN1376 = 1'b0;
wire  _GEN1377 = 1'b1;
wire  _GEN1378 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1379 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1380 = io_x[23] ? _GEN1379 : _GEN1378;
wire  _GEN1381 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1382 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1383 = io_x[23] ? _GEN1382 : _GEN1381;
wire  _GEN1384 = io_x[19] ? _GEN1383 : _GEN1380;
wire  _GEN1385 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1386 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1387 = io_x[23] ? _GEN1386 : _GEN1385;
wire  _GEN1388 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1389 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1390 = io_x[23] ? _GEN1389 : _GEN1388;
wire  _GEN1391 = io_x[19] ? _GEN1390 : _GEN1387;
wire  _GEN1392 = io_x[31] ? _GEN1391 : _GEN1384;
wire  _GEN1393 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1394 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1395 = io_x[23] ? _GEN1394 : _GEN1393;
wire  _GEN1396 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1397 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1398 = io_x[23] ? _GEN1397 : _GEN1396;
wire  _GEN1399 = io_x[19] ? _GEN1398 : _GEN1395;
wire  _GEN1400 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1401 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1402 = io_x[23] ? _GEN1401 : _GEN1400;
wire  _GEN1403 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1404 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1405 = io_x[23] ? _GEN1404 : _GEN1403;
wire  _GEN1406 = io_x[19] ? _GEN1405 : _GEN1402;
wire  _GEN1407 = io_x[31] ? _GEN1406 : _GEN1399;
wire  _GEN1408 = io_x[27] ? _GEN1407 : _GEN1392;
wire  _GEN1409 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1410 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1411 = io_x[23] ? _GEN1410 : _GEN1409;
wire  _GEN1412 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1413 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1414 = io_x[23] ? _GEN1413 : _GEN1412;
wire  _GEN1415 = io_x[19] ? _GEN1414 : _GEN1411;
wire  _GEN1416 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1417 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1418 = io_x[23] ? _GEN1417 : _GEN1416;
wire  _GEN1419 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1420 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1421 = io_x[23] ? _GEN1420 : _GEN1419;
wire  _GEN1422 = io_x[19] ? _GEN1421 : _GEN1418;
wire  _GEN1423 = io_x[31] ? _GEN1422 : _GEN1415;
wire  _GEN1424 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1425 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1426 = io_x[23] ? _GEN1425 : _GEN1424;
wire  _GEN1427 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1428 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1429 = io_x[23] ? _GEN1428 : _GEN1427;
wire  _GEN1430 = io_x[19] ? _GEN1429 : _GEN1426;
wire  _GEN1431 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1432 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1433 = io_x[23] ? _GEN1432 : _GEN1431;
wire  _GEN1434 = io_x[77] ? _GEN1376 : _GEN1377;
wire  _GEN1435 = io_x[77] ? _GEN1377 : _GEN1376;
wire  _GEN1436 = io_x[23] ? _GEN1435 : _GEN1434;
wire  _GEN1437 = io_x[19] ? _GEN1436 : _GEN1433;
wire  _GEN1438 = io_x[31] ? _GEN1437 : _GEN1430;
wire  _GEN1439 = io_x[27] ? _GEN1438 : _GEN1423;
wire  _GEN1440 = io_x[45] ? _GEN1439 : _GEN1408;
assign io_y[18] = _GEN1440;
wire  _GEN1441 = 1'b0;
wire  _GEN1442 = 1'b1;
wire  _GEN1443 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1444 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1445 = io_x[22] ? _GEN1444 : _GEN1443;
wire  _GEN1446 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1447 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1448 = io_x[22] ? _GEN1447 : _GEN1446;
wire  _GEN1449 = io_x[18] ? _GEN1448 : _GEN1445;
wire  _GEN1450 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1451 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1452 = io_x[22] ? _GEN1451 : _GEN1450;
wire  _GEN1453 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1454 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1455 = io_x[22] ? _GEN1454 : _GEN1453;
wire  _GEN1456 = io_x[18] ? _GEN1455 : _GEN1452;
wire  _GEN1457 = io_x[75] ? _GEN1456 : _GEN1449;
wire  _GEN1458 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1459 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1460 = io_x[22] ? _GEN1459 : _GEN1458;
wire  _GEN1461 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1462 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1463 = io_x[22] ? _GEN1462 : _GEN1461;
wire  _GEN1464 = io_x[18] ? _GEN1463 : _GEN1460;
wire  _GEN1465 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1466 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1467 = io_x[22] ? _GEN1466 : _GEN1465;
wire  _GEN1468 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1469 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1470 = io_x[22] ? _GEN1469 : _GEN1468;
wire  _GEN1471 = io_x[18] ? _GEN1470 : _GEN1467;
wire  _GEN1472 = io_x[75] ? _GEN1471 : _GEN1464;
wire  _GEN1473 = io_x[30] ? _GEN1472 : _GEN1457;
wire  _GEN1474 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1475 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1476 = io_x[22] ? _GEN1475 : _GEN1474;
wire  _GEN1477 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1478 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1479 = io_x[22] ? _GEN1478 : _GEN1477;
wire  _GEN1480 = io_x[18] ? _GEN1479 : _GEN1476;
wire  _GEN1481 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1482 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1483 = io_x[22] ? _GEN1482 : _GEN1481;
wire  _GEN1484 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1485 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1486 = io_x[22] ? _GEN1485 : _GEN1484;
wire  _GEN1487 = io_x[18] ? _GEN1486 : _GEN1483;
wire  _GEN1488 = io_x[75] ? _GEN1487 : _GEN1480;
wire  _GEN1489 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1490 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1491 = io_x[22] ? _GEN1490 : _GEN1489;
wire  _GEN1492 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1493 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1494 = io_x[22] ? _GEN1493 : _GEN1492;
wire  _GEN1495 = io_x[18] ? _GEN1494 : _GEN1491;
wire  _GEN1496 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1497 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1498 = io_x[22] ? _GEN1497 : _GEN1496;
wire  _GEN1499 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1500 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1501 = io_x[22] ? _GEN1500 : _GEN1499;
wire  _GEN1502 = io_x[18] ? _GEN1501 : _GEN1498;
wire  _GEN1503 = io_x[75] ? _GEN1502 : _GEN1495;
wire  _GEN1504 = io_x[30] ? _GEN1503 : _GEN1488;
wire  _GEN1505 = io_x[26] ? _GEN1504 : _GEN1473;
wire  _GEN1506 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1507 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1508 = io_x[22] ? _GEN1507 : _GEN1506;
wire  _GEN1509 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1510 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1511 = io_x[22] ? _GEN1510 : _GEN1509;
wire  _GEN1512 = io_x[18] ? _GEN1511 : _GEN1508;
wire  _GEN1513 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1514 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1515 = io_x[22] ? _GEN1514 : _GEN1513;
wire  _GEN1516 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1517 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1518 = io_x[22] ? _GEN1517 : _GEN1516;
wire  _GEN1519 = io_x[18] ? _GEN1518 : _GEN1515;
wire  _GEN1520 = io_x[75] ? _GEN1519 : _GEN1512;
wire  _GEN1521 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1522 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1523 = io_x[22] ? _GEN1522 : _GEN1521;
wire  _GEN1524 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1525 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1526 = io_x[22] ? _GEN1525 : _GEN1524;
wire  _GEN1527 = io_x[18] ? _GEN1526 : _GEN1523;
wire  _GEN1528 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1529 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1530 = io_x[22] ? _GEN1529 : _GEN1528;
wire  _GEN1531 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1532 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1533 = io_x[22] ? _GEN1532 : _GEN1531;
wire  _GEN1534 = io_x[18] ? _GEN1533 : _GEN1530;
wire  _GEN1535 = io_x[75] ? _GEN1534 : _GEN1527;
wire  _GEN1536 = io_x[30] ? _GEN1535 : _GEN1520;
wire  _GEN1537 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1538 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1539 = io_x[22] ? _GEN1538 : _GEN1537;
wire  _GEN1540 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1541 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1542 = io_x[22] ? _GEN1541 : _GEN1540;
wire  _GEN1543 = io_x[18] ? _GEN1542 : _GEN1539;
wire  _GEN1544 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1545 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1546 = io_x[22] ? _GEN1545 : _GEN1544;
wire  _GEN1547 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1548 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1549 = io_x[22] ? _GEN1548 : _GEN1547;
wire  _GEN1550 = io_x[18] ? _GEN1549 : _GEN1546;
wire  _GEN1551 = io_x[75] ? _GEN1550 : _GEN1543;
wire  _GEN1552 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1553 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1554 = io_x[22] ? _GEN1553 : _GEN1552;
wire  _GEN1555 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1556 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1557 = io_x[22] ? _GEN1556 : _GEN1555;
wire  _GEN1558 = io_x[18] ? _GEN1557 : _GEN1554;
wire  _GEN1559 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1560 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1561 = io_x[22] ? _GEN1560 : _GEN1559;
wire  _GEN1562 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1563 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1564 = io_x[22] ? _GEN1563 : _GEN1562;
wire  _GEN1565 = io_x[18] ? _GEN1564 : _GEN1561;
wire  _GEN1566 = io_x[75] ? _GEN1565 : _GEN1558;
wire  _GEN1567 = io_x[30] ? _GEN1566 : _GEN1551;
wire  _GEN1568 = io_x[26] ? _GEN1567 : _GEN1536;
wire  _GEN1569 = io_x[73] ? _GEN1568 : _GEN1505;
wire  _GEN1570 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1571 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1572 = io_x[22] ? _GEN1571 : _GEN1570;
wire  _GEN1573 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1574 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1575 = io_x[22] ? _GEN1574 : _GEN1573;
wire  _GEN1576 = io_x[18] ? _GEN1575 : _GEN1572;
wire  _GEN1577 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1578 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1579 = io_x[22] ? _GEN1578 : _GEN1577;
wire  _GEN1580 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1581 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1582 = io_x[22] ? _GEN1581 : _GEN1580;
wire  _GEN1583 = io_x[18] ? _GEN1582 : _GEN1579;
wire  _GEN1584 = io_x[75] ? _GEN1583 : _GEN1576;
wire  _GEN1585 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1586 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1587 = io_x[22] ? _GEN1586 : _GEN1585;
wire  _GEN1588 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1589 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1590 = io_x[22] ? _GEN1589 : _GEN1588;
wire  _GEN1591 = io_x[18] ? _GEN1590 : _GEN1587;
wire  _GEN1592 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1593 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1594 = io_x[22] ? _GEN1593 : _GEN1592;
wire  _GEN1595 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1596 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1597 = io_x[22] ? _GEN1596 : _GEN1595;
wire  _GEN1598 = io_x[18] ? _GEN1597 : _GEN1594;
wire  _GEN1599 = io_x[75] ? _GEN1598 : _GEN1591;
wire  _GEN1600 = io_x[30] ? _GEN1599 : _GEN1584;
wire  _GEN1601 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1602 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1603 = io_x[22] ? _GEN1602 : _GEN1601;
wire  _GEN1604 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1605 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1606 = io_x[22] ? _GEN1605 : _GEN1604;
wire  _GEN1607 = io_x[18] ? _GEN1606 : _GEN1603;
wire  _GEN1608 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1609 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1610 = io_x[22] ? _GEN1609 : _GEN1608;
wire  _GEN1611 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1612 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1613 = io_x[22] ? _GEN1612 : _GEN1611;
wire  _GEN1614 = io_x[18] ? _GEN1613 : _GEN1610;
wire  _GEN1615 = io_x[75] ? _GEN1614 : _GEN1607;
wire  _GEN1616 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1617 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1618 = io_x[22] ? _GEN1617 : _GEN1616;
wire  _GEN1619 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1620 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1621 = io_x[22] ? _GEN1620 : _GEN1619;
wire  _GEN1622 = io_x[18] ? _GEN1621 : _GEN1618;
wire  _GEN1623 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1624 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1625 = io_x[22] ? _GEN1624 : _GEN1623;
wire  _GEN1626 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1627 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1628 = io_x[22] ? _GEN1627 : _GEN1626;
wire  _GEN1629 = io_x[18] ? _GEN1628 : _GEN1625;
wire  _GEN1630 = io_x[75] ? _GEN1629 : _GEN1622;
wire  _GEN1631 = io_x[30] ? _GEN1630 : _GEN1615;
wire  _GEN1632 = io_x[26] ? _GEN1631 : _GEN1600;
wire  _GEN1633 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1634 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1635 = io_x[22] ? _GEN1634 : _GEN1633;
wire  _GEN1636 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1637 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1638 = io_x[22] ? _GEN1637 : _GEN1636;
wire  _GEN1639 = io_x[18] ? _GEN1638 : _GEN1635;
wire  _GEN1640 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1641 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1642 = io_x[22] ? _GEN1641 : _GEN1640;
wire  _GEN1643 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1644 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1645 = io_x[22] ? _GEN1644 : _GEN1643;
wire  _GEN1646 = io_x[18] ? _GEN1645 : _GEN1642;
wire  _GEN1647 = io_x[75] ? _GEN1646 : _GEN1639;
wire  _GEN1648 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1649 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1650 = io_x[22] ? _GEN1649 : _GEN1648;
wire  _GEN1651 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1652 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1653 = io_x[22] ? _GEN1652 : _GEN1651;
wire  _GEN1654 = io_x[18] ? _GEN1653 : _GEN1650;
wire  _GEN1655 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1656 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1657 = io_x[22] ? _GEN1656 : _GEN1655;
wire  _GEN1658 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1659 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1660 = io_x[22] ? _GEN1659 : _GEN1658;
wire  _GEN1661 = io_x[18] ? _GEN1660 : _GEN1657;
wire  _GEN1662 = io_x[75] ? _GEN1661 : _GEN1654;
wire  _GEN1663 = io_x[30] ? _GEN1662 : _GEN1647;
wire  _GEN1664 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1665 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1666 = io_x[22] ? _GEN1665 : _GEN1664;
wire  _GEN1667 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1668 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1669 = io_x[22] ? _GEN1668 : _GEN1667;
wire  _GEN1670 = io_x[18] ? _GEN1669 : _GEN1666;
wire  _GEN1671 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1672 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1673 = io_x[22] ? _GEN1672 : _GEN1671;
wire  _GEN1674 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1675 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1676 = io_x[22] ? _GEN1675 : _GEN1674;
wire  _GEN1677 = io_x[18] ? _GEN1676 : _GEN1673;
wire  _GEN1678 = io_x[75] ? _GEN1677 : _GEN1670;
wire  _GEN1679 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1680 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1681 = io_x[22] ? _GEN1680 : _GEN1679;
wire  _GEN1682 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1683 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1684 = io_x[22] ? _GEN1683 : _GEN1682;
wire  _GEN1685 = io_x[18] ? _GEN1684 : _GEN1681;
wire  _GEN1686 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1687 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1688 = io_x[22] ? _GEN1687 : _GEN1686;
wire  _GEN1689 = io_x[76] ? _GEN1441 : _GEN1442;
wire  _GEN1690 = io_x[76] ? _GEN1442 : _GEN1441;
wire  _GEN1691 = io_x[22] ? _GEN1690 : _GEN1689;
wire  _GEN1692 = io_x[18] ? _GEN1691 : _GEN1688;
wire  _GEN1693 = io_x[75] ? _GEN1692 : _GEN1685;
wire  _GEN1694 = io_x[30] ? _GEN1693 : _GEN1678;
wire  _GEN1695 = io_x[26] ? _GEN1694 : _GEN1663;
wire  _GEN1696 = io_x[73] ? _GEN1695 : _GEN1632;
wire  _GEN1697 = io_x[38] ? _GEN1696 : _GEN1569;
assign io_y[17] = _GEN1697;
wire  _GEN1698 = 1'b0;
wire  _GEN1699 = 1'b1;
wire  _GEN1700 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1701 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1702 = io_x[17] ? _GEN1701 : _GEN1700;
wire  _GEN1703 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1704 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1705 = io_x[17] ? _GEN1704 : _GEN1703;
wire  _GEN1706 = io_x[75] ? _GEN1705 : _GEN1702;
wire  _GEN1707 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1708 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1709 = io_x[17] ? _GEN1708 : _GEN1707;
wire  _GEN1710 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1711 = 1'b0;
wire  _GEN1712 = io_x[17] ? _GEN1711 : _GEN1710;
wire  _GEN1713 = io_x[75] ? _GEN1712 : _GEN1709;
wire  _GEN1714 = io_x[25] ? _GEN1713 : _GEN1706;
wire  _GEN1715 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1716 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1717 = io_x[17] ? _GEN1716 : _GEN1715;
wire  _GEN1718 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1719 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1720 = io_x[17] ? _GEN1719 : _GEN1718;
wire  _GEN1721 = io_x[75] ? _GEN1720 : _GEN1717;
wire  _GEN1722 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1723 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1724 = io_x[17] ? _GEN1723 : _GEN1722;
wire  _GEN1725 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1726 = io_x[17] ? _GEN1711 : _GEN1725;
wire  _GEN1727 = io_x[75] ? _GEN1726 : _GEN1724;
wire  _GEN1728 = io_x[25] ? _GEN1727 : _GEN1721;
wire  _GEN1729 = io_x[37] ? _GEN1728 : _GEN1714;
wire  _GEN1730 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1731 = 1'b1;
wire  _GEN1732 = io_x[17] ? _GEN1731 : _GEN1730;
wire  _GEN1733 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1734 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1735 = io_x[17] ? _GEN1734 : _GEN1733;
wire  _GEN1736 = io_x[75] ? _GEN1735 : _GEN1732;
wire  _GEN1737 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN1738 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1739 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1740 = io_x[17] ? _GEN1739 : _GEN1738;
wire  _GEN1741 = io_x[75] ? _GEN1740 : _GEN1737;
wire  _GEN1742 = io_x[25] ? _GEN1741 : _GEN1736;
wire  _GEN1743 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1744 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1745 = io_x[17] ? _GEN1744 : _GEN1743;
wire  _GEN1746 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1747 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1748 = io_x[17] ? _GEN1747 : _GEN1746;
wire  _GEN1749 = io_x[75] ? _GEN1748 : _GEN1745;
wire  _GEN1750 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1751 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1752 = io_x[17] ? _GEN1751 : _GEN1750;
wire  _GEN1753 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1754 = io_x[17] ? _GEN1731 : _GEN1753;
wire  _GEN1755 = io_x[75] ? _GEN1754 : _GEN1752;
wire  _GEN1756 = io_x[25] ? _GEN1755 : _GEN1749;
wire  _GEN1757 = io_x[37] ? _GEN1756 : _GEN1742;
wire  _GEN1758 = io_x[39] ? _GEN1757 : _GEN1729;
wire  _GEN1759 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1760 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1761 = io_x[17] ? _GEN1760 : _GEN1759;
wire  _GEN1762 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1763 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1764 = io_x[17] ? _GEN1763 : _GEN1762;
wire  _GEN1765 = io_x[75] ? _GEN1764 : _GEN1761;
wire  _GEN1766 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1767 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1768 = io_x[17] ? _GEN1767 : _GEN1766;
wire  _GEN1769 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1770 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1771 = io_x[17] ? _GEN1770 : _GEN1769;
wire  _GEN1772 = io_x[75] ? _GEN1771 : _GEN1768;
wire  _GEN1773 = io_x[25] ? _GEN1772 : _GEN1765;
wire  _GEN1774 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1775 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1776 = io_x[17] ? _GEN1775 : _GEN1774;
wire  _GEN1777 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1778 = io_x[17] ? _GEN1711 : _GEN1777;
wire  _GEN1779 = io_x[75] ? _GEN1778 : _GEN1776;
wire  _GEN1780 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1781 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1782 = io_x[17] ? _GEN1781 : _GEN1780;
wire  _GEN1783 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1784 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1785 = io_x[17] ? _GEN1784 : _GEN1783;
wire  _GEN1786 = io_x[75] ? _GEN1785 : _GEN1782;
wire  _GEN1787 = io_x[25] ? _GEN1786 : _GEN1779;
wire  _GEN1788 = io_x[37] ? _GEN1787 : _GEN1773;
wire  _GEN1789 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1790 = io_x[17] ? _GEN1731 : _GEN1789;
wire  _GEN1791 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1792 = io_x[17] ? _GEN1711 : _GEN1791;
wire  _GEN1793 = io_x[75] ? _GEN1792 : _GEN1790;
wire  _GEN1794 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN1795 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1796 = io_x[17] ? _GEN1795 : _GEN1731;
wire  _GEN1797 = io_x[75] ? _GEN1796 : _GEN1794;
wire  _GEN1798 = io_x[25] ? _GEN1797 : _GEN1793;
wire  _GEN1799 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1800 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1801 = io_x[17] ? _GEN1800 : _GEN1799;
wire  _GEN1802 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1803 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1804 = io_x[17] ? _GEN1803 : _GEN1802;
wire  _GEN1805 = io_x[75] ? _GEN1804 : _GEN1801;
wire  _GEN1806 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1807 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1808 = io_x[17] ? _GEN1807 : _GEN1806;
wire  _GEN1809 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1810 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1811 = io_x[17] ? _GEN1810 : _GEN1809;
wire  _GEN1812 = io_x[75] ? _GEN1811 : _GEN1808;
wire  _GEN1813 = io_x[25] ? _GEN1812 : _GEN1805;
wire  _GEN1814 = io_x[37] ? _GEN1813 : _GEN1798;
wire  _GEN1815 = io_x[39] ? _GEN1814 : _GEN1788;
wire  _GEN1816 = io_x[72] ? _GEN1815 : _GEN1758;
wire  _GEN1817 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1818 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1819 = io_x[17] ? _GEN1818 : _GEN1817;
wire  _GEN1820 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1821 = io_x[17] ? _GEN1711 : _GEN1820;
wire  _GEN1822 = io_x[75] ? _GEN1821 : _GEN1819;
wire  _GEN1823 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1824 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1825 = io_x[17] ? _GEN1824 : _GEN1823;
wire  _GEN1826 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1827 = io_x[17] ? _GEN1731 : _GEN1826;
wire  _GEN1828 = io_x[75] ? _GEN1827 : _GEN1825;
wire  _GEN1829 = io_x[25] ? _GEN1828 : _GEN1822;
wire  _GEN1830 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1831 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1832 = io_x[17] ? _GEN1831 : _GEN1830;
wire  _GEN1833 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1834 = io_x[17] ? _GEN1731 : _GEN1833;
wire  _GEN1835 = io_x[75] ? _GEN1834 : _GEN1832;
wire  _GEN1836 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1837 = io_x[17] ? _GEN1836 : _GEN1711;
wire  _GEN1838 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1839 = io_x[17] ? _GEN1731 : _GEN1838;
wire  _GEN1840 = io_x[75] ? _GEN1839 : _GEN1837;
wire  _GEN1841 = io_x[25] ? _GEN1840 : _GEN1835;
wire  _GEN1842 = io_x[37] ? _GEN1841 : _GEN1829;
wire  _GEN1843 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1844 = io_x[17] ? _GEN1711 : _GEN1843;
wire  _GEN1845 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1846 = io_x[17] ? _GEN1731 : _GEN1845;
wire  _GEN1847 = io_x[75] ? _GEN1846 : _GEN1844;
wire  _GEN1848 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN1849 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1850 = io_x[17] ? _GEN1731 : _GEN1849;
wire  _GEN1851 = io_x[75] ? _GEN1850 : _GEN1848;
wire  _GEN1852 = io_x[25] ? _GEN1851 : _GEN1847;
wire  _GEN1853 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1854 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1855 = io_x[17] ? _GEN1854 : _GEN1853;
wire  _GEN1856 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1857 = io_x[17] ? _GEN1731 : _GEN1856;
wire  _GEN1858 = io_x[75] ? _GEN1857 : _GEN1855;
wire  _GEN1859 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1860 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1861 = io_x[17] ? _GEN1860 : _GEN1859;
wire  _GEN1862 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1863 = io_x[17] ? _GEN1731 : _GEN1862;
wire  _GEN1864 = io_x[75] ? _GEN1863 : _GEN1861;
wire  _GEN1865 = io_x[25] ? _GEN1864 : _GEN1858;
wire  _GEN1866 = io_x[37] ? _GEN1865 : _GEN1852;
wire  _GEN1867 = io_x[39] ? _GEN1866 : _GEN1842;
wire  _GEN1868 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1869 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1870 = io_x[17] ? _GEN1869 : _GEN1868;
wire  _GEN1871 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1872 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1873 = io_x[17] ? _GEN1872 : _GEN1871;
wire  _GEN1874 = io_x[75] ? _GEN1873 : _GEN1870;
wire  _GEN1875 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1876 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1877 = io_x[17] ? _GEN1876 : _GEN1875;
wire  _GEN1878 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1879 = io_x[17] ? _GEN1731 : _GEN1878;
wire  _GEN1880 = io_x[75] ? _GEN1879 : _GEN1877;
wire  _GEN1881 = io_x[25] ? _GEN1880 : _GEN1874;
wire  _GEN1882 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1883 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1884 = io_x[17] ? _GEN1883 : _GEN1882;
wire  _GEN1885 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1886 = io_x[17] ? _GEN1711 : _GEN1885;
wire  _GEN1887 = io_x[75] ? _GEN1886 : _GEN1884;
wire  _GEN1888 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1889 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1890 = io_x[17] ? _GEN1889 : _GEN1888;
wire  _GEN1891 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1892 = io_x[17] ? _GEN1711 : _GEN1891;
wire  _GEN1893 = io_x[75] ? _GEN1892 : _GEN1890;
wire  _GEN1894 = io_x[25] ? _GEN1893 : _GEN1887;
wire  _GEN1895 = io_x[37] ? _GEN1894 : _GEN1881;
wire  _GEN1896 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1897 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1898 = io_x[17] ? _GEN1897 : _GEN1896;
wire  _GEN1899 = 1'b1;
wire  _GEN1900 = io_x[75] ? _GEN1899 : _GEN1898;
wire  _GEN1901 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1902 = io_x[17] ? _GEN1731 : _GEN1901;
wire  _GEN1903 = 1'b0;
wire  _GEN1904 = io_x[75] ? _GEN1903 : _GEN1902;
wire  _GEN1905 = io_x[25] ? _GEN1904 : _GEN1900;
wire  _GEN1906 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1907 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1908 = io_x[17] ? _GEN1907 : _GEN1906;
wire  _GEN1909 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1910 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1911 = io_x[17] ? _GEN1910 : _GEN1909;
wire  _GEN1912 = io_x[75] ? _GEN1911 : _GEN1908;
wire  _GEN1913 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1914 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1915 = io_x[17] ? _GEN1914 : _GEN1913;
wire  _GEN1916 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1917 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1918 = io_x[17] ? _GEN1917 : _GEN1916;
wire  _GEN1919 = io_x[75] ? _GEN1918 : _GEN1915;
wire  _GEN1920 = io_x[25] ? _GEN1919 : _GEN1912;
wire  _GEN1921 = io_x[37] ? _GEN1920 : _GEN1905;
wire  _GEN1922 = io_x[39] ? _GEN1921 : _GEN1895;
wire  _GEN1923 = io_x[72] ? _GEN1922 : _GEN1867;
wire  _GEN1924 = io_x[29] ? _GEN1923 : _GEN1816;
wire  _GEN1925 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1926 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1927 = io_x[17] ? _GEN1926 : _GEN1925;
wire  _GEN1928 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1929 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1930 = io_x[17] ? _GEN1929 : _GEN1928;
wire  _GEN1931 = io_x[75] ? _GEN1930 : _GEN1927;
wire  _GEN1932 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1933 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1934 = io_x[17] ? _GEN1933 : _GEN1932;
wire  _GEN1935 = io_x[75] ? _GEN1899 : _GEN1934;
wire  _GEN1936 = io_x[25] ? _GEN1935 : _GEN1931;
wire  _GEN1937 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1938 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1939 = io_x[17] ? _GEN1938 : _GEN1937;
wire  _GEN1940 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1941 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1942 = io_x[17] ? _GEN1941 : _GEN1940;
wire  _GEN1943 = io_x[75] ? _GEN1942 : _GEN1939;
wire  _GEN1944 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1945 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1946 = io_x[17] ? _GEN1945 : _GEN1944;
wire  _GEN1947 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN1948 = io_x[75] ? _GEN1947 : _GEN1946;
wire  _GEN1949 = io_x[25] ? _GEN1948 : _GEN1943;
wire  _GEN1950 = io_x[37] ? _GEN1949 : _GEN1936;
wire  _GEN1951 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1952 = io_x[17] ? _GEN1951 : _GEN1711;
wire  _GEN1953 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1954 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1955 = io_x[17] ? _GEN1954 : _GEN1953;
wire  _GEN1956 = io_x[75] ? _GEN1955 : _GEN1952;
wire  _GEN1957 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1958 = io_x[17] ? _GEN1731 : _GEN1957;
wire  _GEN1959 = io_x[75] ? _GEN1958 : _GEN1903;
wire  _GEN1960 = io_x[25] ? _GEN1959 : _GEN1956;
wire  _GEN1961 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1962 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1963 = io_x[17] ? _GEN1962 : _GEN1961;
wire  _GEN1964 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1965 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1966 = io_x[17] ? _GEN1965 : _GEN1964;
wire  _GEN1967 = io_x[75] ? _GEN1966 : _GEN1963;
wire  _GEN1968 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1969 = io_x[17] ? _GEN1711 : _GEN1968;
wire  _GEN1970 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1971 = io_x[17] ? _GEN1970 : _GEN1711;
wire  _GEN1972 = io_x[75] ? _GEN1971 : _GEN1969;
wire  _GEN1973 = io_x[25] ? _GEN1972 : _GEN1967;
wire  _GEN1974 = io_x[37] ? _GEN1973 : _GEN1960;
wire  _GEN1975 = io_x[39] ? _GEN1974 : _GEN1950;
wire  _GEN1976 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1977 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1978 = io_x[17] ? _GEN1977 : _GEN1976;
wire  _GEN1979 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1980 = io_x[17] ? _GEN1979 : _GEN1731;
wire  _GEN1981 = io_x[75] ? _GEN1980 : _GEN1978;
wire  _GEN1982 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1983 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1984 = io_x[17] ? _GEN1983 : _GEN1982;
wire  _GEN1985 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1986 = io_x[17] ? _GEN1985 : _GEN1731;
wire  _GEN1987 = io_x[75] ? _GEN1986 : _GEN1984;
wire  _GEN1988 = io_x[25] ? _GEN1987 : _GEN1981;
wire  _GEN1989 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1990 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1991 = io_x[17] ? _GEN1990 : _GEN1989;
wire  _GEN1992 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1993 = io_x[17] ? _GEN1992 : _GEN1731;
wire  _GEN1994 = io_x[75] ? _GEN1993 : _GEN1991;
wire  _GEN1995 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN1996 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN1997 = io_x[17] ? _GEN1996 : _GEN1995;
wire  _GEN1998 = io_x[75] ? _GEN1899 : _GEN1997;
wire  _GEN1999 = io_x[25] ? _GEN1998 : _GEN1994;
wire  _GEN2000 = io_x[37] ? _GEN1999 : _GEN1988;
wire  _GEN2001 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2002 = io_x[17] ? _GEN2001 : _GEN1711;
wire  _GEN2003 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2004 = io_x[17] ? _GEN2003 : _GEN1731;
wire  _GEN2005 = io_x[75] ? _GEN2004 : _GEN2002;
wire  _GEN2006 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2007 = io_x[17] ? _GEN2006 : _GEN1731;
wire  _GEN2008 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2009 = io_x[17] ? _GEN2008 : _GEN1731;
wire  _GEN2010 = io_x[75] ? _GEN2009 : _GEN2007;
wire  _GEN2011 = io_x[25] ? _GEN2010 : _GEN2005;
wire  _GEN2012 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2013 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2014 = io_x[17] ? _GEN2013 : _GEN2012;
wire  _GEN2015 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2016 = io_x[17] ? _GEN1711 : _GEN2015;
wire  _GEN2017 = io_x[75] ? _GEN2016 : _GEN2014;
wire  _GEN2018 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2019 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2020 = io_x[17] ? _GEN2019 : _GEN2018;
wire  _GEN2021 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2022 = io_x[17] ? _GEN1731 : _GEN2021;
wire  _GEN2023 = io_x[75] ? _GEN2022 : _GEN2020;
wire  _GEN2024 = io_x[25] ? _GEN2023 : _GEN2017;
wire  _GEN2025 = io_x[37] ? _GEN2024 : _GEN2011;
wire  _GEN2026 = io_x[39] ? _GEN2025 : _GEN2000;
wire  _GEN2027 = io_x[72] ? _GEN2026 : _GEN1975;
wire  _GEN2028 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2029 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2030 = io_x[17] ? _GEN2029 : _GEN2028;
wire  _GEN2031 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2032 = io_x[17] ? _GEN2031 : _GEN1731;
wire  _GEN2033 = io_x[75] ? _GEN2032 : _GEN2030;
wire  _GEN2034 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2035 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2036 = io_x[17] ? _GEN2035 : _GEN2034;
wire  _GEN2037 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2038 = io_x[17] ? _GEN2037 : _GEN1731;
wire  _GEN2039 = io_x[75] ? _GEN2038 : _GEN2036;
wire  _GEN2040 = io_x[25] ? _GEN2039 : _GEN2033;
wire  _GEN2041 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2042 = io_x[17] ? _GEN2041 : _GEN1711;
wire  _GEN2043 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2044 = io_x[17] ? _GEN1731 : _GEN2043;
wire  _GEN2045 = io_x[75] ? _GEN2044 : _GEN2042;
wire  _GEN2046 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN2047 = io_x[75] ? _GEN1899 : _GEN2046;
wire  _GEN2048 = io_x[25] ? _GEN2047 : _GEN2045;
wire  _GEN2049 = io_x[37] ? _GEN2048 : _GEN2040;
wire  _GEN2050 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2051 = io_x[17] ? _GEN2050 : _GEN1731;
wire  _GEN2052 = io_x[75] ? _GEN1899 : _GEN2051;
wire  _GEN2053 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2054 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2055 = io_x[17] ? _GEN2054 : _GEN2053;
wire  _GEN2056 = io_x[75] ? _GEN1899 : _GEN2055;
wire  _GEN2057 = io_x[25] ? _GEN2056 : _GEN2052;
wire  _GEN2058 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2059 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2060 = io_x[17] ? _GEN2059 : _GEN2058;
wire  _GEN2061 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2062 = io_x[17] ? _GEN1711 : _GEN2061;
wire  _GEN2063 = io_x[75] ? _GEN2062 : _GEN2060;
wire  _GEN2064 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2065 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2066 = io_x[17] ? _GEN2065 : _GEN2064;
wire  _GEN2067 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2068 = io_x[17] ? _GEN2067 : _GEN1731;
wire  _GEN2069 = io_x[75] ? _GEN2068 : _GEN2066;
wire  _GEN2070 = io_x[25] ? _GEN2069 : _GEN2063;
wire  _GEN2071 = io_x[37] ? _GEN2070 : _GEN2057;
wire  _GEN2072 = io_x[39] ? _GEN2071 : _GEN2049;
wire  _GEN2073 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2074 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2075 = io_x[17] ? _GEN2074 : _GEN2073;
wire  _GEN2076 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN2077 = io_x[75] ? _GEN2076 : _GEN2075;
wire  _GEN2078 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2079 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2080 = io_x[17] ? _GEN2079 : _GEN2078;
wire  _GEN2081 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2082 = io_x[17] ? _GEN2081 : _GEN1731;
wire  _GEN2083 = io_x[75] ? _GEN2082 : _GEN2080;
wire  _GEN2084 = io_x[25] ? _GEN2083 : _GEN2077;
wire  _GEN2085 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2086 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2087 = io_x[17] ? _GEN2086 : _GEN2085;
wire  _GEN2088 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2089 = io_x[17] ? _GEN2088 : _GEN1731;
wire  _GEN2090 = io_x[75] ? _GEN2089 : _GEN2087;
wire  _GEN2091 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2092 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2093 = io_x[17] ? _GEN2092 : _GEN2091;
wire  _GEN2094 = io_x[75] ? _GEN1903 : _GEN2093;
wire  _GEN2095 = io_x[25] ? _GEN2094 : _GEN2090;
wire  _GEN2096 = io_x[37] ? _GEN2095 : _GEN2084;
wire  _GEN2097 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2098 = io_x[17] ? _GEN2097 : _GEN1711;
wire  _GEN2099 = io_x[75] ? _GEN1903 : _GEN2098;
wire  _GEN2100 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2101 = io_x[17] ? _GEN2100 : _GEN1731;
wire  _GEN2102 = io_x[75] ? _GEN1899 : _GEN2101;
wire  _GEN2103 = io_x[25] ? _GEN2102 : _GEN2099;
wire  _GEN2104 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2105 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2106 = io_x[17] ? _GEN2105 : _GEN2104;
wire  _GEN2107 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2108 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2109 = io_x[17] ? _GEN2108 : _GEN2107;
wire  _GEN2110 = io_x[75] ? _GEN2109 : _GEN2106;
wire  _GEN2111 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2112 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2113 = io_x[17] ? _GEN2112 : _GEN2111;
wire  _GEN2114 = io_x[75] ? _GEN1899 : _GEN2113;
wire  _GEN2115 = io_x[25] ? _GEN2114 : _GEN2110;
wire  _GEN2116 = io_x[37] ? _GEN2115 : _GEN2103;
wire  _GEN2117 = io_x[39] ? _GEN2116 : _GEN2096;
wire  _GEN2118 = io_x[72] ? _GEN2117 : _GEN2072;
wire  _GEN2119 = io_x[29] ? _GEN2118 : _GEN2027;
wire  _GEN2120 = io_x[18] ? _GEN2119 : _GEN1924;
wire  _GEN2121 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2122 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2123 = io_x[17] ? _GEN2122 : _GEN2121;
wire  _GEN2124 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2125 = io_x[17] ? _GEN2124 : _GEN1731;
wire  _GEN2126 = io_x[75] ? _GEN2125 : _GEN2123;
wire  _GEN2127 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2128 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2129 = io_x[17] ? _GEN2128 : _GEN2127;
wire  _GEN2130 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2131 = io_x[17] ? _GEN1731 : _GEN2130;
wire  _GEN2132 = io_x[75] ? _GEN2131 : _GEN2129;
wire  _GEN2133 = io_x[25] ? _GEN2132 : _GEN2126;
wire  _GEN2134 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2135 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2136 = io_x[17] ? _GEN2135 : _GEN2134;
wire  _GEN2137 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2138 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2139 = io_x[17] ? _GEN2138 : _GEN2137;
wire  _GEN2140 = io_x[75] ? _GEN2139 : _GEN2136;
wire  _GEN2141 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2142 = io_x[17] ? _GEN1731 : _GEN2141;
wire  _GEN2143 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2144 = io_x[17] ? _GEN1711 : _GEN2143;
wire  _GEN2145 = io_x[75] ? _GEN2144 : _GEN2142;
wire  _GEN2146 = io_x[25] ? _GEN2145 : _GEN2140;
wire  _GEN2147 = io_x[37] ? _GEN2146 : _GEN2133;
wire  _GEN2148 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2149 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2150 = io_x[17] ? _GEN2149 : _GEN2148;
wire  _GEN2151 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2152 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2153 = io_x[17] ? _GEN2152 : _GEN2151;
wire  _GEN2154 = io_x[75] ? _GEN2153 : _GEN2150;
wire  _GEN2155 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2156 = io_x[17] ? _GEN1731 : _GEN2155;
wire  _GEN2157 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2158 = io_x[17] ? _GEN1711 : _GEN2157;
wire  _GEN2159 = io_x[75] ? _GEN2158 : _GEN2156;
wire  _GEN2160 = io_x[25] ? _GEN2159 : _GEN2154;
wire  _GEN2161 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2162 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2163 = io_x[17] ? _GEN2162 : _GEN2161;
wire  _GEN2164 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2165 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2166 = io_x[17] ? _GEN2165 : _GEN2164;
wire  _GEN2167 = io_x[75] ? _GEN2166 : _GEN2163;
wire  _GEN2168 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2169 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2170 = io_x[17] ? _GEN2169 : _GEN2168;
wire  _GEN2171 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2172 = io_x[17] ? _GEN1731 : _GEN2171;
wire  _GEN2173 = io_x[75] ? _GEN2172 : _GEN2170;
wire  _GEN2174 = io_x[25] ? _GEN2173 : _GEN2167;
wire  _GEN2175 = io_x[37] ? _GEN2174 : _GEN2160;
wire  _GEN2176 = io_x[39] ? _GEN2175 : _GEN2147;
wire  _GEN2177 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2178 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2179 = io_x[17] ? _GEN2178 : _GEN2177;
wire  _GEN2180 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2181 = io_x[17] ? _GEN1731 : _GEN2180;
wire  _GEN2182 = io_x[75] ? _GEN2181 : _GEN2179;
wire  _GEN2183 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2184 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2185 = io_x[17] ? _GEN2184 : _GEN2183;
wire  _GEN2186 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2187 = io_x[17] ? _GEN2186 : _GEN1711;
wire  _GEN2188 = io_x[75] ? _GEN2187 : _GEN2185;
wire  _GEN2189 = io_x[25] ? _GEN2188 : _GEN2182;
wire  _GEN2190 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2191 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2192 = io_x[17] ? _GEN2191 : _GEN2190;
wire  _GEN2193 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2194 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2195 = io_x[17] ? _GEN2194 : _GEN2193;
wire  _GEN2196 = io_x[75] ? _GEN2195 : _GEN2192;
wire  _GEN2197 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2198 = io_x[17] ? _GEN2197 : _GEN1731;
wire  _GEN2199 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2200 = io_x[17] ? _GEN1731 : _GEN2199;
wire  _GEN2201 = io_x[75] ? _GEN2200 : _GEN2198;
wire  _GEN2202 = io_x[25] ? _GEN2201 : _GEN2196;
wire  _GEN2203 = io_x[37] ? _GEN2202 : _GEN2189;
wire  _GEN2204 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2205 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2206 = io_x[17] ? _GEN2205 : _GEN2204;
wire  _GEN2207 = io_x[75] ? _GEN1899 : _GEN2206;
wire  _GEN2208 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN2209 = io_x[75] ? _GEN2208 : _GEN1903;
wire  _GEN2210 = io_x[25] ? _GEN2209 : _GEN2207;
wire  _GEN2211 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2212 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2213 = io_x[17] ? _GEN2212 : _GEN2211;
wire  _GEN2214 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2215 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2216 = io_x[17] ? _GEN2215 : _GEN2214;
wire  _GEN2217 = io_x[75] ? _GEN2216 : _GEN2213;
wire  _GEN2218 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2219 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2220 = io_x[17] ? _GEN2219 : _GEN2218;
wire  _GEN2221 = io_x[75] ? _GEN1903 : _GEN2220;
wire  _GEN2222 = io_x[25] ? _GEN2221 : _GEN2217;
wire  _GEN2223 = io_x[37] ? _GEN2222 : _GEN2210;
wire  _GEN2224 = io_x[39] ? _GEN2223 : _GEN2203;
wire  _GEN2225 = io_x[72] ? _GEN2224 : _GEN2176;
wire  _GEN2226 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2227 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2228 = io_x[17] ? _GEN2227 : _GEN2226;
wire  _GEN2229 = io_x[75] ? _GEN1899 : _GEN2228;
wire  _GEN2230 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2231 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2232 = io_x[17] ? _GEN2231 : _GEN2230;
wire  _GEN2233 = io_x[75] ? _GEN1903 : _GEN2232;
wire  _GEN2234 = io_x[25] ? _GEN2233 : _GEN2229;
wire  _GEN2235 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2236 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2237 = io_x[17] ? _GEN2236 : _GEN2235;
wire  _GEN2238 = io_x[75] ? _GEN1903 : _GEN2237;
wire  _GEN2239 = 1'b0;
wire  _GEN2240 = io_x[25] ? _GEN2239 : _GEN2238;
wire  _GEN2241 = io_x[37] ? _GEN2240 : _GEN2234;
wire  _GEN2242 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2243 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2244 = io_x[17] ? _GEN2243 : _GEN2242;
wire  _GEN2245 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2246 = io_x[17] ? _GEN1711 : _GEN2245;
wire  _GEN2247 = io_x[75] ? _GEN2246 : _GEN2244;
wire  _GEN2248 = io_x[25] ? _GEN2239 : _GEN2247;
wire  _GEN2249 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2250 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2251 = io_x[17] ? _GEN2250 : _GEN2249;
wire  _GEN2252 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2253 = io_x[17] ? _GEN1711 : _GEN2252;
wire  _GEN2254 = io_x[75] ? _GEN2253 : _GEN2251;
wire  _GEN2255 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2256 = io_x[17] ? _GEN1711 : _GEN2255;
wire  _GEN2257 = io_x[75] ? _GEN1899 : _GEN2256;
wire  _GEN2258 = io_x[25] ? _GEN2257 : _GEN2254;
wire  _GEN2259 = io_x[37] ? _GEN2258 : _GEN2248;
wire  _GEN2260 = io_x[39] ? _GEN2259 : _GEN2241;
wire  _GEN2261 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2262 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2263 = io_x[17] ? _GEN2262 : _GEN2261;
wire  _GEN2264 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2265 = io_x[17] ? _GEN1731 : _GEN2264;
wire  _GEN2266 = io_x[75] ? _GEN2265 : _GEN2263;
wire  _GEN2267 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2268 = io_x[17] ? _GEN1711 : _GEN2267;
wire  _GEN2269 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2270 = io_x[17] ? _GEN1731 : _GEN2269;
wire  _GEN2271 = io_x[75] ? _GEN2270 : _GEN2268;
wire  _GEN2272 = io_x[25] ? _GEN2271 : _GEN2266;
wire  _GEN2273 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2274 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2275 = io_x[17] ? _GEN2274 : _GEN2273;
wire  _GEN2276 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2277 = io_x[17] ? _GEN1731 : _GEN2276;
wire  _GEN2278 = io_x[75] ? _GEN2277 : _GEN2275;
wire  _GEN2279 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2280 = io_x[17] ? _GEN1731 : _GEN2279;
wire  _GEN2281 = io_x[75] ? _GEN1903 : _GEN2280;
wire  _GEN2282 = io_x[25] ? _GEN2281 : _GEN2278;
wire  _GEN2283 = io_x[37] ? _GEN2282 : _GEN2272;
wire  _GEN2284 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2285 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2286 = io_x[17] ? _GEN2285 : _GEN2284;
wire  _GEN2287 = io_x[75] ? _GEN1903 : _GEN2286;
wire  _GEN2288 = 1'b1;
wire  _GEN2289 = io_x[25] ? _GEN2288 : _GEN2287;
wire  _GEN2290 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2291 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2292 = io_x[17] ? _GEN2291 : _GEN2290;
wire  _GEN2293 = io_x[75] ? _GEN1899 : _GEN2292;
wire  _GEN2294 = io_x[25] ? _GEN2239 : _GEN2293;
wire  _GEN2295 = io_x[37] ? _GEN2294 : _GEN2289;
wire  _GEN2296 = io_x[39] ? _GEN2295 : _GEN2283;
wire  _GEN2297 = io_x[72] ? _GEN2296 : _GEN2260;
wire  _GEN2298 = io_x[29] ? _GEN2297 : _GEN2225;
wire  _GEN2299 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2300 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2301 = io_x[17] ? _GEN2300 : _GEN2299;
wire  _GEN2302 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2303 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2304 = io_x[17] ? _GEN2303 : _GEN2302;
wire  _GEN2305 = io_x[75] ? _GEN2304 : _GEN2301;
wire  _GEN2306 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2307 = io_x[17] ? _GEN2306 : _GEN1711;
wire  _GEN2308 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2309 = io_x[17] ? _GEN2308 : _GEN1731;
wire  _GEN2310 = io_x[75] ? _GEN2309 : _GEN2307;
wire  _GEN2311 = io_x[25] ? _GEN2310 : _GEN2305;
wire  _GEN2312 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2313 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2314 = io_x[17] ? _GEN2313 : _GEN2312;
wire  _GEN2315 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2316 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2317 = io_x[17] ? _GEN2316 : _GEN2315;
wire  _GEN2318 = io_x[75] ? _GEN2317 : _GEN2314;
wire  _GEN2319 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2320 = io_x[17] ? _GEN2319 : _GEN1711;
wire  _GEN2321 = io_x[75] ? _GEN1899 : _GEN2320;
wire  _GEN2322 = io_x[25] ? _GEN2321 : _GEN2318;
wire  _GEN2323 = io_x[37] ? _GEN2322 : _GEN2311;
wire  _GEN2324 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2325 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2326 = io_x[17] ? _GEN2325 : _GEN2324;
wire  _GEN2327 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2328 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2329 = io_x[17] ? _GEN2328 : _GEN2327;
wire  _GEN2330 = io_x[75] ? _GEN2329 : _GEN2326;
wire  _GEN2331 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2332 = io_x[17] ? _GEN2331 : _GEN1731;
wire  _GEN2333 = io_x[75] ? _GEN1899 : _GEN2332;
wire  _GEN2334 = io_x[25] ? _GEN2333 : _GEN2330;
wire  _GEN2335 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2336 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2337 = io_x[17] ? _GEN2336 : _GEN2335;
wire  _GEN2338 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2339 = io_x[17] ? _GEN2338 : _GEN1711;
wire  _GEN2340 = io_x[75] ? _GEN2339 : _GEN2337;
wire  _GEN2341 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2342 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2343 = io_x[17] ? _GEN2342 : _GEN2341;
wire  _GEN2344 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2345 = io_x[17] ? _GEN2344 : _GEN1731;
wire  _GEN2346 = io_x[75] ? _GEN2345 : _GEN2343;
wire  _GEN2347 = io_x[25] ? _GEN2346 : _GEN2340;
wire  _GEN2348 = io_x[37] ? _GEN2347 : _GEN2334;
wire  _GEN2349 = io_x[39] ? _GEN2348 : _GEN2323;
wire  _GEN2350 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2351 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2352 = io_x[17] ? _GEN2351 : _GEN2350;
wire  _GEN2353 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2354 = io_x[17] ? _GEN2353 : _GEN1711;
wire  _GEN2355 = io_x[75] ? _GEN2354 : _GEN2352;
wire  _GEN2356 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2357 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2358 = io_x[17] ? _GEN2357 : _GEN2356;
wire  _GEN2359 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2360 = io_x[17] ? _GEN2359 : _GEN1731;
wire  _GEN2361 = io_x[75] ? _GEN2360 : _GEN2358;
wire  _GEN2362 = io_x[25] ? _GEN2361 : _GEN2355;
wire  _GEN2363 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2364 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2365 = io_x[17] ? _GEN2364 : _GEN2363;
wire  _GEN2366 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2367 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2368 = io_x[17] ? _GEN2367 : _GEN2366;
wire  _GEN2369 = io_x[75] ? _GEN2368 : _GEN2365;
wire  _GEN2370 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2371 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2372 = io_x[17] ? _GEN2371 : _GEN2370;
wire  _GEN2373 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2374 = io_x[17] ? _GEN2373 : _GEN1711;
wire  _GEN2375 = io_x[75] ? _GEN2374 : _GEN2372;
wire  _GEN2376 = io_x[25] ? _GEN2375 : _GEN2369;
wire  _GEN2377 = io_x[37] ? _GEN2376 : _GEN2362;
wire  _GEN2378 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2379 = io_x[17] ? _GEN2378 : _GEN1731;
wire  _GEN2380 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2381 = io_x[17] ? _GEN2380 : _GEN1711;
wire  _GEN2382 = io_x[75] ? _GEN2381 : _GEN2379;
wire  _GEN2383 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2384 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2385 = io_x[17] ? _GEN2384 : _GEN2383;
wire  _GEN2386 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2387 = io_x[17] ? _GEN2386 : _GEN1731;
wire  _GEN2388 = io_x[75] ? _GEN2387 : _GEN2385;
wire  _GEN2389 = io_x[25] ? _GEN2388 : _GEN2382;
wire  _GEN2390 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2391 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2392 = io_x[17] ? _GEN2391 : _GEN2390;
wire  _GEN2393 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2394 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2395 = io_x[17] ? _GEN2394 : _GEN2393;
wire  _GEN2396 = io_x[75] ? _GEN2395 : _GEN2392;
wire  _GEN2397 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2398 = io_x[17] ? _GEN2397 : _GEN1711;
wire  _GEN2399 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2400 = io_x[17] ? _GEN2399 : _GEN1731;
wire  _GEN2401 = io_x[75] ? _GEN2400 : _GEN2398;
wire  _GEN2402 = io_x[25] ? _GEN2401 : _GEN2396;
wire  _GEN2403 = io_x[37] ? _GEN2402 : _GEN2389;
wire  _GEN2404 = io_x[39] ? _GEN2403 : _GEN2377;
wire  _GEN2405 = io_x[72] ? _GEN2404 : _GEN2349;
wire  _GEN2406 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2407 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2408 = io_x[17] ? _GEN2407 : _GEN2406;
wire  _GEN2409 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2410 = io_x[17] ? _GEN2409 : _GEN1711;
wire  _GEN2411 = io_x[75] ? _GEN2410 : _GEN2408;
wire  _GEN2412 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2413 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2414 = io_x[17] ? _GEN2413 : _GEN2412;
wire  _GEN2415 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN2416 = io_x[75] ? _GEN2415 : _GEN2414;
wire  _GEN2417 = io_x[25] ? _GEN2416 : _GEN2411;
wire  _GEN2418 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2419 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2420 = io_x[17] ? _GEN2419 : _GEN2418;
wire  _GEN2421 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2422 = io_x[17] ? _GEN2421 : _GEN1711;
wire  _GEN2423 = io_x[75] ? _GEN2422 : _GEN2420;
wire  _GEN2424 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2425 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2426 = io_x[17] ? _GEN2425 : _GEN2424;
wire  _GEN2427 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2428 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2429 = io_x[17] ? _GEN2428 : _GEN2427;
wire  _GEN2430 = io_x[75] ? _GEN2429 : _GEN2426;
wire  _GEN2431 = io_x[25] ? _GEN2430 : _GEN2423;
wire  _GEN2432 = io_x[37] ? _GEN2431 : _GEN2417;
wire  _GEN2433 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2434 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2435 = io_x[17] ? _GEN2434 : _GEN2433;
wire  _GEN2436 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2437 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2438 = io_x[17] ? _GEN2437 : _GEN2436;
wire  _GEN2439 = io_x[75] ? _GEN2438 : _GEN2435;
wire  _GEN2440 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2441 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2442 = io_x[17] ? _GEN2441 : _GEN2440;
wire  _GEN2443 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2444 = io_x[17] ? _GEN1731 : _GEN2443;
wire  _GEN2445 = io_x[75] ? _GEN2444 : _GEN2442;
wire  _GEN2446 = io_x[25] ? _GEN2445 : _GEN2439;
wire  _GEN2447 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2448 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2449 = io_x[17] ? _GEN2448 : _GEN2447;
wire  _GEN2450 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2451 = io_x[17] ? _GEN2450 : _GEN1731;
wire  _GEN2452 = io_x[75] ? _GEN2451 : _GEN2449;
wire  _GEN2453 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2454 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2455 = io_x[17] ? _GEN2454 : _GEN2453;
wire  _GEN2456 = io_x[75] ? _GEN1903 : _GEN2455;
wire  _GEN2457 = io_x[25] ? _GEN2456 : _GEN2452;
wire  _GEN2458 = io_x[37] ? _GEN2457 : _GEN2446;
wire  _GEN2459 = io_x[39] ? _GEN2458 : _GEN2432;
wire  _GEN2460 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2461 = io_x[17] ? _GEN2460 : _GEN1731;
wire  _GEN2462 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2463 = io_x[17] ? _GEN2462 : _GEN1731;
wire  _GEN2464 = io_x[75] ? _GEN2463 : _GEN2461;
wire  _GEN2465 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2466 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2467 = io_x[17] ? _GEN2466 : _GEN2465;
wire  _GEN2468 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2469 = io_x[17] ? _GEN2468 : _GEN1711;
wire  _GEN2470 = io_x[75] ? _GEN2469 : _GEN2467;
wire  _GEN2471 = io_x[25] ? _GEN2470 : _GEN2464;
wire  _GEN2472 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2473 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2474 = io_x[17] ? _GEN2473 : _GEN2472;
wire  _GEN2475 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2476 = io_x[17] ? _GEN2475 : _GEN1731;
wire  _GEN2477 = io_x[75] ? _GEN2476 : _GEN2474;
wire  _GEN2478 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2479 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2480 = io_x[17] ? _GEN2479 : _GEN2478;
wire  _GEN2481 = io_x[75] ? _GEN1903 : _GEN2480;
wire  _GEN2482 = io_x[25] ? _GEN2481 : _GEN2477;
wire  _GEN2483 = io_x[37] ? _GEN2482 : _GEN2471;
wire  _GEN2484 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2485 = io_x[17] ? _GEN2484 : _GEN1731;
wire  _GEN2486 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2487 = io_x[17] ? _GEN2486 : _GEN1731;
wire  _GEN2488 = io_x[75] ? _GEN2487 : _GEN2485;
wire  _GEN2489 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2490 = io_x[17] ? _GEN2489 : _GEN1731;
wire  _GEN2491 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2492 = io_x[17] ? _GEN2491 : _GEN1711;
wire  _GEN2493 = io_x[75] ? _GEN2492 : _GEN2490;
wire  _GEN2494 = io_x[25] ? _GEN2493 : _GEN2488;
wire  _GEN2495 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2496 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2497 = io_x[17] ? _GEN2496 : _GEN2495;
wire  _GEN2498 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2499 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2500 = io_x[17] ? _GEN2499 : _GEN2498;
wire  _GEN2501 = io_x[75] ? _GEN2500 : _GEN2497;
wire  _GEN2502 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2503 = io_x[17] ? _GEN2502 : _GEN1731;
wire  _GEN2504 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2505 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2506 = io_x[17] ? _GEN2505 : _GEN2504;
wire  _GEN2507 = io_x[75] ? _GEN2506 : _GEN2503;
wire  _GEN2508 = io_x[25] ? _GEN2507 : _GEN2501;
wire  _GEN2509 = io_x[37] ? _GEN2508 : _GEN2494;
wire  _GEN2510 = io_x[39] ? _GEN2509 : _GEN2483;
wire  _GEN2511 = io_x[72] ? _GEN2510 : _GEN2459;
wire  _GEN2512 = io_x[29] ? _GEN2511 : _GEN2405;
wire  _GEN2513 = io_x[18] ? _GEN2512 : _GEN2298;
wire  _GEN2514 = io_x[19] ? _GEN2513 : _GEN2120;
wire  _GEN2515 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2516 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2517 = io_x[17] ? _GEN2516 : _GEN2515;
wire  _GEN2518 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2519 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2520 = io_x[17] ? _GEN2519 : _GEN2518;
wire  _GEN2521 = io_x[75] ? _GEN2520 : _GEN2517;
wire  _GEN2522 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2523 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2524 = io_x[17] ? _GEN2523 : _GEN2522;
wire  _GEN2525 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2526 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2527 = io_x[17] ? _GEN2526 : _GEN2525;
wire  _GEN2528 = io_x[75] ? _GEN2527 : _GEN2524;
wire  _GEN2529 = io_x[25] ? _GEN2528 : _GEN2521;
wire  _GEN2530 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2531 = io_x[17] ? _GEN2530 : _GEN1711;
wire  _GEN2532 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2533 = io_x[17] ? _GEN1731 : _GEN2532;
wire  _GEN2534 = io_x[75] ? _GEN2533 : _GEN2531;
wire  _GEN2535 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2536 = io_x[17] ? _GEN2535 : _GEN1731;
wire  _GEN2537 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2538 = io_x[17] ? _GEN1731 : _GEN2537;
wire  _GEN2539 = io_x[75] ? _GEN2538 : _GEN2536;
wire  _GEN2540 = io_x[25] ? _GEN2539 : _GEN2534;
wire  _GEN2541 = io_x[37] ? _GEN2540 : _GEN2529;
wire  _GEN2542 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2543 = io_x[17] ? _GEN1731 : _GEN2542;
wire  _GEN2544 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2545 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2546 = io_x[17] ? _GEN2545 : _GEN2544;
wire  _GEN2547 = io_x[75] ? _GEN2546 : _GEN2543;
wire  _GEN2548 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2549 = io_x[17] ? _GEN1731 : _GEN2548;
wire  _GEN2550 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2551 = io_x[17] ? _GEN1731 : _GEN2550;
wire  _GEN2552 = io_x[75] ? _GEN2551 : _GEN2549;
wire  _GEN2553 = io_x[25] ? _GEN2552 : _GEN2547;
wire  _GEN2554 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2555 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2556 = io_x[17] ? _GEN2555 : _GEN2554;
wire  _GEN2557 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2558 = io_x[17] ? _GEN1731 : _GEN2557;
wire  _GEN2559 = io_x[75] ? _GEN2558 : _GEN2556;
wire  _GEN2560 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2561 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2562 = io_x[17] ? _GEN2561 : _GEN2560;
wire  _GEN2563 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2564 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2565 = io_x[17] ? _GEN2564 : _GEN2563;
wire  _GEN2566 = io_x[75] ? _GEN2565 : _GEN2562;
wire  _GEN2567 = io_x[25] ? _GEN2566 : _GEN2559;
wire  _GEN2568 = io_x[37] ? _GEN2567 : _GEN2553;
wire  _GEN2569 = io_x[39] ? _GEN2568 : _GEN2541;
wire  _GEN2570 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2571 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2572 = io_x[17] ? _GEN2571 : _GEN2570;
wire  _GEN2573 = io_x[75] ? _GEN1899 : _GEN2572;
wire  _GEN2574 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2575 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2576 = io_x[17] ? _GEN2575 : _GEN2574;
wire  _GEN2577 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2578 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2579 = io_x[17] ? _GEN2578 : _GEN2577;
wire  _GEN2580 = io_x[75] ? _GEN2579 : _GEN2576;
wire  _GEN2581 = io_x[25] ? _GEN2580 : _GEN2573;
wire  _GEN2582 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2583 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2584 = io_x[17] ? _GEN2583 : _GEN2582;
wire  _GEN2585 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2586 = io_x[17] ? _GEN1731 : _GEN2585;
wire  _GEN2587 = io_x[75] ? _GEN2586 : _GEN2584;
wire  _GEN2588 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2589 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2590 = io_x[17] ? _GEN2589 : _GEN2588;
wire  _GEN2591 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2592 = io_x[17] ? _GEN1711 : _GEN2591;
wire  _GEN2593 = io_x[75] ? _GEN2592 : _GEN2590;
wire  _GEN2594 = io_x[25] ? _GEN2593 : _GEN2587;
wire  _GEN2595 = io_x[37] ? _GEN2594 : _GEN2581;
wire  _GEN2596 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2597 = io_x[17] ? _GEN1711 : _GEN2596;
wire  _GEN2598 = io_x[75] ? _GEN1899 : _GEN2597;
wire  _GEN2599 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2600 = io_x[17] ? _GEN1711 : _GEN2599;
wire  _GEN2601 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN2602 = io_x[75] ? _GEN2601 : _GEN2600;
wire  _GEN2603 = io_x[25] ? _GEN2602 : _GEN2598;
wire  _GEN2604 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2605 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2606 = io_x[17] ? _GEN2605 : _GEN2604;
wire  _GEN2607 = io_x[75] ? _GEN1899 : _GEN2606;
wire  _GEN2608 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2609 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2610 = io_x[17] ? _GEN2609 : _GEN2608;
wire  _GEN2611 = io_x[75] ? _GEN1899 : _GEN2610;
wire  _GEN2612 = io_x[25] ? _GEN2611 : _GEN2607;
wire  _GEN2613 = io_x[37] ? _GEN2612 : _GEN2603;
wire  _GEN2614 = io_x[39] ? _GEN2613 : _GEN2595;
wire  _GEN2615 = io_x[72] ? _GEN2614 : _GEN2569;
wire  _GEN2616 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2617 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2618 = io_x[17] ? _GEN2617 : _GEN2616;
wire  _GEN2619 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2620 = io_x[17] ? _GEN1731 : _GEN2619;
wire  _GEN2621 = io_x[75] ? _GEN2620 : _GEN2618;
wire  _GEN2622 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2623 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2624 = io_x[17] ? _GEN2623 : _GEN2622;
wire  _GEN2625 = io_x[75] ? _GEN1903 : _GEN2624;
wire  _GEN2626 = io_x[25] ? _GEN2625 : _GEN2621;
wire  _GEN2627 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2628 = io_x[17] ? _GEN1731 : _GEN2627;
wire  _GEN2629 = io_x[75] ? _GEN2628 : _GEN1903;
wire  _GEN2630 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2631 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2632 = io_x[17] ? _GEN2631 : _GEN2630;
wire  _GEN2633 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2634 = io_x[17] ? _GEN1731 : _GEN2633;
wire  _GEN2635 = io_x[75] ? _GEN2634 : _GEN2632;
wire  _GEN2636 = io_x[25] ? _GEN2635 : _GEN2629;
wire  _GEN2637 = io_x[37] ? _GEN2636 : _GEN2626;
wire  _GEN2638 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2639 = io_x[17] ? _GEN1731 : _GEN2638;
wire  _GEN2640 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2641 = io_x[17] ? _GEN1731 : _GEN2640;
wire  _GEN2642 = io_x[75] ? _GEN2641 : _GEN2639;
wire  _GEN2643 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2644 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2645 = io_x[17] ? _GEN2644 : _GEN2643;
wire  _GEN2646 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2647 = io_x[17] ? _GEN1731 : _GEN2646;
wire  _GEN2648 = io_x[75] ? _GEN2647 : _GEN2645;
wire  _GEN2649 = io_x[25] ? _GEN2648 : _GEN2642;
wire  _GEN2650 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2651 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2652 = io_x[17] ? _GEN2651 : _GEN2650;
wire  _GEN2653 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2654 = io_x[17] ? _GEN1731 : _GEN2653;
wire  _GEN2655 = io_x[75] ? _GEN2654 : _GEN2652;
wire  _GEN2656 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2657 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2658 = io_x[17] ? _GEN2657 : _GEN2656;
wire  _GEN2659 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2660 = io_x[17] ? _GEN1731 : _GEN2659;
wire  _GEN2661 = io_x[75] ? _GEN2660 : _GEN2658;
wire  _GEN2662 = io_x[25] ? _GEN2661 : _GEN2655;
wire  _GEN2663 = io_x[37] ? _GEN2662 : _GEN2649;
wire  _GEN2664 = io_x[39] ? _GEN2663 : _GEN2637;
wire  _GEN2665 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2666 = io_x[17] ? _GEN1711 : _GEN2665;
wire  _GEN2667 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2668 = io_x[17] ? _GEN1731 : _GEN2667;
wire  _GEN2669 = io_x[75] ? _GEN2668 : _GEN2666;
wire  _GEN2670 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2671 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2672 = io_x[17] ? _GEN2671 : _GEN2670;
wire  _GEN2673 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2674 = io_x[17] ? _GEN1731 : _GEN2673;
wire  _GEN2675 = io_x[75] ? _GEN2674 : _GEN2672;
wire  _GEN2676 = io_x[25] ? _GEN2675 : _GEN2669;
wire  _GEN2677 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2678 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2679 = io_x[17] ? _GEN2678 : _GEN2677;
wire  _GEN2680 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2681 = io_x[17] ? _GEN1731 : _GEN2680;
wire  _GEN2682 = io_x[75] ? _GEN2681 : _GEN2679;
wire  _GEN2683 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2684 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2685 = io_x[17] ? _GEN2684 : _GEN2683;
wire  _GEN2686 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2687 = io_x[17] ? _GEN1731 : _GEN2686;
wire  _GEN2688 = io_x[75] ? _GEN2687 : _GEN2685;
wire  _GEN2689 = io_x[25] ? _GEN2688 : _GEN2682;
wire  _GEN2690 = io_x[37] ? _GEN2689 : _GEN2676;
wire  _GEN2691 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2692 = io_x[17] ? _GEN1731 : _GEN2691;
wire  _GEN2693 = io_x[75] ? _GEN1899 : _GEN2692;
wire  _GEN2694 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2695 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2696 = io_x[17] ? _GEN2695 : _GEN2694;
wire  _GEN2697 = io_x[75] ? _GEN1899 : _GEN2696;
wire  _GEN2698 = io_x[25] ? _GEN2697 : _GEN2693;
wire  _GEN2699 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2700 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2701 = io_x[17] ? _GEN2700 : _GEN2699;
wire  _GEN2702 = io_x[75] ? _GEN1899 : _GEN2701;
wire  _GEN2703 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2704 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2705 = io_x[17] ? _GEN2704 : _GEN2703;
wire  _GEN2706 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2707 = io_x[17] ? _GEN2706 : _GEN1731;
wire  _GEN2708 = io_x[75] ? _GEN2707 : _GEN2705;
wire  _GEN2709 = io_x[25] ? _GEN2708 : _GEN2702;
wire  _GEN2710 = io_x[37] ? _GEN2709 : _GEN2698;
wire  _GEN2711 = io_x[39] ? _GEN2710 : _GEN2690;
wire  _GEN2712 = io_x[72] ? _GEN2711 : _GEN2664;
wire  _GEN2713 = io_x[29] ? _GEN2712 : _GEN2615;
wire  _GEN2714 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2715 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2716 = io_x[17] ? _GEN2715 : _GEN2714;
wire  _GEN2717 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN2718 = io_x[75] ? _GEN2717 : _GEN2716;
wire  _GEN2719 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2720 = io_x[17] ? _GEN2719 : _GEN1731;
wire  _GEN2721 = io_x[75] ? _GEN1903 : _GEN2720;
wire  _GEN2722 = io_x[25] ? _GEN2721 : _GEN2718;
wire  _GEN2723 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2724 = io_x[17] ? _GEN1731 : _GEN2723;
wire  _GEN2725 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2726 = io_x[17] ? _GEN1711 : _GEN2725;
wire  _GEN2727 = io_x[75] ? _GEN2726 : _GEN2724;
wire  _GEN2728 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2729 = io_x[17] ? _GEN2728 : _GEN1731;
wire  _GEN2730 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2731 = io_x[17] ? _GEN2730 : _GEN1731;
wire  _GEN2732 = io_x[75] ? _GEN2731 : _GEN2729;
wire  _GEN2733 = io_x[25] ? _GEN2732 : _GEN2727;
wire  _GEN2734 = io_x[37] ? _GEN2733 : _GEN2722;
wire  _GEN2735 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2736 = io_x[17] ? _GEN2735 : _GEN1731;
wire  _GEN2737 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2738 = io_x[17] ? _GEN1711 : _GEN2737;
wire  _GEN2739 = io_x[75] ? _GEN2738 : _GEN2736;
wire  _GEN2740 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2741 = io_x[17] ? _GEN2740 : _GEN1731;
wire  _GEN2742 = io_x[75] ? _GEN2741 : _GEN1903;
wire  _GEN2743 = io_x[25] ? _GEN2742 : _GEN2739;
wire  _GEN2744 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2745 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2746 = io_x[17] ? _GEN2745 : _GEN2744;
wire  _GEN2747 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2748 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2749 = io_x[17] ? _GEN2748 : _GEN2747;
wire  _GEN2750 = io_x[75] ? _GEN2749 : _GEN2746;
wire  _GEN2751 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2752 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2753 = io_x[17] ? _GEN2752 : _GEN2751;
wire  _GEN2754 = io_x[75] ? _GEN1903 : _GEN2753;
wire  _GEN2755 = io_x[25] ? _GEN2754 : _GEN2750;
wire  _GEN2756 = io_x[37] ? _GEN2755 : _GEN2743;
wire  _GEN2757 = io_x[39] ? _GEN2756 : _GEN2734;
wire  _GEN2758 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2759 = io_x[17] ? _GEN1731 : _GEN2758;
wire  _GEN2760 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2761 = io_x[17] ? _GEN1711 : _GEN2760;
wire  _GEN2762 = io_x[75] ? _GEN2761 : _GEN2759;
wire  _GEN2763 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2764 = io_x[17] ? _GEN2763 : _GEN1731;
wire  _GEN2765 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2766 = io_x[17] ? _GEN2765 : _GEN1731;
wire  _GEN2767 = io_x[75] ? _GEN2766 : _GEN2764;
wire  _GEN2768 = io_x[25] ? _GEN2767 : _GEN2762;
wire  _GEN2769 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2770 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2771 = io_x[17] ? _GEN2770 : _GEN2769;
wire  _GEN2772 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2773 = io_x[17] ? _GEN2772 : _GEN1731;
wire  _GEN2774 = io_x[75] ? _GEN2773 : _GEN2771;
wire  _GEN2775 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2776 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2777 = io_x[17] ? _GEN2776 : _GEN2775;
wire  _GEN2778 = io_x[75] ? _GEN1899 : _GEN2777;
wire  _GEN2779 = io_x[25] ? _GEN2778 : _GEN2774;
wire  _GEN2780 = io_x[37] ? _GEN2779 : _GEN2768;
wire  _GEN2781 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2782 = io_x[17] ? _GEN2781 : _GEN1731;
wire  _GEN2783 = io_x[75] ? _GEN1903 : _GEN2782;
wire  _GEN2784 = io_x[25] ? _GEN2783 : _GEN2288;
wire  _GEN2785 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2786 = io_x[17] ? _GEN1731 : _GEN2785;
wire  _GEN2787 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2788 = io_x[17] ? _GEN1731 : _GEN2787;
wire  _GEN2789 = io_x[75] ? _GEN2788 : _GEN2786;
wire  _GEN2790 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2791 = io_x[17] ? _GEN2790 : _GEN1731;
wire  _GEN2792 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN2793 = io_x[75] ? _GEN2792 : _GEN2791;
wire  _GEN2794 = io_x[25] ? _GEN2793 : _GEN2789;
wire  _GEN2795 = io_x[37] ? _GEN2794 : _GEN2784;
wire  _GEN2796 = io_x[39] ? _GEN2795 : _GEN2780;
wire  _GEN2797 = io_x[72] ? _GEN2796 : _GEN2757;
wire  _GEN2798 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2799 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2800 = io_x[17] ? _GEN2799 : _GEN2798;
wire  _GEN2801 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN2802 = io_x[75] ? _GEN2801 : _GEN2800;
wire  _GEN2803 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2804 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2805 = io_x[17] ? _GEN2804 : _GEN2803;
wire  _GEN2806 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN2807 = io_x[75] ? _GEN2806 : _GEN2805;
wire  _GEN2808 = io_x[25] ? _GEN2807 : _GEN2802;
wire  _GEN2809 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2810 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2811 = io_x[17] ? _GEN2810 : _GEN2809;
wire  _GEN2812 = io_x[75] ? _GEN1903 : _GEN2811;
wire  _GEN2813 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2814 = io_x[17] ? _GEN2813 : _GEN1731;
wire  _GEN2815 = io_x[75] ? _GEN1899 : _GEN2814;
wire  _GEN2816 = io_x[25] ? _GEN2815 : _GEN2812;
wire  _GEN2817 = io_x[37] ? _GEN2816 : _GEN2808;
wire  _GEN2818 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2819 = io_x[17] ? _GEN1731 : _GEN2818;
wire  _GEN2820 = io_x[75] ? _GEN2819 : _GEN1899;
wire  _GEN2821 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2822 = io_x[17] ? _GEN2821 : _GEN1711;
wire  _GEN2823 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2824 = io_x[17] ? _GEN1731 : _GEN2823;
wire  _GEN2825 = io_x[75] ? _GEN2824 : _GEN2822;
wire  _GEN2826 = io_x[25] ? _GEN2825 : _GEN2820;
wire  _GEN2827 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2828 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2829 = io_x[17] ? _GEN2828 : _GEN2827;
wire  _GEN2830 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2831 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2832 = io_x[17] ? _GEN2831 : _GEN2830;
wire  _GEN2833 = io_x[75] ? _GEN2832 : _GEN2829;
wire  _GEN2834 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2835 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2836 = io_x[17] ? _GEN2835 : _GEN2834;
wire  _GEN2837 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2838 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2839 = io_x[17] ? _GEN2838 : _GEN2837;
wire  _GEN2840 = io_x[75] ? _GEN2839 : _GEN2836;
wire  _GEN2841 = io_x[25] ? _GEN2840 : _GEN2833;
wire  _GEN2842 = io_x[37] ? _GEN2841 : _GEN2826;
wire  _GEN2843 = io_x[39] ? _GEN2842 : _GEN2817;
wire  _GEN2844 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2845 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2846 = io_x[17] ? _GEN2845 : _GEN2844;
wire  _GEN2847 = io_x[75] ? _GEN1899 : _GEN2846;
wire  _GEN2848 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2849 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2850 = io_x[17] ? _GEN2849 : _GEN2848;
wire  _GEN2851 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2852 = io_x[17] ? _GEN2851 : _GEN1731;
wire  _GEN2853 = io_x[75] ? _GEN2852 : _GEN2850;
wire  _GEN2854 = io_x[25] ? _GEN2853 : _GEN2847;
wire  _GEN2855 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2856 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2857 = io_x[17] ? _GEN2856 : _GEN2855;
wire  _GEN2858 = io_x[75] ? _GEN1899 : _GEN2857;
wire  _GEN2859 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2860 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2861 = io_x[17] ? _GEN2860 : _GEN2859;
wire  _GEN2862 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2863 = io_x[17] ? _GEN1711 : _GEN2862;
wire  _GEN2864 = io_x[75] ? _GEN2863 : _GEN2861;
wire  _GEN2865 = io_x[25] ? _GEN2864 : _GEN2858;
wire  _GEN2866 = io_x[37] ? _GEN2865 : _GEN2854;
wire  _GEN2867 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN2868 = io_x[75] ? _GEN2867 : _GEN1899;
wire  _GEN2869 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2870 = io_x[17] ? _GEN2869 : _GEN1731;
wire  _GEN2871 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2872 = io_x[17] ? _GEN2871 : _GEN1731;
wire  _GEN2873 = io_x[75] ? _GEN2872 : _GEN2870;
wire  _GEN2874 = io_x[25] ? _GEN2873 : _GEN2868;
wire  _GEN2875 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2876 = io_x[17] ? _GEN1711 : _GEN2875;
wire  _GEN2877 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2878 = io_x[17] ? _GEN1731 : _GEN2877;
wire  _GEN2879 = io_x[75] ? _GEN2878 : _GEN2876;
wire  _GEN2880 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2881 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2882 = io_x[17] ? _GEN2881 : _GEN2880;
wire  _GEN2883 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2884 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2885 = io_x[17] ? _GEN2884 : _GEN2883;
wire  _GEN2886 = io_x[75] ? _GEN2885 : _GEN2882;
wire  _GEN2887 = io_x[25] ? _GEN2886 : _GEN2879;
wire  _GEN2888 = io_x[37] ? _GEN2887 : _GEN2874;
wire  _GEN2889 = io_x[39] ? _GEN2888 : _GEN2866;
wire  _GEN2890 = io_x[72] ? _GEN2889 : _GEN2843;
wire  _GEN2891 = io_x[29] ? _GEN2890 : _GEN2797;
wire  _GEN2892 = io_x[18] ? _GEN2891 : _GEN2713;
wire  _GEN2893 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2894 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2895 = io_x[17] ? _GEN2894 : _GEN2893;
wire  _GEN2896 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2897 = io_x[17] ? _GEN1731 : _GEN2896;
wire  _GEN2898 = io_x[75] ? _GEN2897 : _GEN2895;
wire  _GEN2899 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2900 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2901 = io_x[17] ? _GEN2900 : _GEN2899;
wire  _GEN2902 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN2903 = io_x[75] ? _GEN2902 : _GEN2901;
wire  _GEN2904 = io_x[25] ? _GEN2903 : _GEN2898;
wire  _GEN2905 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2906 = io_x[17] ? _GEN1731 : _GEN2905;
wire  _GEN2907 = io_x[75] ? _GEN1899 : _GEN2906;
wire  _GEN2908 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2909 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2910 = io_x[17] ? _GEN2909 : _GEN2908;
wire  _GEN2911 = io_x[75] ? _GEN1899 : _GEN2910;
wire  _GEN2912 = io_x[25] ? _GEN2911 : _GEN2907;
wire  _GEN2913 = io_x[37] ? _GEN2912 : _GEN2904;
wire  _GEN2914 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2915 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2916 = io_x[17] ? _GEN2915 : _GEN2914;
wire  _GEN2917 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2918 = io_x[17] ? _GEN1731 : _GEN2917;
wire  _GEN2919 = io_x[75] ? _GEN2918 : _GEN2916;
wire  _GEN2920 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2921 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2922 = io_x[17] ? _GEN2921 : _GEN2920;
wire  _GEN2923 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2924 = io_x[17] ? _GEN1731 : _GEN2923;
wire  _GEN2925 = io_x[75] ? _GEN2924 : _GEN2922;
wire  _GEN2926 = io_x[25] ? _GEN2925 : _GEN2919;
wire  _GEN2927 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2928 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2929 = io_x[17] ? _GEN2928 : _GEN2927;
wire  _GEN2930 = io_x[75] ? _GEN1899 : _GEN2929;
wire  _GEN2931 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2932 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2933 = io_x[17] ? _GEN2932 : _GEN2931;
wire  _GEN2934 = io_x[75] ? _GEN1903 : _GEN2933;
wire  _GEN2935 = io_x[25] ? _GEN2934 : _GEN2930;
wire  _GEN2936 = io_x[37] ? _GEN2935 : _GEN2926;
wire  _GEN2937 = io_x[39] ? _GEN2936 : _GEN2913;
wire  _GEN2938 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2939 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2940 = io_x[17] ? _GEN2939 : _GEN2938;
wire  _GEN2941 = io_x[75] ? _GEN1899 : _GEN2940;
wire  _GEN2942 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2943 = io_x[17] ? _GEN1711 : _GEN2942;
wire  _GEN2944 = io_x[75] ? _GEN1903 : _GEN2943;
wire  _GEN2945 = io_x[25] ? _GEN2944 : _GEN2941;
wire  _GEN2946 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2947 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2948 = io_x[17] ? _GEN2947 : _GEN2946;
wire  _GEN2949 = io_x[75] ? _GEN1899 : _GEN2948;
wire  _GEN2950 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2951 = io_x[17] ? _GEN1711 : _GEN2950;
wire  _GEN2952 = io_x[75] ? _GEN1903 : _GEN2951;
wire  _GEN2953 = io_x[25] ? _GEN2952 : _GEN2949;
wire  _GEN2954 = io_x[37] ? _GEN2953 : _GEN2945;
wire  _GEN2955 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2956 = io_x[17] ? _GEN1731 : _GEN2955;
wire  _GEN2957 = io_x[75] ? _GEN1899 : _GEN2956;
wire  _GEN2958 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2959 = io_x[17] ? _GEN1731 : _GEN2958;
wire  _GEN2960 = io_x[75] ? _GEN1903 : _GEN2959;
wire  _GEN2961 = io_x[25] ? _GEN2960 : _GEN2957;
wire  _GEN2962 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2963 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2964 = io_x[17] ? _GEN2963 : _GEN2962;
wire  _GEN2965 = io_x[75] ? _GEN1899 : _GEN2964;
wire  _GEN2966 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN2967 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN2968 = io_x[75] ? _GEN2967 : _GEN2966;
wire  _GEN2969 = io_x[25] ? _GEN2968 : _GEN2965;
wire  _GEN2970 = io_x[37] ? _GEN2969 : _GEN2961;
wire  _GEN2971 = io_x[39] ? _GEN2970 : _GEN2954;
wire  _GEN2972 = io_x[72] ? _GEN2971 : _GEN2937;
wire  _GEN2973 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2974 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2975 = io_x[17] ? _GEN2974 : _GEN2973;
wire  _GEN2976 = io_x[75] ? _GEN1903 : _GEN2975;
wire  _GEN2977 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2978 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2979 = io_x[17] ? _GEN2978 : _GEN2977;
wire  _GEN2980 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2981 = io_x[17] ? _GEN1731 : _GEN2980;
wire  _GEN2982 = io_x[75] ? _GEN2981 : _GEN2979;
wire  _GEN2983 = io_x[25] ? _GEN2982 : _GEN2976;
wire  _GEN2984 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2985 = io_x[17] ? _GEN2984 : _GEN1731;
wire  _GEN2986 = io_x[75] ? _GEN1903 : _GEN2985;
wire  _GEN2987 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2988 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2989 = io_x[17] ? _GEN2988 : _GEN2987;
wire  _GEN2990 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN2991 = io_x[17] ? _GEN1731 : _GEN2990;
wire  _GEN2992 = io_x[75] ? _GEN2991 : _GEN2989;
wire  _GEN2993 = io_x[25] ? _GEN2992 : _GEN2986;
wire  _GEN2994 = io_x[37] ? _GEN2993 : _GEN2983;
wire  _GEN2995 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2996 = io_x[17] ? _GEN2995 : _GEN1731;
wire  _GEN2997 = io_x[75] ? _GEN1903 : _GEN2996;
wire  _GEN2998 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN2999 = io_x[17] ? _GEN1711 : _GEN2998;
wire  _GEN3000 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3001 = io_x[75] ? _GEN3000 : _GEN2999;
wire  _GEN3002 = io_x[25] ? _GEN3001 : _GEN2997;
wire  _GEN3003 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3004 = io_x[17] ? _GEN1711 : _GEN3003;
wire  _GEN3005 = io_x[75] ? _GEN1903 : _GEN3004;
wire  _GEN3006 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3007 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3008 = io_x[17] ? _GEN3007 : _GEN3006;
wire  _GEN3009 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3010 = io_x[17] ? _GEN1731 : _GEN3009;
wire  _GEN3011 = io_x[75] ? _GEN3010 : _GEN3008;
wire  _GEN3012 = io_x[25] ? _GEN3011 : _GEN3005;
wire  _GEN3013 = io_x[37] ? _GEN3012 : _GEN3002;
wire  _GEN3014 = io_x[39] ? _GEN3013 : _GEN2994;
wire  _GEN3015 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3016 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3017 = io_x[17] ? _GEN3016 : _GEN3015;
wire  _GEN3018 = io_x[75] ? _GEN1899 : _GEN3017;
wire  _GEN3019 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3020 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3021 = io_x[17] ? _GEN3020 : _GEN3019;
wire  _GEN3022 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3023 = io_x[75] ? _GEN3022 : _GEN3021;
wire  _GEN3024 = io_x[25] ? _GEN3023 : _GEN3018;
wire  _GEN3025 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3026 = io_x[17] ? _GEN3025 : _GEN1731;
wire  _GEN3027 = io_x[75] ? _GEN1899 : _GEN3026;
wire  _GEN3028 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3029 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3030 = io_x[17] ? _GEN3029 : _GEN3028;
wire  _GEN3031 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3032 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3033 = io_x[17] ? _GEN3032 : _GEN3031;
wire  _GEN3034 = io_x[75] ? _GEN3033 : _GEN3030;
wire  _GEN3035 = io_x[25] ? _GEN3034 : _GEN3027;
wire  _GEN3036 = io_x[37] ? _GEN3035 : _GEN3024;
wire  _GEN3037 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3038 = io_x[17] ? _GEN3037 : _GEN1711;
wire  _GEN3039 = io_x[75] ? _GEN1903 : _GEN3038;
wire  _GEN3040 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3041 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3042 = io_x[17] ? _GEN3041 : _GEN3040;
wire  _GEN3043 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3044 = io_x[17] ? _GEN1731 : _GEN3043;
wire  _GEN3045 = io_x[75] ? _GEN3044 : _GEN3042;
wire  _GEN3046 = io_x[25] ? _GEN3045 : _GEN3039;
wire  _GEN3047 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3048 = io_x[17] ? _GEN1711 : _GEN3047;
wire  _GEN3049 = io_x[75] ? _GEN1903 : _GEN3048;
wire  _GEN3050 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN3051 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3052 = io_x[17] ? _GEN1731 : _GEN3051;
wire  _GEN3053 = io_x[75] ? _GEN3052 : _GEN3050;
wire  _GEN3054 = io_x[25] ? _GEN3053 : _GEN3049;
wire  _GEN3055 = io_x[37] ? _GEN3054 : _GEN3046;
wire  _GEN3056 = io_x[39] ? _GEN3055 : _GEN3036;
wire  _GEN3057 = io_x[72] ? _GEN3056 : _GEN3014;
wire  _GEN3058 = io_x[29] ? _GEN3057 : _GEN2972;
wire  _GEN3059 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3060 = io_x[17] ? _GEN3059 : _GEN1711;
wire  _GEN3061 = io_x[75] ? _GEN1903 : _GEN3060;
wire  _GEN3062 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3063 = io_x[17] ? _GEN3062 : _GEN1731;
wire  _GEN3064 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3065 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3066 = io_x[17] ? _GEN3065 : _GEN3064;
wire  _GEN3067 = io_x[75] ? _GEN3066 : _GEN3063;
wire  _GEN3068 = io_x[25] ? _GEN3067 : _GEN3061;
wire  _GEN3069 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3070 = io_x[17] ? _GEN3069 : _GEN1711;
wire  _GEN3071 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3072 = io_x[17] ? _GEN3071 : _GEN1731;
wire  _GEN3073 = io_x[75] ? _GEN3072 : _GEN3070;
wire  _GEN3074 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3075 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3076 = io_x[17] ? _GEN3075 : _GEN3074;
wire  _GEN3077 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3078 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3079 = io_x[17] ? _GEN3078 : _GEN3077;
wire  _GEN3080 = io_x[75] ? _GEN3079 : _GEN3076;
wire  _GEN3081 = io_x[25] ? _GEN3080 : _GEN3073;
wire  _GEN3082 = io_x[37] ? _GEN3081 : _GEN3068;
wire  _GEN3083 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3084 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3085 = io_x[17] ? _GEN3084 : _GEN3083;
wire  _GEN3086 = io_x[75] ? _GEN1899 : _GEN3085;
wire  _GEN3087 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3088 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3089 = io_x[17] ? _GEN3088 : _GEN3087;
wire  _GEN3090 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3091 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3092 = io_x[17] ? _GEN3091 : _GEN3090;
wire  _GEN3093 = io_x[75] ? _GEN3092 : _GEN3089;
wire  _GEN3094 = io_x[25] ? _GEN3093 : _GEN3086;
wire  _GEN3095 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3096 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3097 = io_x[17] ? _GEN3096 : _GEN3095;
wire  _GEN3098 = io_x[75] ? _GEN1899 : _GEN3097;
wire  _GEN3099 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3100 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3101 = io_x[17] ? _GEN3100 : _GEN3099;
wire  _GEN3102 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3103 = io_x[17] ? _GEN3102 : _GEN1731;
wire  _GEN3104 = io_x[75] ? _GEN3103 : _GEN3101;
wire  _GEN3105 = io_x[25] ? _GEN3104 : _GEN3098;
wire  _GEN3106 = io_x[37] ? _GEN3105 : _GEN3094;
wire  _GEN3107 = io_x[39] ? _GEN3106 : _GEN3082;
wire  _GEN3108 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3109 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3110 = io_x[17] ? _GEN3109 : _GEN3108;
wire  _GEN3111 = io_x[75] ? _GEN1899 : _GEN3110;
wire  _GEN3112 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3113 = io_x[17] ? _GEN3112 : _GEN1731;
wire  _GEN3114 = io_x[75] ? _GEN1899 : _GEN3113;
wire  _GEN3115 = io_x[25] ? _GEN3114 : _GEN3111;
wire  _GEN3116 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3117 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3118 = io_x[17] ? _GEN3117 : _GEN3116;
wire  _GEN3119 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3120 = io_x[17] ? _GEN3119 : _GEN1731;
wire  _GEN3121 = io_x[75] ? _GEN3120 : _GEN3118;
wire  _GEN3122 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3123 = io_x[17] ? _GEN3122 : _GEN1731;
wire  _GEN3124 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3125 = io_x[17] ? _GEN1711 : _GEN3124;
wire  _GEN3126 = io_x[75] ? _GEN3125 : _GEN3123;
wire  _GEN3127 = io_x[25] ? _GEN3126 : _GEN3121;
wire  _GEN3128 = io_x[37] ? _GEN3127 : _GEN3115;
wire  _GEN3129 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3130 = io_x[17] ? _GEN3129 : _GEN1711;
wire  _GEN3131 = io_x[75] ? _GEN1903 : _GEN3130;
wire  _GEN3132 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3133 = io_x[17] ? _GEN3132 : _GEN1711;
wire  _GEN3134 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3135 = io_x[17] ? _GEN3134 : _GEN1731;
wire  _GEN3136 = io_x[75] ? _GEN3135 : _GEN3133;
wire  _GEN3137 = io_x[25] ? _GEN3136 : _GEN3131;
wire  _GEN3138 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3139 = io_x[17] ? _GEN3138 : _GEN1711;
wire  _GEN3140 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3141 = io_x[17] ? _GEN3140 : _GEN1731;
wire  _GEN3142 = io_x[75] ? _GEN3141 : _GEN3139;
wire  _GEN3143 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3144 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3145 = io_x[17] ? _GEN3144 : _GEN3143;
wire  _GEN3146 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3147 = io_x[17] ? _GEN3146 : _GEN1711;
wire  _GEN3148 = io_x[75] ? _GEN3147 : _GEN3145;
wire  _GEN3149 = io_x[25] ? _GEN3148 : _GEN3142;
wire  _GEN3150 = io_x[37] ? _GEN3149 : _GEN3137;
wire  _GEN3151 = io_x[39] ? _GEN3150 : _GEN3128;
wire  _GEN3152 = io_x[72] ? _GEN3151 : _GEN3107;
wire  _GEN3153 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3154 = io_x[17] ? _GEN3153 : _GEN1731;
wire  _GEN3155 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3156 = io_x[17] ? _GEN3155 : _GEN1731;
wire  _GEN3157 = io_x[75] ? _GEN3156 : _GEN3154;
wire  _GEN3158 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3159 = io_x[17] ? _GEN3158 : _GEN1731;
wire  _GEN3160 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3161 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3162 = io_x[17] ? _GEN3161 : _GEN3160;
wire  _GEN3163 = io_x[75] ? _GEN3162 : _GEN3159;
wire  _GEN3164 = io_x[25] ? _GEN3163 : _GEN3157;
wire  _GEN3165 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3166 = io_x[17] ? _GEN3165 : _GEN1711;
wire  _GEN3167 = io_x[75] ? _GEN1903 : _GEN3166;
wire  _GEN3168 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3169 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3170 = io_x[17] ? _GEN3169 : _GEN3168;
wire  _GEN3171 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3172 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3173 = io_x[17] ? _GEN3172 : _GEN3171;
wire  _GEN3174 = io_x[75] ? _GEN3173 : _GEN3170;
wire  _GEN3175 = io_x[25] ? _GEN3174 : _GEN3167;
wire  _GEN3176 = io_x[37] ? _GEN3175 : _GEN3164;
wire  _GEN3177 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3178 = io_x[17] ? _GEN3177 : _GEN1731;
wire  _GEN3179 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3180 = io_x[17] ? _GEN3179 : _GEN1731;
wire  _GEN3181 = io_x[75] ? _GEN3180 : _GEN3178;
wire  _GEN3182 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3183 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3184 = io_x[17] ? _GEN3183 : _GEN3182;
wire  _GEN3185 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3186 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3187 = io_x[17] ? _GEN3186 : _GEN3185;
wire  _GEN3188 = io_x[75] ? _GEN3187 : _GEN3184;
wire  _GEN3189 = io_x[25] ? _GEN3188 : _GEN3181;
wire  _GEN3190 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3191 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3192 = io_x[17] ? _GEN3191 : _GEN3190;
wire  _GEN3193 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3194 = io_x[17] ? _GEN3193 : _GEN1731;
wire  _GEN3195 = io_x[75] ? _GEN3194 : _GEN3192;
wire  _GEN3196 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3197 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3198 = io_x[17] ? _GEN3197 : _GEN3196;
wire  _GEN3199 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3200 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3201 = io_x[17] ? _GEN3200 : _GEN3199;
wire  _GEN3202 = io_x[75] ? _GEN3201 : _GEN3198;
wire  _GEN3203 = io_x[25] ? _GEN3202 : _GEN3195;
wire  _GEN3204 = io_x[37] ? _GEN3203 : _GEN3189;
wire  _GEN3205 = io_x[39] ? _GEN3204 : _GEN3176;
wire  _GEN3206 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3207 = io_x[17] ? _GEN3206 : _GEN1731;
wire  _GEN3208 = io_x[75] ? _GEN1903 : _GEN3207;
wire  _GEN3209 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3210 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3211 = io_x[17] ? _GEN3210 : _GEN3209;
wire  _GEN3212 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3213 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3214 = io_x[17] ? _GEN3213 : _GEN3212;
wire  _GEN3215 = io_x[75] ? _GEN3214 : _GEN3211;
wire  _GEN3216 = io_x[25] ? _GEN3215 : _GEN3208;
wire  _GEN3217 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3218 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3219 = io_x[17] ? _GEN3218 : _GEN3217;
wire  _GEN3220 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN3221 = io_x[75] ? _GEN3220 : _GEN3219;
wire  _GEN3222 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3223 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3224 = io_x[17] ? _GEN3223 : _GEN3222;
wire  _GEN3225 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3226 = io_x[17] ? _GEN3225 : _GEN1711;
wire  _GEN3227 = io_x[75] ? _GEN3226 : _GEN3224;
wire  _GEN3228 = io_x[25] ? _GEN3227 : _GEN3221;
wire  _GEN3229 = io_x[37] ? _GEN3228 : _GEN3216;
wire  _GEN3230 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3231 = io_x[17] ? _GEN3230 : _GEN1711;
wire  _GEN3232 = io_x[75] ? _GEN1899 : _GEN3231;
wire  _GEN3233 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3234 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3235 = io_x[17] ? _GEN3234 : _GEN3233;
wire  _GEN3236 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3237 = io_x[17] ? _GEN3236 : _GEN1711;
wire  _GEN3238 = io_x[75] ? _GEN3237 : _GEN3235;
wire  _GEN3239 = io_x[25] ? _GEN3238 : _GEN3232;
wire  _GEN3240 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3241 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3242 = io_x[17] ? _GEN3241 : _GEN3240;
wire  _GEN3243 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3244 = io_x[17] ? _GEN1711 : _GEN3243;
wire  _GEN3245 = io_x[75] ? _GEN3244 : _GEN3242;
wire  _GEN3246 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3247 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3248 = io_x[17] ? _GEN3247 : _GEN3246;
wire  _GEN3249 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3250 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3251 = io_x[17] ? _GEN3250 : _GEN3249;
wire  _GEN3252 = io_x[75] ? _GEN3251 : _GEN3248;
wire  _GEN3253 = io_x[25] ? _GEN3252 : _GEN3245;
wire  _GEN3254 = io_x[37] ? _GEN3253 : _GEN3239;
wire  _GEN3255 = io_x[39] ? _GEN3254 : _GEN3229;
wire  _GEN3256 = io_x[72] ? _GEN3255 : _GEN3205;
wire  _GEN3257 = io_x[29] ? _GEN3256 : _GEN3152;
wire  _GEN3258 = io_x[18] ? _GEN3257 : _GEN3058;
wire  _GEN3259 = io_x[19] ? _GEN3258 : _GEN2892;
wire  _GEN3260 = io_x[24] ? _GEN3259 : _GEN2514;
wire  _GEN3261 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3262 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3263 = io_x[17] ? _GEN3262 : _GEN3261;
wire  _GEN3264 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3265 = io_x[17] ? _GEN3264 : _GEN1731;
wire  _GEN3266 = io_x[75] ? _GEN3265 : _GEN3263;
wire  _GEN3267 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3268 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3269 = io_x[17] ? _GEN3268 : _GEN3267;
wire  _GEN3270 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN3271 = io_x[75] ? _GEN3270 : _GEN3269;
wire  _GEN3272 = io_x[25] ? _GEN3271 : _GEN3266;
wire  _GEN3273 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3274 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3275 = io_x[17] ? _GEN3274 : _GEN3273;
wire  _GEN3276 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3277 = io_x[17] ? _GEN1731 : _GEN3276;
wire  _GEN3278 = io_x[75] ? _GEN3277 : _GEN3275;
wire  _GEN3279 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3280 = io_x[17] ? _GEN1731 : _GEN3279;
wire  _GEN3281 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3282 = io_x[17] ? _GEN1731 : _GEN3281;
wire  _GEN3283 = io_x[75] ? _GEN3282 : _GEN3280;
wire  _GEN3284 = io_x[25] ? _GEN3283 : _GEN3278;
wire  _GEN3285 = io_x[37] ? _GEN3284 : _GEN3272;
wire  _GEN3286 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3287 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3288 = io_x[17] ? _GEN3287 : _GEN3286;
wire  _GEN3289 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3290 = io_x[17] ? _GEN1731 : _GEN3289;
wire  _GEN3291 = io_x[75] ? _GEN3290 : _GEN3288;
wire  _GEN3292 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3293 = io_x[17] ? _GEN1711 : _GEN3292;
wire  _GEN3294 = io_x[75] ? _GEN1903 : _GEN3293;
wire  _GEN3295 = io_x[25] ? _GEN3294 : _GEN3291;
wire  _GEN3296 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3297 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3298 = io_x[17] ? _GEN3297 : _GEN3296;
wire  _GEN3299 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3300 = io_x[17] ? _GEN3299 : _GEN1731;
wire  _GEN3301 = io_x[75] ? _GEN3300 : _GEN3298;
wire  _GEN3302 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3303 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3304 = io_x[17] ? _GEN3303 : _GEN3302;
wire  _GEN3305 = io_x[75] ? _GEN1899 : _GEN3304;
wire  _GEN3306 = io_x[25] ? _GEN3305 : _GEN3301;
wire  _GEN3307 = io_x[37] ? _GEN3306 : _GEN3295;
wire  _GEN3308 = io_x[39] ? _GEN3307 : _GEN3285;
wire  _GEN3309 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3310 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3311 = io_x[17] ? _GEN3310 : _GEN3309;
wire  _GEN3312 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3313 = io_x[17] ? _GEN3312 : _GEN1731;
wire  _GEN3314 = io_x[75] ? _GEN3313 : _GEN3311;
wire  _GEN3315 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3316 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3317 = io_x[17] ? _GEN3316 : _GEN3315;
wire  _GEN3318 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3319 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3320 = io_x[17] ? _GEN3319 : _GEN3318;
wire  _GEN3321 = io_x[75] ? _GEN3320 : _GEN3317;
wire  _GEN3322 = io_x[25] ? _GEN3321 : _GEN3314;
wire  _GEN3323 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3324 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3325 = io_x[17] ? _GEN3324 : _GEN3323;
wire  _GEN3326 = io_x[75] ? _GEN1899 : _GEN3325;
wire  _GEN3327 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3328 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3329 = io_x[17] ? _GEN3328 : _GEN3327;
wire  _GEN3330 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3331 = io_x[17] ? _GEN1731 : _GEN3330;
wire  _GEN3332 = io_x[75] ? _GEN3331 : _GEN3329;
wire  _GEN3333 = io_x[25] ? _GEN3332 : _GEN3326;
wire  _GEN3334 = io_x[37] ? _GEN3333 : _GEN3322;
wire  _GEN3335 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3336 = io_x[17] ? _GEN1711 : _GEN3335;
wire  _GEN3337 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3338 = io_x[17] ? _GEN3337 : _GEN1731;
wire  _GEN3339 = io_x[75] ? _GEN3338 : _GEN3336;
wire  _GEN3340 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3341 = io_x[17] ? _GEN1711 : _GEN3340;
wire  _GEN3342 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3343 = io_x[17] ? _GEN3342 : _GEN1731;
wire  _GEN3344 = io_x[75] ? _GEN3343 : _GEN3341;
wire  _GEN3345 = io_x[25] ? _GEN3344 : _GEN3339;
wire  _GEN3346 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3347 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3348 = io_x[17] ? _GEN3347 : _GEN3346;
wire  _GEN3349 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3350 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3351 = io_x[17] ? _GEN3350 : _GEN3349;
wire  _GEN3352 = io_x[75] ? _GEN3351 : _GEN3348;
wire  _GEN3353 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3354 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3355 = io_x[17] ? _GEN3354 : _GEN3353;
wire  _GEN3356 = io_x[75] ? _GEN1899 : _GEN3355;
wire  _GEN3357 = io_x[25] ? _GEN3356 : _GEN3352;
wire  _GEN3358 = io_x[37] ? _GEN3357 : _GEN3345;
wire  _GEN3359 = io_x[39] ? _GEN3358 : _GEN3334;
wire  _GEN3360 = io_x[72] ? _GEN3359 : _GEN3308;
wire  _GEN3361 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3362 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3363 = io_x[17] ? _GEN3362 : _GEN3361;
wire  _GEN3364 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3365 = io_x[17] ? _GEN3364 : _GEN1731;
wire  _GEN3366 = io_x[75] ? _GEN3365 : _GEN3363;
wire  _GEN3367 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3368 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3369 = io_x[17] ? _GEN3368 : _GEN3367;
wire  _GEN3370 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3371 = io_x[17] ? _GEN1731 : _GEN3370;
wire  _GEN3372 = io_x[75] ? _GEN3371 : _GEN3369;
wire  _GEN3373 = io_x[25] ? _GEN3372 : _GEN3366;
wire  _GEN3374 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3375 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3376 = io_x[17] ? _GEN3375 : _GEN3374;
wire  _GEN3377 = io_x[75] ? _GEN1899 : _GEN3376;
wire  _GEN3378 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3379 = io_x[17] ? _GEN3378 : _GEN1731;
wire  _GEN3380 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3381 = io_x[75] ? _GEN3380 : _GEN3379;
wire  _GEN3382 = io_x[25] ? _GEN3381 : _GEN3377;
wire  _GEN3383 = io_x[37] ? _GEN3382 : _GEN3373;
wire  _GEN3384 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3385 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3386 = io_x[17] ? _GEN1711 : _GEN3385;
wire  _GEN3387 = io_x[75] ? _GEN3386 : _GEN3384;
wire  _GEN3388 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3389 = io_x[17] ? _GEN1731 : _GEN3388;
wire  _GEN3390 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3391 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3392 = io_x[17] ? _GEN3391 : _GEN3390;
wire  _GEN3393 = io_x[75] ? _GEN3392 : _GEN3389;
wire  _GEN3394 = io_x[25] ? _GEN3393 : _GEN3387;
wire  _GEN3395 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3396 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3397 = io_x[17] ? _GEN3396 : _GEN3395;
wire  _GEN3398 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3399 = io_x[17] ? _GEN1731 : _GEN3398;
wire  _GEN3400 = io_x[75] ? _GEN3399 : _GEN3397;
wire  _GEN3401 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3402 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3403 = io_x[17] ? _GEN3402 : _GEN3401;
wire  _GEN3404 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3405 = io_x[75] ? _GEN3404 : _GEN3403;
wire  _GEN3406 = io_x[25] ? _GEN3405 : _GEN3400;
wire  _GEN3407 = io_x[37] ? _GEN3406 : _GEN3394;
wire  _GEN3408 = io_x[39] ? _GEN3407 : _GEN3383;
wire  _GEN3409 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3410 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3411 = io_x[17] ? _GEN3410 : _GEN3409;
wire  _GEN3412 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3413 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3414 = io_x[17] ? _GEN3413 : _GEN3412;
wire  _GEN3415 = io_x[75] ? _GEN3414 : _GEN3411;
wire  _GEN3416 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3417 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3418 = io_x[17] ? _GEN3417 : _GEN3416;
wire  _GEN3419 = io_x[75] ? _GEN1899 : _GEN3418;
wire  _GEN3420 = io_x[25] ? _GEN3419 : _GEN3415;
wire  _GEN3421 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3422 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3423 = io_x[17] ? _GEN3422 : _GEN3421;
wire  _GEN3424 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3425 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3426 = io_x[17] ? _GEN3425 : _GEN3424;
wire  _GEN3427 = io_x[75] ? _GEN3426 : _GEN3423;
wire  _GEN3428 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3429 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3430 = io_x[17] ? _GEN3429 : _GEN3428;
wire  _GEN3431 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3432 = io_x[17] ? _GEN3431 : _GEN1731;
wire  _GEN3433 = io_x[75] ? _GEN3432 : _GEN3430;
wire  _GEN3434 = io_x[25] ? _GEN3433 : _GEN3427;
wire  _GEN3435 = io_x[37] ? _GEN3434 : _GEN3420;
wire  _GEN3436 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN3437 = io_x[75] ? _GEN3436 : _GEN1903;
wire  _GEN3438 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3439 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3440 = io_x[17] ? _GEN3439 : _GEN3438;
wire  _GEN3441 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3442 = io_x[75] ? _GEN3441 : _GEN3440;
wire  _GEN3443 = io_x[25] ? _GEN3442 : _GEN3437;
wire  _GEN3444 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3445 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3446 = io_x[17] ? _GEN3445 : _GEN3444;
wire  _GEN3447 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3448 = io_x[17] ? _GEN1731 : _GEN3447;
wire  _GEN3449 = io_x[75] ? _GEN3448 : _GEN3446;
wire  _GEN3450 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3451 = io_x[17] ? _GEN3450 : _GEN1711;
wire  _GEN3452 = io_x[75] ? _GEN1903 : _GEN3451;
wire  _GEN3453 = io_x[25] ? _GEN3452 : _GEN3449;
wire  _GEN3454 = io_x[37] ? _GEN3453 : _GEN3443;
wire  _GEN3455 = io_x[39] ? _GEN3454 : _GEN3435;
wire  _GEN3456 = io_x[72] ? _GEN3455 : _GEN3408;
wire  _GEN3457 = io_x[29] ? _GEN3456 : _GEN3360;
wire  _GEN3458 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3459 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3460 = io_x[17] ? _GEN3459 : _GEN3458;
wire  _GEN3461 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3462 = io_x[17] ? _GEN1731 : _GEN3461;
wire  _GEN3463 = io_x[75] ? _GEN3462 : _GEN3460;
wire  _GEN3464 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3465 = io_x[17] ? _GEN1711 : _GEN3464;
wire  _GEN3466 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3467 = io_x[17] ? _GEN3466 : _GEN1731;
wire  _GEN3468 = io_x[75] ? _GEN3467 : _GEN3465;
wire  _GEN3469 = io_x[25] ? _GEN3468 : _GEN3463;
wire  _GEN3470 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3471 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3472 = io_x[17] ? _GEN3471 : _GEN3470;
wire  _GEN3473 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3474 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3475 = io_x[17] ? _GEN3474 : _GEN3473;
wire  _GEN3476 = io_x[75] ? _GEN3475 : _GEN3472;
wire  _GEN3477 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3478 = io_x[17] ? _GEN3477 : _GEN1711;
wire  _GEN3479 = io_x[75] ? _GEN1903 : _GEN3478;
wire  _GEN3480 = io_x[25] ? _GEN3479 : _GEN3476;
wire  _GEN3481 = io_x[37] ? _GEN3480 : _GEN3469;
wire  _GEN3482 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3483 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3484 = io_x[17] ? _GEN3483 : _GEN3482;
wire  _GEN3485 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3486 = io_x[17] ? _GEN1731 : _GEN3485;
wire  _GEN3487 = io_x[75] ? _GEN3486 : _GEN3484;
wire  _GEN3488 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3489 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3490 = io_x[17] ? _GEN3489 : _GEN3488;
wire  _GEN3491 = io_x[75] ? _GEN1899 : _GEN3490;
wire  _GEN3492 = io_x[25] ? _GEN3491 : _GEN3487;
wire  _GEN3493 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3494 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3495 = io_x[17] ? _GEN3494 : _GEN3493;
wire  _GEN3496 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3497 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3498 = io_x[17] ? _GEN3497 : _GEN3496;
wire  _GEN3499 = io_x[75] ? _GEN3498 : _GEN3495;
wire  _GEN3500 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3501 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3502 = io_x[17] ? _GEN3501 : _GEN3500;
wire  _GEN3503 = io_x[75] ? _GEN1903 : _GEN3502;
wire  _GEN3504 = io_x[25] ? _GEN3503 : _GEN3499;
wire  _GEN3505 = io_x[37] ? _GEN3504 : _GEN3492;
wire  _GEN3506 = io_x[39] ? _GEN3505 : _GEN3481;
wire  _GEN3507 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3508 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3509 = io_x[17] ? _GEN3508 : _GEN3507;
wire  _GEN3510 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3511 = io_x[17] ? _GEN3510 : _GEN1711;
wire  _GEN3512 = io_x[75] ? _GEN3511 : _GEN3509;
wire  _GEN3513 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3514 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3515 = io_x[17] ? _GEN3514 : _GEN3513;
wire  _GEN3516 = io_x[75] ? _GEN1899 : _GEN3515;
wire  _GEN3517 = io_x[25] ? _GEN3516 : _GEN3512;
wire  _GEN3518 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3519 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3520 = io_x[17] ? _GEN3519 : _GEN3518;
wire  _GEN3521 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3522 = io_x[17] ? _GEN1711 : _GEN3521;
wire  _GEN3523 = io_x[75] ? _GEN3522 : _GEN3520;
wire  _GEN3524 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3525 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3526 = io_x[17] ? _GEN3525 : _GEN3524;
wire  _GEN3527 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3528 = io_x[75] ? _GEN3527 : _GEN3526;
wire  _GEN3529 = io_x[25] ? _GEN3528 : _GEN3523;
wire  _GEN3530 = io_x[37] ? _GEN3529 : _GEN3517;
wire  _GEN3531 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3532 = io_x[17] ? _GEN3531 : _GEN1731;
wire  _GEN3533 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3534 = io_x[17] ? _GEN3533 : _GEN1711;
wire  _GEN3535 = io_x[75] ? _GEN3534 : _GEN3532;
wire  _GEN3536 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3537 = io_x[17] ? _GEN3536 : _GEN1711;
wire  _GEN3538 = io_x[75] ? _GEN1903 : _GEN3537;
wire  _GEN3539 = io_x[25] ? _GEN3538 : _GEN3535;
wire  _GEN3540 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3541 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3542 = io_x[17] ? _GEN3541 : _GEN3540;
wire  _GEN3543 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3544 = io_x[17] ? _GEN1731 : _GEN3543;
wire  _GEN3545 = io_x[75] ? _GEN3544 : _GEN3542;
wire  _GEN3546 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3547 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3548 = io_x[17] ? _GEN3547 : _GEN3546;
wire  _GEN3549 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3550 = io_x[17] ? _GEN3549 : _GEN1711;
wire  _GEN3551 = io_x[75] ? _GEN3550 : _GEN3548;
wire  _GEN3552 = io_x[25] ? _GEN3551 : _GEN3545;
wire  _GEN3553 = io_x[37] ? _GEN3552 : _GEN3539;
wire  _GEN3554 = io_x[39] ? _GEN3553 : _GEN3530;
wire  _GEN3555 = io_x[72] ? _GEN3554 : _GEN3506;
wire  _GEN3556 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3557 = io_x[17] ? _GEN1731 : _GEN3556;
wire  _GEN3558 = io_x[75] ? _GEN1899 : _GEN3557;
wire  _GEN3559 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3560 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3561 = io_x[17] ? _GEN3560 : _GEN3559;
wire  _GEN3562 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3563 = io_x[17] ? _GEN3562 : _GEN1731;
wire  _GEN3564 = io_x[75] ? _GEN3563 : _GEN3561;
wire  _GEN3565 = io_x[25] ? _GEN3564 : _GEN3558;
wire  _GEN3566 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3567 = io_x[17] ? _GEN1731 : _GEN3566;
wire  _GEN3568 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3569 = io_x[17] ? _GEN3568 : _GEN1711;
wire  _GEN3570 = io_x[75] ? _GEN3569 : _GEN3567;
wire  _GEN3571 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3572 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3573 = io_x[17] ? _GEN3572 : _GEN3571;
wire  _GEN3574 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3575 = io_x[17] ? _GEN3574 : _GEN1731;
wire  _GEN3576 = io_x[75] ? _GEN3575 : _GEN3573;
wire  _GEN3577 = io_x[25] ? _GEN3576 : _GEN3570;
wire  _GEN3578 = io_x[37] ? _GEN3577 : _GEN3565;
wire  _GEN3579 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3580 = io_x[17] ? _GEN1731 : _GEN3579;
wire  _GEN3581 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3582 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3583 = io_x[17] ? _GEN3582 : _GEN3581;
wire  _GEN3584 = io_x[75] ? _GEN3583 : _GEN3580;
wire  _GEN3585 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3586 = io_x[17] ? _GEN3585 : _GEN1731;
wire  _GEN3587 = io_x[75] ? _GEN3586 : _GEN1903;
wire  _GEN3588 = io_x[25] ? _GEN3587 : _GEN3584;
wire  _GEN3589 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3590 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3591 = io_x[17] ? _GEN3590 : _GEN3589;
wire  _GEN3592 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3593 = io_x[17] ? _GEN3592 : _GEN1711;
wire  _GEN3594 = io_x[75] ? _GEN3593 : _GEN3591;
wire  _GEN3595 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3596 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3597 = io_x[17] ? _GEN3596 : _GEN3595;
wire  _GEN3598 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3599 = io_x[17] ? _GEN3598 : _GEN1711;
wire  _GEN3600 = io_x[75] ? _GEN3599 : _GEN3597;
wire  _GEN3601 = io_x[25] ? _GEN3600 : _GEN3594;
wire  _GEN3602 = io_x[37] ? _GEN3601 : _GEN3588;
wire  _GEN3603 = io_x[39] ? _GEN3602 : _GEN3578;
wire  _GEN3604 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3605 = io_x[17] ? _GEN1711 : _GEN3604;
wire  _GEN3606 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3607 = io_x[17] ? _GEN3606 : _GEN1731;
wire  _GEN3608 = io_x[75] ? _GEN3607 : _GEN3605;
wire  _GEN3609 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3610 = io_x[17] ? _GEN3609 : _GEN1731;
wire  _GEN3611 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3612 = io_x[17] ? _GEN1731 : _GEN3611;
wire  _GEN3613 = io_x[75] ? _GEN3612 : _GEN3610;
wire  _GEN3614 = io_x[25] ? _GEN3613 : _GEN3608;
wire  _GEN3615 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3616 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3617 = io_x[17] ? _GEN3616 : _GEN3615;
wire  _GEN3618 = io_x[75] ? _GEN1899 : _GEN3617;
wire  _GEN3619 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3620 = io_x[17] ? _GEN1731 : _GEN3619;
wire  _GEN3621 = io_x[75] ? _GEN1899 : _GEN3620;
wire  _GEN3622 = io_x[25] ? _GEN3621 : _GEN3618;
wire  _GEN3623 = io_x[37] ? _GEN3622 : _GEN3614;
wire  _GEN3624 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3625 = io_x[17] ? _GEN3624 : _GEN1731;
wire  _GEN3626 = io_x[75] ? _GEN3625 : _GEN1899;
wire  _GEN3627 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3628 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3629 = io_x[17] ? _GEN3628 : _GEN3627;
wire  _GEN3630 = io_x[75] ? _GEN3629 : _GEN1899;
wire  _GEN3631 = io_x[25] ? _GEN3630 : _GEN3626;
wire  _GEN3632 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3633 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3634 = io_x[17] ? _GEN3633 : _GEN3632;
wire  _GEN3635 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3636 = io_x[17] ? _GEN1711 : _GEN3635;
wire  _GEN3637 = io_x[75] ? _GEN3636 : _GEN3634;
wire  _GEN3638 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3639 = io_x[17] ? _GEN3638 : _GEN1731;
wire  _GEN3640 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3641 = io_x[17] ? _GEN1731 : _GEN3640;
wire  _GEN3642 = io_x[75] ? _GEN3641 : _GEN3639;
wire  _GEN3643 = io_x[25] ? _GEN3642 : _GEN3637;
wire  _GEN3644 = io_x[37] ? _GEN3643 : _GEN3631;
wire  _GEN3645 = io_x[39] ? _GEN3644 : _GEN3623;
wire  _GEN3646 = io_x[72] ? _GEN3645 : _GEN3603;
wire  _GEN3647 = io_x[29] ? _GEN3646 : _GEN3555;
wire  _GEN3648 = io_x[18] ? _GEN3647 : _GEN3457;
wire  _GEN3649 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3650 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3651 = io_x[17] ? _GEN3650 : _GEN3649;
wire  _GEN3652 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3653 = io_x[17] ? _GEN1731 : _GEN3652;
wire  _GEN3654 = io_x[75] ? _GEN3653 : _GEN3651;
wire  _GEN3655 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3656 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3657 = io_x[17] ? _GEN3656 : _GEN3655;
wire  _GEN3658 = io_x[75] ? _GEN1899 : _GEN3657;
wire  _GEN3659 = io_x[25] ? _GEN3658 : _GEN3654;
wire  _GEN3660 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN3661 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3662 = io_x[17] ? _GEN1731 : _GEN3661;
wire  _GEN3663 = io_x[75] ? _GEN3662 : _GEN3660;
wire  _GEN3664 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3665 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3666 = io_x[17] ? _GEN3665 : _GEN3664;
wire  _GEN3667 = io_x[75] ? _GEN3666 : _GEN1903;
wire  _GEN3668 = io_x[25] ? _GEN3667 : _GEN3663;
wire  _GEN3669 = io_x[37] ? _GEN3668 : _GEN3659;
wire  _GEN3670 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3671 = io_x[17] ? _GEN1731 : _GEN3670;
wire  _GEN3672 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3673 = io_x[17] ? _GEN1731 : _GEN3672;
wire  _GEN3674 = io_x[75] ? _GEN3673 : _GEN3671;
wire  _GEN3675 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3676 = io_x[75] ? _GEN1899 : _GEN3675;
wire  _GEN3677 = io_x[25] ? _GEN3676 : _GEN3674;
wire  _GEN3678 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3679 = io_x[17] ? _GEN1711 : _GEN3678;
wire  _GEN3680 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3681 = io_x[75] ? _GEN3680 : _GEN3679;
wire  _GEN3682 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3683 = io_x[17] ? _GEN1731 : _GEN3682;
wire  _GEN3684 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3685 = io_x[17] ? _GEN3684 : _GEN1731;
wire  _GEN3686 = io_x[75] ? _GEN3685 : _GEN3683;
wire  _GEN3687 = io_x[25] ? _GEN3686 : _GEN3681;
wire  _GEN3688 = io_x[37] ? _GEN3687 : _GEN3677;
wire  _GEN3689 = io_x[39] ? _GEN3688 : _GEN3669;
wire  _GEN3690 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3691 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3692 = io_x[17] ? _GEN3691 : _GEN3690;
wire  _GEN3693 = io_x[75] ? _GEN1903 : _GEN3692;
wire  _GEN3694 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3695 = io_x[17] ? _GEN1731 : _GEN3694;
wire  _GEN3696 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3697 = io_x[17] ? _GEN1731 : _GEN3696;
wire  _GEN3698 = io_x[75] ? _GEN3697 : _GEN3695;
wire  _GEN3699 = io_x[25] ? _GEN3698 : _GEN3693;
wire  _GEN3700 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3701 = io_x[17] ? _GEN1711 : _GEN3700;
wire  _GEN3702 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3703 = io_x[75] ? _GEN3702 : _GEN3701;
wire  _GEN3704 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3705 = io_x[17] ? _GEN1731 : _GEN3704;
wire  _GEN3706 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3707 = io_x[17] ? _GEN3706 : _GEN1731;
wire  _GEN3708 = io_x[75] ? _GEN3707 : _GEN3705;
wire  _GEN3709 = io_x[25] ? _GEN3708 : _GEN3703;
wire  _GEN3710 = io_x[37] ? _GEN3709 : _GEN3699;
wire  _GEN3711 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3712 = io_x[17] ? _GEN1731 : _GEN3711;
wire  _GEN3713 = io_x[75] ? _GEN1903 : _GEN3712;
wire  _GEN3714 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3715 = io_x[17] ? _GEN3714 : _GEN1711;
wire  _GEN3716 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3717 = io_x[75] ? _GEN3716 : _GEN3715;
wire  _GEN3718 = io_x[25] ? _GEN3717 : _GEN3713;
wire  _GEN3719 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3720 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3721 = io_x[17] ? _GEN3720 : _GEN3719;
wire  _GEN3722 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3723 = io_x[17] ? _GEN1731 : _GEN3722;
wire  _GEN3724 = io_x[75] ? _GEN3723 : _GEN3721;
wire  _GEN3725 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3726 = io_x[17] ? _GEN1731 : _GEN3725;
wire  _GEN3727 = io_x[75] ? _GEN1899 : _GEN3726;
wire  _GEN3728 = io_x[25] ? _GEN3727 : _GEN3724;
wire  _GEN3729 = io_x[37] ? _GEN3728 : _GEN3718;
wire  _GEN3730 = io_x[39] ? _GEN3729 : _GEN3710;
wire  _GEN3731 = io_x[72] ? _GEN3730 : _GEN3689;
wire  _GEN3732 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3733 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3734 = io_x[17] ? _GEN3733 : _GEN3732;
wire  _GEN3735 = io_x[75] ? _GEN1899 : _GEN3734;
wire  _GEN3736 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3737 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3738 = io_x[17] ? _GEN3737 : _GEN3736;
wire  _GEN3739 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3740 = io_x[17] ? _GEN3739 : _GEN1731;
wire  _GEN3741 = io_x[75] ? _GEN3740 : _GEN3738;
wire  _GEN3742 = io_x[25] ? _GEN3741 : _GEN3735;
wire  _GEN3743 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3744 = io_x[17] ? _GEN1731 : _GEN3743;
wire  _GEN3745 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3746 = io_x[17] ? _GEN1731 : _GEN3745;
wire  _GEN3747 = io_x[75] ? _GEN3746 : _GEN3744;
wire  _GEN3748 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN3749 = io_x[75] ? _GEN1899 : _GEN3748;
wire  _GEN3750 = io_x[25] ? _GEN3749 : _GEN3747;
wire  _GEN3751 = io_x[37] ? _GEN3750 : _GEN3742;
wire  _GEN3752 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3753 = io_x[17] ? _GEN1731 : _GEN3752;
wire  _GEN3754 = io_x[75] ? _GEN3753 : _GEN1903;
wire  _GEN3755 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN3756 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3757 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3758 = io_x[17] ? _GEN3757 : _GEN3756;
wire  _GEN3759 = io_x[75] ? _GEN3758 : _GEN3755;
wire  _GEN3760 = io_x[25] ? _GEN3759 : _GEN3754;
wire  _GEN3761 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3762 = io_x[17] ? _GEN1711 : _GEN3761;
wire  _GEN3763 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3764 = io_x[17] ? _GEN1731 : _GEN3763;
wire  _GEN3765 = io_x[75] ? _GEN3764 : _GEN3762;
wire  _GEN3766 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3767 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3768 = io_x[17] ? _GEN3767 : _GEN3766;
wire  _GEN3769 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3770 = io_x[75] ? _GEN3769 : _GEN3768;
wire  _GEN3771 = io_x[25] ? _GEN3770 : _GEN3765;
wire  _GEN3772 = io_x[37] ? _GEN3771 : _GEN3760;
wire  _GEN3773 = io_x[39] ? _GEN3772 : _GEN3751;
wire  _GEN3774 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3775 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3776 = io_x[17] ? _GEN3775 : _GEN3774;
wire  _GEN3777 = io_x[75] ? _GEN1903 : _GEN3776;
wire  _GEN3778 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN3779 = io_x[25] ? _GEN3778 : _GEN3777;
wire  _GEN3780 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3781 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3782 = io_x[17] ? _GEN3781 : _GEN3780;
wire  _GEN3783 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3784 = io_x[17] ? _GEN1731 : _GEN3783;
wire  _GEN3785 = io_x[75] ? _GEN3784 : _GEN3782;
wire  _GEN3786 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3787 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3788 = io_x[17] ? _GEN3787 : _GEN3786;
wire  _GEN3789 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3790 = io_x[17] ? _GEN3789 : _GEN1731;
wire  _GEN3791 = io_x[75] ? _GEN3790 : _GEN3788;
wire  _GEN3792 = io_x[25] ? _GEN3791 : _GEN3785;
wire  _GEN3793 = io_x[37] ? _GEN3792 : _GEN3779;
wire  _GEN3794 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3795 = io_x[17] ? _GEN3794 : _GEN1711;
wire  _GEN3796 = io_x[75] ? _GEN1903 : _GEN3795;
wire  _GEN3797 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3798 = io_x[17] ? _GEN3797 : _GEN1731;
wire  _GEN3799 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3800 = io_x[17] ? _GEN3799 : _GEN1731;
wire  _GEN3801 = io_x[75] ? _GEN3800 : _GEN3798;
wire  _GEN3802 = io_x[25] ? _GEN3801 : _GEN3796;
wire  _GEN3803 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3804 = io_x[17] ? _GEN1731 : _GEN3803;
wire  _GEN3805 = io_x[75] ? _GEN1903 : _GEN3804;
wire  _GEN3806 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3807 = io_x[17] ? _GEN1711 : _GEN3806;
wire  _GEN3808 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3809 = io_x[17] ? _GEN3808 : _GEN1731;
wire  _GEN3810 = io_x[75] ? _GEN3809 : _GEN3807;
wire  _GEN3811 = io_x[25] ? _GEN3810 : _GEN3805;
wire  _GEN3812 = io_x[37] ? _GEN3811 : _GEN3802;
wire  _GEN3813 = io_x[39] ? _GEN3812 : _GEN3793;
wire  _GEN3814 = io_x[72] ? _GEN3813 : _GEN3773;
wire  _GEN3815 = io_x[29] ? _GEN3814 : _GEN3731;
wire  _GEN3816 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3817 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3818 = io_x[17] ? _GEN3817 : _GEN3816;
wire  _GEN3819 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3820 = io_x[17] ? _GEN3819 : _GEN1731;
wire  _GEN3821 = io_x[75] ? _GEN3820 : _GEN3818;
wire  _GEN3822 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3823 = io_x[17] ? _GEN3822 : _GEN1711;
wire  _GEN3824 = io_x[75] ? _GEN1903 : _GEN3823;
wire  _GEN3825 = io_x[25] ? _GEN3824 : _GEN3821;
wire  _GEN3826 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3827 = io_x[17] ? _GEN1711 : _GEN3826;
wire  _GEN3828 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3829 = io_x[17] ? _GEN3828 : _GEN1731;
wire  _GEN3830 = io_x[75] ? _GEN3829 : _GEN3827;
wire  _GEN3831 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3832 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3833 = io_x[17] ? _GEN3832 : _GEN3831;
wire  _GEN3834 = io_x[75] ? _GEN1903 : _GEN3833;
wire  _GEN3835 = io_x[25] ? _GEN3834 : _GEN3830;
wire  _GEN3836 = io_x[37] ? _GEN3835 : _GEN3825;
wire  _GEN3837 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3838 = io_x[17] ? _GEN3837 : _GEN1731;
wire  _GEN3839 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3840 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3841 = io_x[17] ? _GEN3840 : _GEN3839;
wire  _GEN3842 = io_x[75] ? _GEN3841 : _GEN3838;
wire  _GEN3843 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3844 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3845 = io_x[17] ? _GEN1711 : _GEN3844;
wire  _GEN3846 = io_x[75] ? _GEN3845 : _GEN3843;
wire  _GEN3847 = io_x[25] ? _GEN3846 : _GEN3842;
wire  _GEN3848 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3849 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3850 = io_x[17] ? _GEN3849 : _GEN3848;
wire  _GEN3851 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3852 = io_x[17] ? _GEN3851 : _GEN1731;
wire  _GEN3853 = io_x[75] ? _GEN3852 : _GEN3850;
wire  _GEN3854 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3855 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3856 = io_x[17] ? _GEN3855 : _GEN3854;
wire  _GEN3857 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3858 = io_x[17] ? _GEN3857 : _GEN1731;
wire  _GEN3859 = io_x[75] ? _GEN3858 : _GEN3856;
wire  _GEN3860 = io_x[25] ? _GEN3859 : _GEN3853;
wire  _GEN3861 = io_x[37] ? _GEN3860 : _GEN3847;
wire  _GEN3862 = io_x[39] ? _GEN3861 : _GEN3836;
wire  _GEN3863 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3864 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3865 = io_x[17] ? _GEN3864 : _GEN3863;
wire  _GEN3866 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3867 = io_x[17] ? _GEN3866 : _GEN1711;
wire  _GEN3868 = io_x[75] ? _GEN3867 : _GEN3865;
wire  _GEN3869 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3870 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3871 = io_x[17] ? _GEN3870 : _GEN3869;
wire  _GEN3872 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN3873 = io_x[75] ? _GEN3872 : _GEN3871;
wire  _GEN3874 = io_x[25] ? _GEN3873 : _GEN3868;
wire  _GEN3875 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3876 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3877 = io_x[17] ? _GEN3876 : _GEN3875;
wire  _GEN3878 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3879 = io_x[17] ? _GEN3878 : _GEN1711;
wire  _GEN3880 = io_x[75] ? _GEN3879 : _GEN3877;
wire  _GEN3881 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3882 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3883 = io_x[17] ? _GEN3882 : _GEN3881;
wire  _GEN3884 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN3885 = io_x[75] ? _GEN3884 : _GEN3883;
wire  _GEN3886 = io_x[25] ? _GEN3885 : _GEN3880;
wire  _GEN3887 = io_x[37] ? _GEN3886 : _GEN3874;
wire  _GEN3888 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3889 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3890 = io_x[17] ? _GEN3889 : _GEN3888;
wire  _GEN3891 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3892 = io_x[75] ? _GEN3891 : _GEN3890;
wire  _GEN3893 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN3894 = io_x[75] ? _GEN1903 : _GEN3893;
wire  _GEN3895 = io_x[25] ? _GEN3894 : _GEN3892;
wire  _GEN3896 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3897 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3898 = io_x[17] ? _GEN3897 : _GEN3896;
wire  _GEN3899 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3900 = io_x[17] ? _GEN1731 : _GEN3899;
wire  _GEN3901 = io_x[75] ? _GEN3900 : _GEN3898;
wire  _GEN3902 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3903 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3904 = io_x[17] ? _GEN3903 : _GEN3902;
wire  _GEN3905 = io_x[75] ? _GEN1903 : _GEN3904;
wire  _GEN3906 = io_x[25] ? _GEN3905 : _GEN3901;
wire  _GEN3907 = io_x[37] ? _GEN3906 : _GEN3895;
wire  _GEN3908 = io_x[39] ? _GEN3907 : _GEN3887;
wire  _GEN3909 = io_x[72] ? _GEN3908 : _GEN3862;
wire  _GEN3910 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3911 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3912 = io_x[17] ? _GEN3911 : _GEN3910;
wire  _GEN3913 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3914 = io_x[17] ? _GEN3913 : _GEN1711;
wire  _GEN3915 = io_x[75] ? _GEN3914 : _GEN3912;
wire  _GEN3916 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3917 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3918 = io_x[17] ? _GEN3917 : _GEN3916;
wire  _GEN3919 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3920 = io_x[17] ? _GEN3919 : _GEN1711;
wire  _GEN3921 = io_x[75] ? _GEN3920 : _GEN3918;
wire  _GEN3922 = io_x[25] ? _GEN3921 : _GEN3915;
wire  _GEN3923 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3924 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3925 = io_x[17] ? _GEN3924 : _GEN3923;
wire  _GEN3926 = io_x[75] ? _GEN1903 : _GEN3925;
wire  _GEN3927 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3928 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3929 = io_x[17] ? _GEN3928 : _GEN3927;
wire  _GEN3930 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3931 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3932 = io_x[17] ? _GEN3931 : _GEN3930;
wire  _GEN3933 = io_x[75] ? _GEN3932 : _GEN3929;
wire  _GEN3934 = io_x[25] ? _GEN3933 : _GEN3926;
wire  _GEN3935 = io_x[37] ? _GEN3934 : _GEN3922;
wire  _GEN3936 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3937 = io_x[17] ? _GEN3936 : _GEN1711;
wire  _GEN3938 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3939 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3940 = io_x[17] ? _GEN3939 : _GEN3938;
wire  _GEN3941 = io_x[75] ? _GEN3940 : _GEN3937;
wire  _GEN3942 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3943 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3944 = io_x[17] ? _GEN3943 : _GEN3942;
wire  _GEN3945 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3946 = io_x[17] ? _GEN3945 : _GEN1711;
wire  _GEN3947 = io_x[75] ? _GEN3946 : _GEN3944;
wire  _GEN3948 = io_x[25] ? _GEN3947 : _GEN3941;
wire  _GEN3949 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3950 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3951 = io_x[17] ? _GEN3950 : _GEN3949;
wire  _GEN3952 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3953 = io_x[17] ? _GEN3952 : _GEN1711;
wire  _GEN3954 = io_x[75] ? _GEN3953 : _GEN3951;
wire  _GEN3955 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3956 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3957 = io_x[17] ? _GEN3956 : _GEN3955;
wire  _GEN3958 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3959 = io_x[17] ? _GEN3958 : _GEN1731;
wire  _GEN3960 = io_x[75] ? _GEN3959 : _GEN3957;
wire  _GEN3961 = io_x[25] ? _GEN3960 : _GEN3954;
wire  _GEN3962 = io_x[37] ? _GEN3961 : _GEN3948;
wire  _GEN3963 = io_x[39] ? _GEN3962 : _GEN3935;
wire  _GEN3964 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3965 = io_x[17] ? _GEN3964 : _GEN1711;
wire  _GEN3966 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3967 = io_x[17] ? _GEN3966 : _GEN1731;
wire  _GEN3968 = io_x[75] ? _GEN3967 : _GEN3965;
wire  _GEN3969 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3970 = io_x[17] ? _GEN3969 : _GEN1711;
wire  _GEN3971 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3972 = io_x[17] ? _GEN3971 : _GEN1731;
wire  _GEN3973 = io_x[75] ? _GEN3972 : _GEN3970;
wire  _GEN3974 = io_x[25] ? _GEN3973 : _GEN3968;
wire  _GEN3975 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3976 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3977 = io_x[17] ? _GEN3976 : _GEN3975;
wire  _GEN3978 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3979 = io_x[17] ? _GEN3978 : _GEN1731;
wire  _GEN3980 = io_x[75] ? _GEN3979 : _GEN3977;
wire  _GEN3981 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3982 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3983 = io_x[17] ? _GEN3982 : _GEN3981;
wire  _GEN3984 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3985 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3986 = io_x[17] ? _GEN3985 : _GEN3984;
wire  _GEN3987 = io_x[75] ? _GEN3986 : _GEN3983;
wire  _GEN3988 = io_x[25] ? _GEN3987 : _GEN3980;
wire  _GEN3989 = io_x[37] ? _GEN3988 : _GEN3974;
wire  _GEN3990 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3991 = io_x[17] ? _GEN3990 : _GEN1711;
wire  _GEN3992 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN3993 = io_x[75] ? _GEN3992 : _GEN3991;
wire  _GEN3994 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN3995 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3996 = io_x[17] ? _GEN3995 : _GEN3994;
wire  _GEN3997 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN3998 = io_x[17] ? _GEN1731 : _GEN3997;
wire  _GEN3999 = io_x[75] ? _GEN3998 : _GEN3996;
wire  _GEN4000 = io_x[25] ? _GEN3999 : _GEN3993;
wire  _GEN4001 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4002 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4003 = io_x[17] ? _GEN4002 : _GEN4001;
wire  _GEN4004 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4005 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4006 = io_x[17] ? _GEN4005 : _GEN4004;
wire  _GEN4007 = io_x[75] ? _GEN4006 : _GEN4003;
wire  _GEN4008 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4009 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4010 = io_x[17] ? _GEN4009 : _GEN4008;
wire  _GEN4011 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4012 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4013 = io_x[17] ? _GEN4012 : _GEN4011;
wire  _GEN4014 = io_x[75] ? _GEN4013 : _GEN4010;
wire  _GEN4015 = io_x[25] ? _GEN4014 : _GEN4007;
wire  _GEN4016 = io_x[37] ? _GEN4015 : _GEN4000;
wire  _GEN4017 = io_x[39] ? _GEN4016 : _GEN3989;
wire  _GEN4018 = io_x[72] ? _GEN4017 : _GEN3963;
wire  _GEN4019 = io_x[29] ? _GEN4018 : _GEN3909;
wire  _GEN4020 = io_x[18] ? _GEN4019 : _GEN3815;
wire  _GEN4021 = io_x[19] ? _GEN4020 : _GEN3648;
wire  _GEN4022 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4023 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4024 = io_x[17] ? _GEN4023 : _GEN4022;
wire  _GEN4025 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN4026 = io_x[75] ? _GEN4025 : _GEN4024;
wire  _GEN4027 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4028 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4029 = io_x[17] ? _GEN4028 : _GEN4027;
wire  _GEN4030 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4031 = io_x[17] ? _GEN1731 : _GEN4030;
wire  _GEN4032 = io_x[75] ? _GEN4031 : _GEN4029;
wire  _GEN4033 = io_x[25] ? _GEN4032 : _GEN4026;
wire  _GEN4034 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4035 = io_x[17] ? _GEN4034 : _GEN1731;
wire  _GEN4036 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4037 = io_x[17] ? _GEN1731 : _GEN4036;
wire  _GEN4038 = io_x[75] ? _GEN4037 : _GEN4035;
wire  _GEN4039 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4040 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4041 = io_x[17] ? _GEN4040 : _GEN4039;
wire  _GEN4042 = io_x[75] ? _GEN1903 : _GEN4041;
wire  _GEN4043 = io_x[25] ? _GEN4042 : _GEN4038;
wire  _GEN4044 = io_x[37] ? _GEN4043 : _GEN4033;
wire  _GEN4045 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4046 = io_x[17] ? _GEN1731 : _GEN4045;
wire  _GEN4047 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4048 = io_x[17] ? _GEN1731 : _GEN4047;
wire  _GEN4049 = io_x[75] ? _GEN4048 : _GEN4046;
wire  _GEN4050 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4051 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4052 = io_x[17] ? _GEN4051 : _GEN4050;
wire  _GEN4053 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN4054 = io_x[75] ? _GEN4053 : _GEN4052;
wire  _GEN4055 = io_x[25] ? _GEN4054 : _GEN4049;
wire  _GEN4056 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4057 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4058 = io_x[17] ? _GEN4057 : _GEN4056;
wire  _GEN4059 = io_x[75] ? _GEN1899 : _GEN4058;
wire  _GEN4060 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4061 = io_x[17] ? _GEN4060 : _GEN1711;
wire  _GEN4062 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4063 = io_x[17] ? _GEN1731 : _GEN4062;
wire  _GEN4064 = io_x[75] ? _GEN4063 : _GEN4061;
wire  _GEN4065 = io_x[25] ? _GEN4064 : _GEN4059;
wire  _GEN4066 = io_x[37] ? _GEN4065 : _GEN4055;
wire  _GEN4067 = io_x[39] ? _GEN4066 : _GEN4044;
wire  _GEN4068 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4069 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4070 = io_x[17] ? _GEN4069 : _GEN4068;
wire  _GEN4071 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4072 = io_x[17] ? _GEN1731 : _GEN4071;
wire  _GEN4073 = io_x[75] ? _GEN4072 : _GEN4070;
wire  _GEN4074 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4075 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4076 = io_x[17] ? _GEN4075 : _GEN4074;
wire  _GEN4077 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4078 = io_x[17] ? _GEN4077 : _GEN1711;
wire  _GEN4079 = io_x[75] ? _GEN4078 : _GEN4076;
wire  _GEN4080 = io_x[25] ? _GEN4079 : _GEN4073;
wire  _GEN4081 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4082 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4083 = io_x[17] ? _GEN4082 : _GEN4081;
wire  _GEN4084 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4085 = io_x[17] ? _GEN1711 : _GEN4084;
wire  _GEN4086 = io_x[75] ? _GEN4085 : _GEN4083;
wire  _GEN4087 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4088 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4089 = io_x[17] ? _GEN4088 : _GEN4087;
wire  _GEN4090 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN4091 = io_x[75] ? _GEN4090 : _GEN4089;
wire  _GEN4092 = io_x[25] ? _GEN4091 : _GEN4086;
wire  _GEN4093 = io_x[37] ? _GEN4092 : _GEN4080;
wire  _GEN4094 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN4095 = io_x[75] ? _GEN1899 : _GEN4094;
wire  _GEN4096 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4097 = io_x[17] ? _GEN1731 : _GEN4096;
wire  _GEN4098 = io_x[75] ? _GEN1903 : _GEN4097;
wire  _GEN4099 = io_x[25] ? _GEN4098 : _GEN4095;
wire  _GEN4100 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4101 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4102 = io_x[17] ? _GEN4101 : _GEN4100;
wire  _GEN4103 = io_x[75] ? _GEN1903 : _GEN4102;
wire  _GEN4104 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4105 = io_x[17] ? _GEN1711 : _GEN4104;
wire  _GEN4106 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4107 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4108 = io_x[17] ? _GEN4107 : _GEN4106;
wire  _GEN4109 = io_x[75] ? _GEN4108 : _GEN4105;
wire  _GEN4110 = io_x[25] ? _GEN4109 : _GEN4103;
wire  _GEN4111 = io_x[37] ? _GEN4110 : _GEN4099;
wire  _GEN4112 = io_x[39] ? _GEN4111 : _GEN4093;
wire  _GEN4113 = io_x[72] ? _GEN4112 : _GEN4067;
wire  _GEN4114 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4115 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4116 = io_x[17] ? _GEN4115 : _GEN4114;
wire  _GEN4117 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4118 = io_x[17] ? _GEN1711 : _GEN4117;
wire  _GEN4119 = io_x[75] ? _GEN4118 : _GEN4116;
wire  _GEN4120 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4121 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4122 = io_x[17] ? _GEN4121 : _GEN4120;
wire  _GEN4123 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4124 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4125 = io_x[17] ? _GEN4124 : _GEN4123;
wire  _GEN4126 = io_x[75] ? _GEN4125 : _GEN4122;
wire  _GEN4127 = io_x[25] ? _GEN4126 : _GEN4119;
wire  _GEN4128 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4129 = io_x[17] ? _GEN1731 : _GEN4128;
wire  _GEN4130 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4131 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4132 = io_x[17] ? _GEN4131 : _GEN4130;
wire  _GEN4133 = io_x[75] ? _GEN4132 : _GEN4129;
wire  _GEN4134 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4135 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4136 = io_x[17] ? _GEN4135 : _GEN4134;
wire  _GEN4137 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4138 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4139 = io_x[17] ? _GEN4138 : _GEN4137;
wire  _GEN4140 = io_x[75] ? _GEN4139 : _GEN4136;
wire  _GEN4141 = io_x[25] ? _GEN4140 : _GEN4133;
wire  _GEN4142 = io_x[37] ? _GEN4141 : _GEN4127;
wire  _GEN4143 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4144 = io_x[17] ? _GEN1731 : _GEN4143;
wire  _GEN4145 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4146 = io_x[17] ? _GEN1711 : _GEN4145;
wire  _GEN4147 = io_x[75] ? _GEN4146 : _GEN4144;
wire  _GEN4148 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4149 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4150 = io_x[17] ? _GEN4149 : _GEN4148;
wire  _GEN4151 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4152 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4153 = io_x[17] ? _GEN4152 : _GEN4151;
wire  _GEN4154 = io_x[75] ? _GEN4153 : _GEN4150;
wire  _GEN4155 = io_x[25] ? _GEN4154 : _GEN4147;
wire  _GEN4156 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4157 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4158 = io_x[17] ? _GEN4157 : _GEN4156;
wire  _GEN4159 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4160 = io_x[17] ? _GEN1731 : _GEN4159;
wire  _GEN4161 = io_x[75] ? _GEN4160 : _GEN4158;
wire  _GEN4162 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4163 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4164 = io_x[17] ? _GEN4163 : _GEN4162;
wire  _GEN4165 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4166 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4167 = io_x[17] ? _GEN4166 : _GEN4165;
wire  _GEN4168 = io_x[75] ? _GEN4167 : _GEN4164;
wire  _GEN4169 = io_x[25] ? _GEN4168 : _GEN4161;
wire  _GEN4170 = io_x[37] ? _GEN4169 : _GEN4155;
wire  _GEN4171 = io_x[39] ? _GEN4170 : _GEN4142;
wire  _GEN4172 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4173 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4174 = io_x[17] ? _GEN4173 : _GEN4172;
wire  _GEN4175 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4176 = io_x[17] ? _GEN1731 : _GEN4175;
wire  _GEN4177 = io_x[75] ? _GEN4176 : _GEN4174;
wire  _GEN4178 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4179 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4180 = io_x[17] ? _GEN4179 : _GEN4178;
wire  _GEN4181 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4182 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4183 = io_x[17] ? _GEN4182 : _GEN4181;
wire  _GEN4184 = io_x[75] ? _GEN4183 : _GEN4180;
wire  _GEN4185 = io_x[25] ? _GEN4184 : _GEN4177;
wire  _GEN4186 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4187 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4188 = io_x[17] ? _GEN4187 : _GEN4186;
wire  _GEN4189 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4190 = io_x[17] ? _GEN1731 : _GEN4189;
wire  _GEN4191 = io_x[75] ? _GEN4190 : _GEN4188;
wire  _GEN4192 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4193 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4194 = io_x[17] ? _GEN4193 : _GEN4192;
wire  _GEN4195 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4196 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4197 = io_x[17] ? _GEN4196 : _GEN4195;
wire  _GEN4198 = io_x[75] ? _GEN4197 : _GEN4194;
wire  _GEN4199 = io_x[25] ? _GEN4198 : _GEN4191;
wire  _GEN4200 = io_x[37] ? _GEN4199 : _GEN4185;
wire  _GEN4201 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4202 = io_x[17] ? _GEN1711 : _GEN4201;
wire  _GEN4203 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4204 = io_x[17] ? _GEN1711 : _GEN4203;
wire  _GEN4205 = io_x[75] ? _GEN4204 : _GEN4202;
wire  _GEN4206 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4207 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4208 = io_x[17] ? _GEN4207 : _GEN4206;
wire  _GEN4209 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4210 = io_x[17] ? _GEN1731 : _GEN4209;
wire  _GEN4211 = io_x[75] ? _GEN4210 : _GEN4208;
wire  _GEN4212 = io_x[25] ? _GEN4211 : _GEN4205;
wire  _GEN4213 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4214 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4215 = io_x[17] ? _GEN4214 : _GEN4213;
wire  _GEN4216 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4217 = io_x[17] ? _GEN1711 : _GEN4216;
wire  _GEN4218 = io_x[75] ? _GEN4217 : _GEN4215;
wire  _GEN4219 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4220 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4221 = io_x[17] ? _GEN4220 : _GEN4219;
wire  _GEN4222 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4223 = io_x[17] ? _GEN1731 : _GEN4222;
wire  _GEN4224 = io_x[75] ? _GEN4223 : _GEN4221;
wire  _GEN4225 = io_x[25] ? _GEN4224 : _GEN4218;
wire  _GEN4226 = io_x[37] ? _GEN4225 : _GEN4212;
wire  _GEN4227 = io_x[39] ? _GEN4226 : _GEN4200;
wire  _GEN4228 = io_x[72] ? _GEN4227 : _GEN4171;
wire  _GEN4229 = io_x[29] ? _GEN4228 : _GEN4113;
wire  _GEN4230 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4231 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4232 = io_x[17] ? _GEN4231 : _GEN4230;
wire  _GEN4233 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4234 = io_x[17] ? _GEN4233 : _GEN1731;
wire  _GEN4235 = io_x[75] ? _GEN4234 : _GEN4232;
wire  _GEN4236 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4237 = io_x[17] ? _GEN4236 : _GEN1711;
wire  _GEN4238 = io_x[75] ? _GEN1903 : _GEN4237;
wire  _GEN4239 = io_x[25] ? _GEN4238 : _GEN4235;
wire  _GEN4240 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4241 = io_x[17] ? _GEN4240 : _GEN1731;
wire  _GEN4242 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4243 = io_x[17] ? _GEN4242 : _GEN1731;
wire  _GEN4244 = io_x[75] ? _GEN4243 : _GEN4241;
wire  _GEN4245 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4246 = io_x[17] ? _GEN4245 : _GEN1711;
wire  _GEN4247 = io_x[75] ? _GEN1903 : _GEN4246;
wire  _GEN4248 = io_x[25] ? _GEN4247 : _GEN4244;
wire  _GEN4249 = io_x[37] ? _GEN4248 : _GEN4239;
wire  _GEN4250 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4251 = io_x[17] ? _GEN1711 : _GEN4250;
wire  _GEN4252 = io_x[75] ? _GEN4251 : _GEN1899;
wire  _GEN4253 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4254 = io_x[17] ? _GEN4253 : _GEN1731;
wire  _GEN4255 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4256 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4257 = io_x[17] ? _GEN4256 : _GEN4255;
wire  _GEN4258 = io_x[75] ? _GEN4257 : _GEN4254;
wire  _GEN4259 = io_x[25] ? _GEN4258 : _GEN4252;
wire  _GEN4260 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4261 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4262 = io_x[17] ? _GEN4261 : _GEN4260;
wire  _GEN4263 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4264 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4265 = io_x[17] ? _GEN4264 : _GEN4263;
wire  _GEN4266 = io_x[75] ? _GEN4265 : _GEN4262;
wire  _GEN4267 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4268 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4269 = io_x[17] ? _GEN4268 : _GEN4267;
wire  _GEN4270 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4271 = io_x[17] ? _GEN4270 : _GEN1731;
wire  _GEN4272 = io_x[75] ? _GEN4271 : _GEN4269;
wire  _GEN4273 = io_x[25] ? _GEN4272 : _GEN4266;
wire  _GEN4274 = io_x[37] ? _GEN4273 : _GEN4259;
wire  _GEN4275 = io_x[39] ? _GEN4274 : _GEN4249;
wire  _GEN4276 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN4277 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4278 = io_x[17] ? _GEN4277 : _GEN1731;
wire  _GEN4279 = io_x[75] ? _GEN4278 : _GEN4276;
wire  _GEN4280 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4281 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4282 = io_x[17] ? _GEN4281 : _GEN4280;
wire  _GEN4283 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4284 = io_x[17] ? _GEN4283 : _GEN1731;
wire  _GEN4285 = io_x[75] ? _GEN4284 : _GEN4282;
wire  _GEN4286 = io_x[25] ? _GEN4285 : _GEN4279;
wire  _GEN4287 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4288 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4289 = io_x[17] ? _GEN4288 : _GEN4287;
wire  _GEN4290 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4291 = io_x[17] ? _GEN4290 : _GEN1731;
wire  _GEN4292 = io_x[75] ? _GEN4291 : _GEN4289;
wire  _GEN4293 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4294 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4295 = io_x[17] ? _GEN4294 : _GEN4293;
wire  _GEN4296 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4297 = io_x[17] ? _GEN4296 : _GEN1711;
wire  _GEN4298 = io_x[75] ? _GEN4297 : _GEN4295;
wire  _GEN4299 = io_x[25] ? _GEN4298 : _GEN4292;
wire  _GEN4300 = io_x[37] ? _GEN4299 : _GEN4286;
wire  _GEN4301 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN4302 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4303 = io_x[17] ? _GEN4302 : _GEN1731;
wire  _GEN4304 = io_x[75] ? _GEN4303 : _GEN4301;
wire  _GEN4305 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4306 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4307 = io_x[17] ? _GEN4306 : _GEN4305;
wire  _GEN4308 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4309 = io_x[17] ? _GEN4308 : _GEN1731;
wire  _GEN4310 = io_x[75] ? _GEN4309 : _GEN4307;
wire  _GEN4311 = io_x[25] ? _GEN4310 : _GEN4304;
wire  _GEN4312 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4313 = io_x[17] ? _GEN4312 : _GEN1711;
wire  _GEN4314 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4315 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4316 = io_x[17] ? _GEN4315 : _GEN4314;
wire  _GEN4317 = io_x[75] ? _GEN4316 : _GEN4313;
wire  _GEN4318 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4319 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4320 = io_x[17] ? _GEN4319 : _GEN4318;
wire  _GEN4321 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN4322 = io_x[75] ? _GEN4321 : _GEN4320;
wire  _GEN4323 = io_x[25] ? _GEN4322 : _GEN4317;
wire  _GEN4324 = io_x[37] ? _GEN4323 : _GEN4311;
wire  _GEN4325 = io_x[39] ? _GEN4324 : _GEN4300;
wire  _GEN4326 = io_x[72] ? _GEN4325 : _GEN4275;
wire  _GEN4327 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4328 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4329 = io_x[17] ? _GEN4328 : _GEN4327;
wire  _GEN4330 = io_x[75] ? _GEN1899 : _GEN4329;
wire  _GEN4331 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4332 = io_x[17] ? _GEN4331 : _GEN1731;
wire  _GEN4333 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4334 = io_x[17] ? _GEN4333 : _GEN1731;
wire  _GEN4335 = io_x[75] ? _GEN4334 : _GEN4332;
wire  _GEN4336 = io_x[25] ? _GEN4335 : _GEN4330;
wire  _GEN4337 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4338 = io_x[17] ? _GEN4337 : _GEN1711;
wire  _GEN4339 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN4340 = io_x[75] ? _GEN4339 : _GEN4338;
wire  _GEN4341 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4342 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4343 = io_x[17] ? _GEN4342 : _GEN4341;
wire  _GEN4344 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4345 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4346 = io_x[17] ? _GEN4345 : _GEN4344;
wire  _GEN4347 = io_x[75] ? _GEN4346 : _GEN4343;
wire  _GEN4348 = io_x[25] ? _GEN4347 : _GEN4340;
wire  _GEN4349 = io_x[37] ? _GEN4348 : _GEN4336;
wire  _GEN4350 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4351 = io_x[17] ? _GEN4350 : _GEN1731;
wire  _GEN4352 = io_x[75] ? _GEN4351 : _GEN1899;
wire  _GEN4353 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4354 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4355 = io_x[17] ? _GEN4354 : _GEN4353;
wire  _GEN4356 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4357 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4358 = io_x[17] ? _GEN4357 : _GEN4356;
wire  _GEN4359 = io_x[75] ? _GEN4358 : _GEN4355;
wire  _GEN4360 = io_x[25] ? _GEN4359 : _GEN4352;
wire  _GEN4361 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4362 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4363 = io_x[17] ? _GEN4362 : _GEN4361;
wire  _GEN4364 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4365 = io_x[17] ? _GEN4364 : _GEN1731;
wire  _GEN4366 = io_x[75] ? _GEN4365 : _GEN4363;
wire  _GEN4367 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4368 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4369 = io_x[17] ? _GEN4368 : _GEN4367;
wire  _GEN4370 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4371 = io_x[17] ? _GEN4370 : _GEN1711;
wire  _GEN4372 = io_x[75] ? _GEN4371 : _GEN4369;
wire  _GEN4373 = io_x[25] ? _GEN4372 : _GEN4366;
wire  _GEN4374 = io_x[37] ? _GEN4373 : _GEN4360;
wire  _GEN4375 = io_x[39] ? _GEN4374 : _GEN4349;
wire  _GEN4376 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4377 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4378 = io_x[17] ? _GEN4377 : _GEN4376;
wire  _GEN4379 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4380 = io_x[17] ? _GEN4379 : _GEN1731;
wire  _GEN4381 = io_x[75] ? _GEN4380 : _GEN4378;
wire  _GEN4382 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4383 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4384 = io_x[17] ? _GEN4383 : _GEN4382;
wire  _GEN4385 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4386 = io_x[17] ? _GEN4385 : _GEN1711;
wire  _GEN4387 = io_x[75] ? _GEN4386 : _GEN4384;
wire  _GEN4388 = io_x[25] ? _GEN4387 : _GEN4381;
wire  _GEN4389 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4390 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4391 = io_x[17] ? _GEN4390 : _GEN4389;
wire  _GEN4392 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4393 = io_x[17] ? _GEN4392 : _GEN1731;
wire  _GEN4394 = io_x[75] ? _GEN4393 : _GEN4391;
wire  _GEN4395 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4396 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4397 = io_x[17] ? _GEN4396 : _GEN4395;
wire  _GEN4398 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4399 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4400 = io_x[17] ? _GEN4399 : _GEN4398;
wire  _GEN4401 = io_x[75] ? _GEN4400 : _GEN4397;
wire  _GEN4402 = io_x[25] ? _GEN4401 : _GEN4394;
wire  _GEN4403 = io_x[37] ? _GEN4402 : _GEN4388;
wire  _GEN4404 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4405 = io_x[17] ? _GEN4404 : _GEN1711;
wire  _GEN4406 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN4407 = io_x[75] ? _GEN4406 : _GEN4405;
wire  _GEN4408 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4409 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4410 = io_x[17] ? _GEN4409 : _GEN4408;
wire  _GEN4411 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4412 = io_x[17] ? _GEN4411 : _GEN1731;
wire  _GEN4413 = io_x[75] ? _GEN4412 : _GEN4410;
wire  _GEN4414 = io_x[25] ? _GEN4413 : _GEN4407;
wire  _GEN4415 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4416 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4417 = io_x[17] ? _GEN4416 : _GEN4415;
wire  _GEN4418 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4419 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4420 = io_x[17] ? _GEN4419 : _GEN4418;
wire  _GEN4421 = io_x[75] ? _GEN4420 : _GEN4417;
wire  _GEN4422 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4423 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4424 = io_x[17] ? _GEN4423 : _GEN4422;
wire  _GEN4425 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4426 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4427 = io_x[17] ? _GEN4426 : _GEN4425;
wire  _GEN4428 = io_x[75] ? _GEN4427 : _GEN4424;
wire  _GEN4429 = io_x[25] ? _GEN4428 : _GEN4421;
wire  _GEN4430 = io_x[37] ? _GEN4429 : _GEN4414;
wire  _GEN4431 = io_x[39] ? _GEN4430 : _GEN4403;
wire  _GEN4432 = io_x[72] ? _GEN4431 : _GEN4375;
wire  _GEN4433 = io_x[29] ? _GEN4432 : _GEN4326;
wire  _GEN4434 = io_x[18] ? _GEN4433 : _GEN4229;
wire  _GEN4435 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4436 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4437 = io_x[17] ? _GEN4436 : _GEN4435;
wire  _GEN4438 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN4439 = io_x[75] ? _GEN4438 : _GEN4437;
wire  _GEN4440 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4441 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4442 = io_x[17] ? _GEN4441 : _GEN4440;
wire  _GEN4443 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4444 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4445 = io_x[17] ? _GEN4444 : _GEN4443;
wire  _GEN4446 = io_x[75] ? _GEN4445 : _GEN4442;
wire  _GEN4447 = io_x[25] ? _GEN4446 : _GEN4439;
wire  _GEN4448 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN4449 = io_x[75] ? _GEN1899 : _GEN4448;
wire  _GEN4450 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4451 = io_x[17] ? _GEN4450 : _GEN1731;
wire  _GEN4452 = io_x[75] ? _GEN4451 : _GEN1899;
wire  _GEN4453 = io_x[25] ? _GEN4452 : _GEN4449;
wire  _GEN4454 = io_x[37] ? _GEN4453 : _GEN4447;
wire  _GEN4455 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4456 = io_x[17] ? _GEN4455 : _GEN1731;
wire  _GEN4457 = io_x[75] ? _GEN1903 : _GEN4456;
wire  _GEN4458 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4459 = io_x[17] ? _GEN1731 : _GEN4458;
wire  _GEN4460 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4461 = io_x[17] ? _GEN1711 : _GEN4460;
wire  _GEN4462 = io_x[75] ? _GEN4461 : _GEN4459;
wire  _GEN4463 = io_x[25] ? _GEN4462 : _GEN4457;
wire  _GEN4464 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4465 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4466 = io_x[17] ? _GEN4465 : _GEN4464;
wire  _GEN4467 = io_x[75] ? _GEN1899 : _GEN4466;
wire  _GEN4468 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4469 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4470 = io_x[17] ? _GEN4469 : _GEN4468;
wire  _GEN4471 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4472 = io_x[17] ? _GEN4471 : _GEN1731;
wire  _GEN4473 = io_x[75] ? _GEN4472 : _GEN4470;
wire  _GEN4474 = io_x[25] ? _GEN4473 : _GEN4467;
wire  _GEN4475 = io_x[37] ? _GEN4474 : _GEN4463;
wire  _GEN4476 = io_x[39] ? _GEN4475 : _GEN4454;
wire  _GEN4477 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4478 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4479 = io_x[17] ? _GEN4478 : _GEN4477;
wire  _GEN4480 = io_x[75] ? _GEN1903 : _GEN4479;
wire  _GEN4481 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4482 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4483 = io_x[17] ? _GEN4482 : _GEN4481;
wire  _GEN4484 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4485 = io_x[17] ? _GEN1711 : _GEN4484;
wire  _GEN4486 = io_x[75] ? _GEN4485 : _GEN4483;
wire  _GEN4487 = io_x[25] ? _GEN4486 : _GEN4480;
wire  _GEN4488 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4489 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4490 = io_x[17] ? _GEN4489 : _GEN4488;
wire  _GEN4491 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4492 = io_x[17] ? _GEN1731 : _GEN4491;
wire  _GEN4493 = io_x[75] ? _GEN4492 : _GEN4490;
wire  _GEN4494 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4495 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4496 = io_x[17] ? _GEN4495 : _GEN4494;
wire  _GEN4497 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4498 = io_x[17] ? _GEN4497 : _GEN1731;
wire  _GEN4499 = io_x[75] ? _GEN4498 : _GEN4496;
wire  _GEN4500 = io_x[25] ? _GEN4499 : _GEN4493;
wire  _GEN4501 = io_x[37] ? _GEN4500 : _GEN4487;
wire  _GEN4502 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4503 = io_x[17] ? _GEN4502 : _GEN1731;
wire  _GEN4504 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4505 = io_x[17] ? _GEN1731 : _GEN4504;
wire  _GEN4506 = io_x[75] ? _GEN4505 : _GEN4503;
wire  _GEN4507 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4508 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4509 = io_x[17] ? _GEN4508 : _GEN4507;
wire  _GEN4510 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN4511 = io_x[75] ? _GEN4510 : _GEN4509;
wire  _GEN4512 = io_x[25] ? _GEN4511 : _GEN4506;
wire  _GEN4513 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4514 = io_x[17] ? _GEN1731 : _GEN4513;
wire  _GEN4515 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4516 = io_x[17] ? _GEN4515 : _GEN1711;
wire  _GEN4517 = io_x[75] ? _GEN4516 : _GEN4514;
wire  _GEN4518 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4519 = io_x[17] ? _GEN4518 : _GEN1731;
wire  _GEN4520 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4521 = io_x[17] ? _GEN1731 : _GEN4520;
wire  _GEN4522 = io_x[75] ? _GEN4521 : _GEN4519;
wire  _GEN4523 = io_x[25] ? _GEN4522 : _GEN4517;
wire  _GEN4524 = io_x[37] ? _GEN4523 : _GEN4512;
wire  _GEN4525 = io_x[39] ? _GEN4524 : _GEN4501;
wire  _GEN4526 = io_x[72] ? _GEN4525 : _GEN4476;
wire  _GEN4527 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4528 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4529 = io_x[17] ? _GEN4528 : _GEN4527;
wire  _GEN4530 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4531 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4532 = io_x[17] ? _GEN4531 : _GEN4530;
wire  _GEN4533 = io_x[75] ? _GEN4532 : _GEN4529;
wire  _GEN4534 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4535 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4536 = io_x[17] ? _GEN4535 : _GEN4534;
wire  _GEN4537 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4538 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4539 = io_x[17] ? _GEN4538 : _GEN4537;
wire  _GEN4540 = io_x[75] ? _GEN4539 : _GEN4536;
wire  _GEN4541 = io_x[25] ? _GEN4540 : _GEN4533;
wire  _GEN4542 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4543 = io_x[17] ? _GEN4542 : _GEN1711;
wire  _GEN4544 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4545 = io_x[17] ? _GEN4544 : _GEN1731;
wire  _GEN4546 = io_x[75] ? _GEN4545 : _GEN4543;
wire  _GEN4547 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4548 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4549 = io_x[17] ? _GEN4548 : _GEN4547;
wire  _GEN4550 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4551 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4552 = io_x[17] ? _GEN4551 : _GEN4550;
wire  _GEN4553 = io_x[75] ? _GEN4552 : _GEN4549;
wire  _GEN4554 = io_x[25] ? _GEN4553 : _GEN4546;
wire  _GEN4555 = io_x[37] ? _GEN4554 : _GEN4541;
wire  _GEN4556 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4557 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4558 = io_x[17] ? _GEN4557 : _GEN4556;
wire  _GEN4559 = io_x[75] ? _GEN1903 : _GEN4558;
wire  _GEN4560 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4561 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4562 = io_x[17] ? _GEN4561 : _GEN4560;
wire  _GEN4563 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4564 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4565 = io_x[17] ? _GEN4564 : _GEN4563;
wire  _GEN4566 = io_x[75] ? _GEN4565 : _GEN4562;
wire  _GEN4567 = io_x[25] ? _GEN4566 : _GEN4559;
wire  _GEN4568 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4569 = io_x[17] ? _GEN1731 : _GEN4568;
wire  _GEN4570 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4571 = io_x[17] ? _GEN4570 : _GEN1731;
wire  _GEN4572 = io_x[75] ? _GEN4571 : _GEN4569;
wire  _GEN4573 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4574 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4575 = io_x[17] ? _GEN4574 : _GEN4573;
wire  _GEN4576 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4577 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4578 = io_x[17] ? _GEN4577 : _GEN4576;
wire  _GEN4579 = io_x[75] ? _GEN4578 : _GEN4575;
wire  _GEN4580 = io_x[25] ? _GEN4579 : _GEN4572;
wire  _GEN4581 = io_x[37] ? _GEN4580 : _GEN4567;
wire  _GEN4582 = io_x[39] ? _GEN4581 : _GEN4555;
wire  _GEN4583 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4584 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4585 = io_x[17] ? _GEN4584 : _GEN4583;
wire  _GEN4586 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4587 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4588 = io_x[17] ? _GEN4587 : _GEN4586;
wire  _GEN4589 = io_x[75] ? _GEN4588 : _GEN4585;
wire  _GEN4590 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4591 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4592 = io_x[17] ? _GEN4591 : _GEN4590;
wire  _GEN4593 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4594 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4595 = io_x[17] ? _GEN4594 : _GEN4593;
wire  _GEN4596 = io_x[75] ? _GEN4595 : _GEN4592;
wire  _GEN4597 = io_x[25] ? _GEN4596 : _GEN4589;
wire  _GEN4598 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4599 = io_x[17] ? _GEN4598 : _GEN1731;
wire  _GEN4600 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4601 = io_x[17] ? _GEN4600 : _GEN1731;
wire  _GEN4602 = io_x[75] ? _GEN4601 : _GEN4599;
wire  _GEN4603 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4604 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4605 = io_x[17] ? _GEN4604 : _GEN4603;
wire  _GEN4606 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4607 = io_x[17] ? _GEN4606 : _GEN1711;
wire  _GEN4608 = io_x[75] ? _GEN4607 : _GEN4605;
wire  _GEN4609 = io_x[25] ? _GEN4608 : _GEN4602;
wire  _GEN4610 = io_x[37] ? _GEN4609 : _GEN4597;
wire  _GEN4611 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4612 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4613 = io_x[17] ? _GEN4612 : _GEN4611;
wire  _GEN4614 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN4615 = io_x[75] ? _GEN4614 : _GEN4613;
wire  _GEN4616 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4617 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4618 = io_x[17] ? _GEN4617 : _GEN4616;
wire  _GEN4619 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4620 = io_x[17] ? _GEN1731 : _GEN4619;
wire  _GEN4621 = io_x[75] ? _GEN4620 : _GEN4618;
wire  _GEN4622 = io_x[25] ? _GEN4621 : _GEN4615;
wire  _GEN4623 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN4624 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN4625 = io_x[75] ? _GEN4624 : _GEN4623;
wire  _GEN4626 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4627 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4628 = io_x[17] ? _GEN4627 : _GEN4626;
wire  _GEN4629 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN4630 = io_x[75] ? _GEN4629 : _GEN4628;
wire  _GEN4631 = io_x[25] ? _GEN4630 : _GEN4625;
wire  _GEN4632 = io_x[37] ? _GEN4631 : _GEN4622;
wire  _GEN4633 = io_x[39] ? _GEN4632 : _GEN4610;
wire  _GEN4634 = io_x[72] ? _GEN4633 : _GEN4582;
wire  _GEN4635 = io_x[29] ? _GEN4634 : _GEN4526;
wire  _GEN4636 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4637 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4638 = io_x[17] ? _GEN4637 : _GEN4636;
wire  _GEN4639 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4640 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4641 = io_x[17] ? _GEN4640 : _GEN4639;
wire  _GEN4642 = io_x[75] ? _GEN4641 : _GEN4638;
wire  _GEN4643 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4644 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4645 = io_x[17] ? _GEN4644 : _GEN4643;
wire  _GEN4646 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4647 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4648 = io_x[17] ? _GEN4647 : _GEN4646;
wire  _GEN4649 = io_x[75] ? _GEN4648 : _GEN4645;
wire  _GEN4650 = io_x[25] ? _GEN4649 : _GEN4642;
wire  _GEN4651 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4652 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4653 = io_x[17] ? _GEN4652 : _GEN4651;
wire  _GEN4654 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4655 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4656 = io_x[17] ? _GEN4655 : _GEN4654;
wire  _GEN4657 = io_x[75] ? _GEN4656 : _GEN4653;
wire  _GEN4658 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4659 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4660 = io_x[17] ? _GEN4659 : _GEN4658;
wire  _GEN4661 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4662 = io_x[17] ? _GEN4661 : _GEN1731;
wire  _GEN4663 = io_x[75] ? _GEN4662 : _GEN4660;
wire  _GEN4664 = io_x[25] ? _GEN4663 : _GEN4657;
wire  _GEN4665 = io_x[37] ? _GEN4664 : _GEN4650;
wire  _GEN4666 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4667 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4668 = io_x[17] ? _GEN4667 : _GEN4666;
wire  _GEN4669 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4670 = io_x[17] ? _GEN4669 : _GEN1731;
wire  _GEN4671 = io_x[75] ? _GEN4670 : _GEN4668;
wire  _GEN4672 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4673 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4674 = io_x[17] ? _GEN4673 : _GEN4672;
wire  _GEN4675 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4676 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4677 = io_x[17] ? _GEN4676 : _GEN4675;
wire  _GEN4678 = io_x[75] ? _GEN4677 : _GEN4674;
wire  _GEN4679 = io_x[25] ? _GEN4678 : _GEN4671;
wire  _GEN4680 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4681 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4682 = io_x[17] ? _GEN4681 : _GEN4680;
wire  _GEN4683 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4684 = io_x[17] ? _GEN4683 : _GEN1731;
wire  _GEN4685 = io_x[75] ? _GEN4684 : _GEN4682;
wire  _GEN4686 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4687 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4688 = io_x[17] ? _GEN4687 : _GEN4686;
wire  _GEN4689 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4690 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4691 = io_x[17] ? _GEN4690 : _GEN4689;
wire  _GEN4692 = io_x[75] ? _GEN4691 : _GEN4688;
wire  _GEN4693 = io_x[25] ? _GEN4692 : _GEN4685;
wire  _GEN4694 = io_x[37] ? _GEN4693 : _GEN4679;
wire  _GEN4695 = io_x[39] ? _GEN4694 : _GEN4665;
wire  _GEN4696 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4697 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4698 = io_x[17] ? _GEN4697 : _GEN4696;
wire  _GEN4699 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4700 = io_x[17] ? _GEN4699 : _GEN1731;
wire  _GEN4701 = io_x[75] ? _GEN4700 : _GEN4698;
wire  _GEN4702 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4703 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4704 = io_x[17] ? _GEN4703 : _GEN4702;
wire  _GEN4705 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4706 = io_x[17] ? _GEN4705 : _GEN1731;
wire  _GEN4707 = io_x[75] ? _GEN4706 : _GEN4704;
wire  _GEN4708 = io_x[25] ? _GEN4707 : _GEN4701;
wire  _GEN4709 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4710 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4711 = io_x[17] ? _GEN4710 : _GEN4709;
wire  _GEN4712 = io_x[75] ? _GEN1899 : _GEN4711;
wire  _GEN4713 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4714 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4715 = io_x[17] ? _GEN4714 : _GEN4713;
wire  _GEN4716 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4717 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4718 = io_x[17] ? _GEN4717 : _GEN4716;
wire  _GEN4719 = io_x[75] ? _GEN4718 : _GEN4715;
wire  _GEN4720 = io_x[25] ? _GEN4719 : _GEN4712;
wire  _GEN4721 = io_x[37] ? _GEN4720 : _GEN4708;
wire  _GEN4722 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4723 = io_x[17] ? _GEN4722 : _GEN1731;
wire  _GEN4724 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4725 = io_x[17] ? _GEN4724 : _GEN1731;
wire  _GEN4726 = io_x[75] ? _GEN4725 : _GEN4723;
wire  _GEN4727 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4728 = io_x[17] ? _GEN4727 : _GEN1711;
wire  _GEN4729 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4730 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4731 = io_x[17] ? _GEN4730 : _GEN4729;
wire  _GEN4732 = io_x[75] ? _GEN4731 : _GEN4728;
wire  _GEN4733 = io_x[25] ? _GEN4732 : _GEN4726;
wire  _GEN4734 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4735 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4736 = io_x[17] ? _GEN4735 : _GEN4734;
wire  _GEN4737 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4738 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4739 = io_x[17] ? _GEN4738 : _GEN4737;
wire  _GEN4740 = io_x[75] ? _GEN4739 : _GEN4736;
wire  _GEN4741 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4742 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4743 = io_x[17] ? _GEN4742 : _GEN4741;
wire  _GEN4744 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4745 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4746 = io_x[17] ? _GEN4745 : _GEN4744;
wire  _GEN4747 = io_x[75] ? _GEN4746 : _GEN4743;
wire  _GEN4748 = io_x[25] ? _GEN4747 : _GEN4740;
wire  _GEN4749 = io_x[37] ? _GEN4748 : _GEN4733;
wire  _GEN4750 = io_x[39] ? _GEN4749 : _GEN4721;
wire  _GEN4751 = io_x[72] ? _GEN4750 : _GEN4695;
wire  _GEN4752 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4753 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4754 = io_x[17] ? _GEN4753 : _GEN4752;
wire  _GEN4755 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4756 = io_x[17] ? _GEN4755 : _GEN1731;
wire  _GEN4757 = io_x[75] ? _GEN4756 : _GEN4754;
wire  _GEN4758 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4759 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4760 = io_x[17] ? _GEN4759 : _GEN4758;
wire  _GEN4761 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4762 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4763 = io_x[17] ? _GEN4762 : _GEN4761;
wire  _GEN4764 = io_x[75] ? _GEN4763 : _GEN4760;
wire  _GEN4765 = io_x[25] ? _GEN4764 : _GEN4757;
wire  _GEN4766 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4767 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4768 = io_x[17] ? _GEN4767 : _GEN4766;
wire  _GEN4769 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4770 = io_x[17] ? _GEN4769 : _GEN1731;
wire  _GEN4771 = io_x[75] ? _GEN4770 : _GEN4768;
wire  _GEN4772 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4773 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4774 = io_x[17] ? _GEN4773 : _GEN4772;
wire  _GEN4775 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4776 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4777 = io_x[17] ? _GEN4776 : _GEN4775;
wire  _GEN4778 = io_x[75] ? _GEN4777 : _GEN4774;
wire  _GEN4779 = io_x[25] ? _GEN4778 : _GEN4771;
wire  _GEN4780 = io_x[37] ? _GEN4779 : _GEN4765;
wire  _GEN4781 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4782 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4783 = io_x[17] ? _GEN4782 : _GEN4781;
wire  _GEN4784 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4785 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4786 = io_x[17] ? _GEN4785 : _GEN4784;
wire  _GEN4787 = io_x[75] ? _GEN4786 : _GEN4783;
wire  _GEN4788 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4789 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4790 = io_x[17] ? _GEN4789 : _GEN4788;
wire  _GEN4791 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4792 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4793 = io_x[17] ? _GEN4792 : _GEN4791;
wire  _GEN4794 = io_x[75] ? _GEN4793 : _GEN4790;
wire  _GEN4795 = io_x[25] ? _GEN4794 : _GEN4787;
wire  _GEN4796 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4797 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4798 = io_x[17] ? _GEN4797 : _GEN4796;
wire  _GEN4799 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4800 = io_x[17] ? _GEN4799 : _GEN1731;
wire  _GEN4801 = io_x[75] ? _GEN4800 : _GEN4798;
wire  _GEN4802 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4803 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4804 = io_x[17] ? _GEN4803 : _GEN4802;
wire  _GEN4805 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4806 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4807 = io_x[17] ? _GEN4806 : _GEN4805;
wire  _GEN4808 = io_x[75] ? _GEN4807 : _GEN4804;
wire  _GEN4809 = io_x[25] ? _GEN4808 : _GEN4801;
wire  _GEN4810 = io_x[37] ? _GEN4809 : _GEN4795;
wire  _GEN4811 = io_x[39] ? _GEN4810 : _GEN4780;
wire  _GEN4812 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4813 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4814 = io_x[17] ? _GEN4813 : _GEN4812;
wire  _GEN4815 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4816 = io_x[17] ? _GEN4815 : _GEN1731;
wire  _GEN4817 = io_x[75] ? _GEN4816 : _GEN4814;
wire  _GEN4818 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4819 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4820 = io_x[17] ? _GEN4819 : _GEN4818;
wire  _GEN4821 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4822 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4823 = io_x[17] ? _GEN4822 : _GEN4821;
wire  _GEN4824 = io_x[75] ? _GEN4823 : _GEN4820;
wire  _GEN4825 = io_x[25] ? _GEN4824 : _GEN4817;
wire  _GEN4826 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4827 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4828 = io_x[17] ? _GEN4827 : _GEN4826;
wire  _GEN4829 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4830 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4831 = io_x[17] ? _GEN4830 : _GEN4829;
wire  _GEN4832 = io_x[75] ? _GEN4831 : _GEN4828;
wire  _GEN4833 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4834 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4835 = io_x[17] ? _GEN4834 : _GEN4833;
wire  _GEN4836 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4837 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4838 = io_x[17] ? _GEN4837 : _GEN4836;
wire  _GEN4839 = io_x[75] ? _GEN4838 : _GEN4835;
wire  _GEN4840 = io_x[25] ? _GEN4839 : _GEN4832;
wire  _GEN4841 = io_x[37] ? _GEN4840 : _GEN4825;
wire  _GEN4842 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4843 = io_x[17] ? _GEN4842 : _GEN1711;
wire  _GEN4844 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4845 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4846 = io_x[17] ? _GEN4845 : _GEN4844;
wire  _GEN4847 = io_x[75] ? _GEN4846 : _GEN4843;
wire  _GEN4848 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4849 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4850 = io_x[17] ? _GEN4849 : _GEN4848;
wire  _GEN4851 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4852 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4853 = io_x[17] ? _GEN4852 : _GEN4851;
wire  _GEN4854 = io_x[75] ? _GEN4853 : _GEN4850;
wire  _GEN4855 = io_x[25] ? _GEN4854 : _GEN4847;
wire  _GEN4856 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4857 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4858 = io_x[17] ? _GEN4857 : _GEN4856;
wire  _GEN4859 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4860 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4861 = io_x[17] ? _GEN4860 : _GEN4859;
wire  _GEN4862 = io_x[75] ? _GEN4861 : _GEN4858;
wire  _GEN4863 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4864 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4865 = io_x[17] ? _GEN4864 : _GEN4863;
wire  _GEN4866 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4867 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4868 = io_x[17] ? _GEN4867 : _GEN4866;
wire  _GEN4869 = io_x[75] ? _GEN4868 : _GEN4865;
wire  _GEN4870 = io_x[25] ? _GEN4869 : _GEN4862;
wire  _GEN4871 = io_x[37] ? _GEN4870 : _GEN4855;
wire  _GEN4872 = io_x[39] ? _GEN4871 : _GEN4841;
wire  _GEN4873 = io_x[72] ? _GEN4872 : _GEN4811;
wire  _GEN4874 = io_x[29] ? _GEN4873 : _GEN4751;
wire  _GEN4875 = io_x[18] ? _GEN4874 : _GEN4635;
wire  _GEN4876 = io_x[19] ? _GEN4875 : _GEN4434;
wire  _GEN4877 = io_x[24] ? _GEN4876 : _GEN4021;
wire  _GEN4878 = io_x[23] ? _GEN4877 : _GEN3260;
wire  _GEN4879 = 1'b1;
wire  _GEN4880 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN4881 = io_x[25] ? _GEN2288 : _GEN4880;
wire  _GEN4882 = io_x[37] ? _GEN4881 : _GEN4879;
wire  _GEN4883 = 1'b1;
wire  _GEN4884 = io_x[39] ? _GEN4883 : _GEN4882;
wire  _GEN4885 = 1'b0;
wire  _GEN4886 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN4887 = 1'b0;
wire  _GEN4888 = io_x[39] ? _GEN4887 : _GEN4886;
wire  _GEN4889 = io_x[72] ? _GEN4888 : _GEN4884;
wire  _GEN4890 = 1'b0;
wire  _GEN4891 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN4892 = io_x[25] ? _GEN4891 : _GEN2288;
wire  _GEN4893 = io_x[37] ? _GEN4885 : _GEN4892;
wire  _GEN4894 = io_x[39] ? _GEN4883 : _GEN4893;
wire  _GEN4895 = io_x[72] ? _GEN4894 : _GEN4890;
wire  _GEN4896 = io_x[29] ? _GEN4895 : _GEN4889;
wire  _GEN4897 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN4898 = io_x[25] ? _GEN2288 : _GEN4897;
wire  _GEN4899 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4900 = io_x[17] ? _GEN4899 : _GEN1711;
wire  _GEN4901 = io_x[75] ? _GEN1899 : _GEN4900;
wire  _GEN4902 = io_x[25] ? _GEN2288 : _GEN4901;
wire  _GEN4903 = io_x[37] ? _GEN4902 : _GEN4898;
wire  _GEN4904 = io_x[39] ? _GEN4883 : _GEN4903;
wire  _GEN4905 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN4906 = io_x[39] ? _GEN4887 : _GEN4905;
wire  _GEN4907 = io_x[72] ? _GEN4906 : _GEN4904;
wire  _GEN4908 = io_x[39] ? _GEN4883 : _GEN4887;
wire  _GEN4909 = io_x[72] ? _GEN4890 : _GEN4908;
wire  _GEN4910 = io_x[29] ? _GEN4909 : _GEN4907;
wire  _GEN4911 = io_x[18] ? _GEN4910 : _GEN4896;
wire  _GEN4912 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4913 = io_x[17] ? _GEN4912 : _GEN1731;
wire  _GEN4914 = io_x[75] ? _GEN1899 : _GEN4913;
wire  _GEN4915 = io_x[25] ? _GEN2288 : _GEN4914;
wire  _GEN4916 = io_x[37] ? _GEN4915 : _GEN4879;
wire  _GEN4917 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN4918 = io_x[37] ? _GEN4917 : _GEN4879;
wire  _GEN4919 = io_x[39] ? _GEN4918 : _GEN4916;
wire  _GEN4920 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN4921 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN4922 = io_x[37] ? _GEN4921 : _GEN4920;
wire  _GEN4923 = io_x[39] ? _GEN4883 : _GEN4922;
wire  _GEN4924 = io_x[72] ? _GEN4923 : _GEN4919;
wire  _GEN4925 = 1'b0;
wire  _GEN4926 = io_x[29] ? _GEN4925 : _GEN4924;
wire  _GEN4927 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4928 = io_x[17] ? _GEN4927 : _GEN1731;
wire  _GEN4929 = io_x[75] ? _GEN1899 : _GEN4928;
wire  _GEN4930 = io_x[25] ? _GEN2288 : _GEN4929;
wire  _GEN4931 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN4932 = io_x[75] ? _GEN1899 : _GEN4931;
wire  _GEN4933 = io_x[25] ? _GEN2288 : _GEN4932;
wire  _GEN4934 = io_x[37] ? _GEN4933 : _GEN4930;
wire  _GEN4935 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4936 = io_x[17] ? _GEN1731 : _GEN4935;
wire  _GEN4937 = io_x[75] ? _GEN1899 : _GEN4936;
wire  _GEN4938 = io_x[25] ? _GEN2288 : _GEN4937;
wire  _GEN4939 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN4940 = io_x[25] ? _GEN2288 : _GEN4939;
wire  _GEN4941 = io_x[37] ? _GEN4940 : _GEN4938;
wire  _GEN4942 = io_x[39] ? _GEN4941 : _GEN4934;
wire  _GEN4943 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN4944 = io_x[25] ? _GEN4943 : _GEN2239;
wire  _GEN4945 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN4946 = io_x[37] ? _GEN4945 : _GEN4944;
wire  _GEN4947 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN4948 = io_x[39] ? _GEN4947 : _GEN4946;
wire  _GEN4949 = io_x[72] ? _GEN4948 : _GEN4942;
wire  _GEN4950 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN4951 = io_x[25] ? _GEN4950 : _GEN2288;
wire  _GEN4952 = io_x[37] ? _GEN4951 : _GEN4885;
wire  _GEN4953 = io_x[39] ? _GEN4883 : _GEN4952;
wire  _GEN4954 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4955 = io_x[17] ? _GEN4954 : _GEN1731;
wire  _GEN4956 = io_x[75] ? _GEN4955 : _GEN1903;
wire  _GEN4957 = io_x[25] ? _GEN2239 : _GEN4956;
wire  _GEN4958 = io_x[37] ? _GEN4879 : _GEN4957;
wire  _GEN4959 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4960 = io_x[17] ? _GEN4959 : _GEN1731;
wire  _GEN4961 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4962 = io_x[17] ? _GEN4961 : _GEN1731;
wire  _GEN4963 = io_x[75] ? _GEN4962 : _GEN4960;
wire  _GEN4964 = io_x[25] ? _GEN2288 : _GEN4963;
wire  _GEN4965 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN4966 = io_x[25] ? _GEN4965 : _GEN2239;
wire  _GEN4967 = io_x[37] ? _GEN4966 : _GEN4964;
wire  _GEN4968 = io_x[39] ? _GEN4967 : _GEN4958;
wire  _GEN4969 = io_x[72] ? _GEN4968 : _GEN4953;
wire  _GEN4970 = io_x[29] ? _GEN4969 : _GEN4949;
wire  _GEN4971 = io_x[18] ? _GEN4970 : _GEN4926;
wire  _GEN4972 = io_x[19] ? _GEN4971 : _GEN4911;
wire  _GEN4973 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN4974 = io_x[17] ? _GEN4973 : _GEN1731;
wire  _GEN4975 = io_x[75] ? _GEN1903 : _GEN4974;
wire  _GEN4976 = io_x[25] ? _GEN2288 : _GEN4975;
wire  _GEN4977 = io_x[37] ? _GEN4976 : _GEN4885;
wire  _GEN4978 = io_x[39] ? _GEN4883 : _GEN4977;
wire  _GEN4979 = 1'b1;
wire  _GEN4980 = io_x[72] ? _GEN4979 : _GEN4978;
wire  _GEN4981 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN4982 = io_x[37] ? _GEN4981 : _GEN4879;
wire  _GEN4983 = io_x[39] ? _GEN4883 : _GEN4982;
wire  _GEN4984 = io_x[39] ? _GEN4887 : _GEN4883;
wire  _GEN4985 = io_x[72] ? _GEN4984 : _GEN4983;
wire  _GEN4986 = io_x[29] ? _GEN4985 : _GEN4980;
wire  _GEN4987 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN4988 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN4989 = io_x[75] ? _GEN1899 : _GEN4988;
wire  _GEN4990 = io_x[25] ? _GEN2288 : _GEN4989;
wire  _GEN4991 = io_x[37] ? _GEN4990 : _GEN4987;
wire  _GEN4992 = io_x[39] ? _GEN4887 : _GEN4991;
wire  _GEN4993 = io_x[72] ? _GEN4890 : _GEN4992;
wire  _GEN4994 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN4995 = io_x[17] ? _GEN4994 : _GEN1731;
wire  _GEN4996 = io_x[75] ? _GEN1899 : _GEN4995;
wire  _GEN4997 = io_x[25] ? _GEN2239 : _GEN4996;
wire  _GEN4998 = io_x[37] ? _GEN4997 : _GEN4879;
wire  _GEN4999 = io_x[39] ? _GEN4887 : _GEN4998;
wire  _GEN5000 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN5001 = io_x[39] ? _GEN4883 : _GEN5000;
wire  _GEN5002 = io_x[72] ? _GEN5001 : _GEN4999;
wire  _GEN5003 = io_x[29] ? _GEN5002 : _GEN4993;
wire  _GEN5004 = io_x[18] ? _GEN5003 : _GEN4986;
wire  _GEN5005 = 1'b1;
wire  _GEN5006 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5007 = io_x[17] ? _GEN1731 : _GEN5006;
wire  _GEN5008 = io_x[75] ? _GEN5007 : _GEN1903;
wire  _GEN5009 = io_x[25] ? _GEN5008 : _GEN2239;
wire  _GEN5010 = io_x[37] ? _GEN4885 : _GEN5009;
wire  _GEN5011 = io_x[39] ? _GEN4887 : _GEN5010;
wire  _GEN5012 = io_x[72] ? _GEN5011 : _GEN4890;
wire  _GEN5013 = io_x[29] ? _GEN5012 : _GEN5005;
wire  _GEN5014 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5015 = io_x[37] ? _GEN4885 : _GEN5014;
wire  _GEN5016 = io_x[39] ? _GEN4887 : _GEN5015;
wire  _GEN5017 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5018 = io_x[75] ? _GEN5017 : _GEN1899;
wire  _GEN5019 = io_x[25] ? _GEN5018 : _GEN2239;
wire  _GEN5020 = io_x[37] ? _GEN4879 : _GEN5019;
wire  _GEN5021 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN5022 = io_x[39] ? _GEN5021 : _GEN5020;
wire  _GEN5023 = io_x[72] ? _GEN5022 : _GEN5016;
wire  _GEN5024 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5025 = io_x[17] ? _GEN5024 : _GEN1731;
wire  _GEN5026 = io_x[75] ? _GEN1899 : _GEN5025;
wire  _GEN5027 = io_x[25] ? _GEN5026 : _GEN2288;
wire  _GEN5028 = io_x[37] ? _GEN5027 : _GEN4879;
wire  _GEN5029 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5030 = io_x[37] ? _GEN4879 : _GEN5029;
wire  _GEN5031 = io_x[39] ? _GEN5030 : _GEN5028;
wire  _GEN5032 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5033 = io_x[25] ? _GEN2239 : _GEN5032;
wire  _GEN5034 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5035 = io_x[17] ? _GEN5034 : _GEN1731;
wire  _GEN5036 = io_x[75] ? _GEN1899 : _GEN5035;
wire  _GEN5037 = io_x[25] ? _GEN5036 : _GEN2288;
wire  _GEN5038 = io_x[37] ? _GEN5037 : _GEN5033;
wire  _GEN5039 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN5040 = io_x[39] ? _GEN5039 : _GEN5038;
wire  _GEN5041 = io_x[72] ? _GEN5040 : _GEN5031;
wire  _GEN5042 = io_x[29] ? _GEN5041 : _GEN5023;
wire  _GEN5043 = io_x[18] ? _GEN5042 : _GEN5013;
wire  _GEN5044 = io_x[19] ? _GEN5043 : _GEN5004;
wire  _GEN5045 = io_x[24] ? _GEN5044 : _GEN4972;
wire  _GEN5046 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5047 = io_x[25] ? _GEN2288 : _GEN5046;
wire  _GEN5048 = io_x[37] ? _GEN5047 : _GEN4879;
wire  _GEN5049 = io_x[39] ? _GEN5048 : _GEN4887;
wire  _GEN5050 = io_x[72] ? _GEN5049 : _GEN4890;
wire  _GEN5051 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN5052 = io_x[39] ? _GEN4883 : _GEN5051;
wire  _GEN5053 = io_x[72] ? _GEN5052 : _GEN4890;
wire  _GEN5054 = io_x[29] ? _GEN5053 : _GEN5050;
wire  _GEN5055 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5056 = io_x[75] ? _GEN1899 : _GEN5055;
wire  _GEN5057 = io_x[25] ? _GEN5056 : _GEN2288;
wire  _GEN5058 = io_x[37] ? _GEN5057 : _GEN4879;
wire  _GEN5059 = io_x[39] ? _GEN5058 : _GEN4887;
wire  _GEN5060 = io_x[72] ? _GEN4890 : _GEN5059;
wire  _GEN5061 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN5062 = io_x[39] ? _GEN4883 : _GEN5061;
wire  _GEN5063 = io_x[72] ? _GEN5062 : _GEN4979;
wire  _GEN5064 = io_x[29] ? _GEN5063 : _GEN5060;
wire  _GEN5065 = io_x[18] ? _GEN5064 : _GEN5054;
wire  _GEN5066 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN5067 = io_x[37] ? _GEN4879 : _GEN5066;
wire  _GEN5068 = io_x[39] ? _GEN4883 : _GEN5067;
wire  _GEN5069 = io_x[72] ? _GEN5068 : _GEN4979;
wire  _GEN5070 = io_x[29] ? _GEN4925 : _GEN5069;
wire  _GEN5071 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5072 = io_x[25] ? _GEN5071 : _GEN2239;
wire  _GEN5073 = io_x[37] ? _GEN4885 : _GEN5072;
wire  _GEN5074 = io_x[39] ? _GEN4887 : _GEN5073;
wire  _GEN5075 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5076 = io_x[17] ? _GEN5075 : _GEN1731;
wire  _GEN5077 = io_x[75] ? _GEN1899 : _GEN5076;
wire  _GEN5078 = io_x[25] ? _GEN5077 : _GEN2288;
wire  _GEN5079 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5080 = io_x[17] ? _GEN5079 : _GEN1731;
wire  _GEN5081 = io_x[75] ? _GEN1903 : _GEN5080;
wire  _GEN5082 = io_x[25] ? _GEN5081 : _GEN2288;
wire  _GEN5083 = io_x[37] ? _GEN5082 : _GEN5078;
wire  _GEN5084 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN5085 = io_x[39] ? _GEN5084 : _GEN5083;
wire  _GEN5086 = io_x[72] ? _GEN5085 : _GEN5074;
wire  _GEN5087 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5088 = io_x[17] ? _GEN5087 : _GEN1731;
wire  _GEN5089 = io_x[75] ? _GEN5088 : _GEN1899;
wire  _GEN5090 = io_x[25] ? _GEN5089 : _GEN2288;
wire  _GEN5091 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5092 = io_x[25] ? _GEN5091 : _GEN2288;
wire  _GEN5093 = io_x[37] ? _GEN5092 : _GEN5090;
wire  _GEN5094 = io_x[39] ? _GEN4883 : _GEN5093;
wire  _GEN5095 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5096 = io_x[17] ? _GEN5095 : _GEN1731;
wire  _GEN5097 = io_x[75] ? _GEN1899 : _GEN5096;
wire  _GEN5098 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5099 = io_x[25] ? _GEN5098 : _GEN5097;
wire  _GEN5100 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5101 = io_x[17] ? _GEN5100 : _GEN1731;
wire  _GEN5102 = io_x[75] ? _GEN1899 : _GEN5101;
wire  _GEN5103 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5104 = io_x[25] ? _GEN5103 : _GEN5102;
wire  _GEN5105 = io_x[37] ? _GEN5104 : _GEN5099;
wire  _GEN5106 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5107 = io_x[75] ? _GEN1899 : _GEN5106;
wire  _GEN5108 = io_x[25] ? _GEN5107 : _GEN2288;
wire  _GEN5109 = io_x[37] ? _GEN4879 : _GEN5108;
wire  _GEN5110 = io_x[39] ? _GEN5109 : _GEN5105;
wire  _GEN5111 = io_x[72] ? _GEN5110 : _GEN5094;
wire  _GEN5112 = io_x[29] ? _GEN5111 : _GEN5086;
wire  _GEN5113 = io_x[18] ? _GEN5112 : _GEN5070;
wire  _GEN5114 = io_x[19] ? _GEN5113 : _GEN5065;
wire  _GEN5115 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5116 = io_x[75] ? _GEN1899 : _GEN5115;
wire  _GEN5117 = io_x[25] ? _GEN5116 : _GEN2288;
wire  _GEN5118 = io_x[37] ? _GEN4879 : _GEN5117;
wire  _GEN5119 = io_x[39] ? _GEN5118 : _GEN4883;
wire  _GEN5120 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5121 = io_x[25] ? _GEN5120 : _GEN2288;
wire  _GEN5122 = io_x[37] ? _GEN4879 : _GEN5121;
wire  _GEN5123 = io_x[39] ? _GEN4887 : _GEN5122;
wire  _GEN5124 = io_x[72] ? _GEN5123 : _GEN5119;
wire  _GEN5125 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5126 = io_x[25] ? _GEN5125 : _GEN2288;
wire  _GEN5127 = io_x[37] ? _GEN5126 : _GEN4885;
wire  _GEN5128 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5129 = io_x[25] ? _GEN5128 : _GEN2288;
wire  _GEN5130 = io_x[37] ? _GEN5129 : _GEN4879;
wire  _GEN5131 = io_x[39] ? _GEN5130 : _GEN5127;
wire  _GEN5132 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5133 = io_x[25] ? _GEN5132 : _GEN2288;
wire  _GEN5134 = io_x[37] ? _GEN5133 : _GEN4879;
wire  _GEN5135 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN5136 = io_x[39] ? _GEN5135 : _GEN5134;
wire  _GEN5137 = io_x[72] ? _GEN5136 : _GEN5131;
wire  _GEN5138 = io_x[29] ? _GEN5137 : _GEN5124;
wire  _GEN5139 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5140 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5141 = io_x[37] ? _GEN5140 : _GEN5139;
wire  _GEN5142 = io_x[39] ? _GEN4883 : _GEN5141;
wire  _GEN5143 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5144 = io_x[25] ? _GEN5143 : _GEN2288;
wire  _GEN5145 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5146 = io_x[37] ? _GEN5145 : _GEN5144;
wire  _GEN5147 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5148 = io_x[17] ? _GEN5147 : _GEN1731;
wire  _GEN5149 = io_x[75] ? _GEN5148 : _GEN1899;
wire  _GEN5150 = io_x[25] ? _GEN5149 : _GEN2288;
wire  _GEN5151 = io_x[37] ? _GEN5150 : _GEN4885;
wire  _GEN5152 = io_x[39] ? _GEN5151 : _GEN5146;
wire  _GEN5153 = io_x[72] ? _GEN5152 : _GEN5142;
wire  _GEN5154 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5155 = io_x[17] ? _GEN5154 : _GEN1731;
wire  _GEN5156 = io_x[75] ? _GEN1899 : _GEN5155;
wire  _GEN5157 = io_x[25] ? _GEN5156 : _GEN2239;
wire  _GEN5158 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5159 = io_x[75] ? _GEN1899 : _GEN5158;
wire  _GEN5160 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5161 = io_x[17] ? _GEN5160 : _GEN1731;
wire  _GEN5162 = io_x[75] ? _GEN1899 : _GEN5161;
wire  _GEN5163 = io_x[25] ? _GEN5162 : _GEN5159;
wire  _GEN5164 = io_x[37] ? _GEN5163 : _GEN5157;
wire  _GEN5165 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5166 = io_x[25] ? _GEN5165 : _GEN2288;
wire  _GEN5167 = io_x[37] ? _GEN5166 : _GEN4879;
wire  _GEN5168 = io_x[39] ? _GEN5167 : _GEN5164;
wire  _GEN5169 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5170 = io_x[75] ? _GEN5169 : _GEN1899;
wire  _GEN5171 = io_x[25] ? _GEN5170 : _GEN2288;
wire  _GEN5172 = io_x[37] ? _GEN4885 : _GEN5171;
wire  _GEN5173 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN5174 = io_x[39] ? _GEN5173 : _GEN5172;
wire  _GEN5175 = io_x[72] ? _GEN5174 : _GEN5168;
wire  _GEN5176 = io_x[29] ? _GEN5175 : _GEN5153;
wire  _GEN5177 = io_x[18] ? _GEN5176 : _GEN5138;
wire  _GEN5178 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN5179 = io_x[39] ? _GEN4883 : _GEN5178;
wire  _GEN5180 = io_x[72] ? _GEN4979 : _GEN5179;
wire  _GEN5181 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5182 = io_x[75] ? _GEN5181 : _GEN1899;
wire  _GEN5183 = io_x[25] ? _GEN5182 : _GEN2288;
wire  _GEN5184 = io_x[37] ? _GEN4885 : _GEN5183;
wire  _GEN5185 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5186 = io_x[75] ? _GEN5185 : _GEN1903;
wire  _GEN5187 = io_x[25] ? _GEN5186 : _GEN2288;
wire  _GEN5188 = io_x[37] ? _GEN5187 : _GEN4879;
wire  _GEN5189 = io_x[39] ? _GEN5188 : _GEN5184;
wire  _GEN5190 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5191 = io_x[17] ? _GEN1731 : _GEN5190;
wire  _GEN5192 = io_x[75] ? _GEN5191 : _GEN1903;
wire  _GEN5193 = io_x[25] ? _GEN5192 : _GEN2288;
wire  _GEN5194 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5195 = io_x[25] ? _GEN5194 : _GEN2239;
wire  _GEN5196 = io_x[37] ? _GEN5195 : _GEN5193;
wire  _GEN5197 = io_x[39] ? _GEN4887 : _GEN5196;
wire  _GEN5198 = io_x[72] ? _GEN5197 : _GEN5189;
wire  _GEN5199 = io_x[29] ? _GEN5198 : _GEN5180;
wire  _GEN5200 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5201 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5202 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5203 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5204 = io_x[17] ? _GEN5203 : _GEN5202;
wire  _GEN5205 = io_x[75] ? _GEN1899 : _GEN5204;
wire  _GEN5206 = io_x[25] ? _GEN5205 : _GEN5201;
wire  _GEN5207 = io_x[37] ? _GEN5206 : _GEN5200;
wire  _GEN5208 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5209 = io_x[75] ? _GEN1903 : _GEN5208;
wire  _GEN5210 = io_x[25] ? _GEN5209 : _GEN2239;
wire  _GEN5211 = io_x[37] ? _GEN4879 : _GEN5210;
wire  _GEN5212 = io_x[39] ? _GEN5211 : _GEN5207;
wire  _GEN5213 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5214 = io_x[25] ? _GEN2239 : _GEN5213;
wire  _GEN5215 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5216 = io_x[25] ? _GEN5215 : _GEN2239;
wire  _GEN5217 = io_x[37] ? _GEN5216 : _GEN5214;
wire  _GEN5218 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5219 = io_x[37] ? _GEN4885 : _GEN5218;
wire  _GEN5220 = io_x[39] ? _GEN5219 : _GEN5217;
wire  _GEN5221 = io_x[72] ? _GEN5220 : _GEN5212;
wire  _GEN5222 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5223 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5224 = io_x[17] ? _GEN5223 : _GEN1711;
wire  _GEN5225 = io_x[75] ? _GEN5224 : _GEN1899;
wire  _GEN5226 = io_x[25] ? _GEN5225 : _GEN5222;
wire  _GEN5227 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5228 = io_x[17] ? _GEN1731 : _GEN5227;
wire  _GEN5229 = io_x[75] ? _GEN1899 : _GEN5228;
wire  _GEN5230 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5231 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5232 = io_x[17] ? _GEN5231 : _GEN5230;
wire  _GEN5233 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5234 = io_x[75] ? _GEN5233 : _GEN5232;
wire  _GEN5235 = io_x[25] ? _GEN5234 : _GEN5229;
wire  _GEN5236 = io_x[37] ? _GEN5235 : _GEN5226;
wire  _GEN5237 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5238 = io_x[17] ? _GEN1731 : _GEN5237;
wire  _GEN5239 = io_x[75] ? _GEN5238 : _GEN1899;
wire  _GEN5240 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5241 = io_x[17] ? _GEN1731 : _GEN5240;
wire  _GEN5242 = io_x[75] ? _GEN5241 : _GEN1899;
wire  _GEN5243 = io_x[25] ? _GEN5242 : _GEN5239;
wire  _GEN5244 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5245 = io_x[17] ? _GEN5244 : _GEN1731;
wire  _GEN5246 = io_x[75] ? _GEN1899 : _GEN5245;
wire  _GEN5247 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5248 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5249 = io_x[17] ? _GEN5248 : _GEN1711;
wire  _GEN5250 = io_x[75] ? _GEN5249 : _GEN5247;
wire  _GEN5251 = io_x[25] ? _GEN5250 : _GEN5246;
wire  _GEN5252 = io_x[37] ? _GEN5251 : _GEN5243;
wire  _GEN5253 = io_x[39] ? _GEN5252 : _GEN5236;
wire  _GEN5254 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5255 = io_x[17] ? _GEN5254 : _GEN1731;
wire  _GEN5256 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5257 = io_x[17] ? _GEN5256 : _GEN1731;
wire  _GEN5258 = io_x[75] ? _GEN5257 : _GEN5255;
wire  _GEN5259 = io_x[25] ? _GEN5258 : _GEN2239;
wire  _GEN5260 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5261 = io_x[17] ? _GEN5260 : _GEN1731;
wire  _GEN5262 = io_x[75] ? _GEN5261 : _GEN1903;
wire  _GEN5263 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5264 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5265 = io_x[17] ? _GEN5264 : _GEN5263;
wire  _GEN5266 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5267 = io_x[17] ? _GEN5266 : _GEN1711;
wire  _GEN5268 = io_x[75] ? _GEN5267 : _GEN5265;
wire  _GEN5269 = io_x[25] ? _GEN5268 : _GEN5262;
wire  _GEN5270 = io_x[37] ? _GEN5269 : _GEN5259;
wire  _GEN5271 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5272 = io_x[17] ? _GEN5271 : _GEN1731;
wire  _GEN5273 = io_x[75] ? _GEN5272 : _GEN1899;
wire  _GEN5274 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5275 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5276 = io_x[17] ? _GEN5275 : _GEN5274;
wire  _GEN5277 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5278 = io_x[17] ? _GEN5277 : _GEN1731;
wire  _GEN5279 = io_x[75] ? _GEN5278 : _GEN5276;
wire  _GEN5280 = io_x[25] ? _GEN5279 : _GEN5273;
wire  _GEN5281 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5282 = io_x[17] ? _GEN5281 : _GEN1711;
wire  _GEN5283 = io_x[75] ? _GEN5282 : _GEN1903;
wire  _GEN5284 = io_x[25] ? _GEN5283 : _GEN2239;
wire  _GEN5285 = io_x[37] ? _GEN5284 : _GEN5280;
wire  _GEN5286 = io_x[39] ? _GEN5285 : _GEN5270;
wire  _GEN5287 = io_x[72] ? _GEN5286 : _GEN5253;
wire  _GEN5288 = io_x[29] ? _GEN5287 : _GEN5221;
wire  _GEN5289 = io_x[18] ? _GEN5288 : _GEN5199;
wire  _GEN5290 = io_x[19] ? _GEN5289 : _GEN5177;
wire  _GEN5291 = io_x[24] ? _GEN5290 : _GEN5114;
wire  _GEN5292 = io_x[23] ? _GEN5291 : _GEN5045;
wire  _GEN5293 = io_x[33] ? _GEN5292 : _GEN4878;
wire  _GEN5294 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5295 = io_x[17] ? _GEN5294 : _GEN1711;
wire  _GEN5296 = io_x[75] ? _GEN1899 : _GEN5295;
wire  _GEN5297 = io_x[25] ? _GEN2288 : _GEN5296;
wire  _GEN5298 = io_x[37] ? _GEN5297 : _GEN4879;
wire  _GEN5299 = io_x[39] ? _GEN4883 : _GEN5298;
wire  _GEN5300 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5301 = io_x[17] ? _GEN5300 : _GEN1731;
wire  _GEN5302 = io_x[75] ? _GEN5301 : _GEN1899;
wire  _GEN5303 = io_x[25] ? _GEN5302 : _GEN2288;
wire  _GEN5304 = io_x[37] ? _GEN4879 : _GEN5303;
wire  _GEN5305 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5306 = io_x[25] ? _GEN5305 : _GEN2288;
wire  _GEN5307 = io_x[37] ? _GEN5306 : _GEN4879;
wire  _GEN5308 = io_x[39] ? _GEN5307 : _GEN5304;
wire  _GEN5309 = io_x[72] ? _GEN5308 : _GEN5299;
wire  _GEN5310 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5311 = io_x[17] ? _GEN5310 : _GEN1731;
wire  _GEN5312 = io_x[75] ? _GEN1899 : _GEN5311;
wire  _GEN5313 = io_x[25] ? _GEN2288 : _GEN5312;
wire  _GEN5314 = io_x[37] ? _GEN4879 : _GEN5313;
wire  _GEN5315 = io_x[39] ? _GEN5314 : _GEN4887;
wire  _GEN5316 = io_x[72] ? _GEN4979 : _GEN5315;
wire  _GEN5317 = io_x[29] ? _GEN5316 : _GEN5309;
wire  _GEN5318 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN5319 = io_x[37] ? _GEN5318 : _GEN4879;
wire  _GEN5320 = io_x[39] ? _GEN4883 : _GEN5319;
wire  _GEN5321 = io_x[72] ? _GEN4890 : _GEN5320;
wire  _GEN5322 = io_x[29] ? _GEN4925 : _GEN5321;
wire  _GEN5323 = io_x[18] ? _GEN5322 : _GEN5317;
wire  _GEN5324 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5325 = io_x[25] ? _GEN2288 : _GEN5324;
wire  _GEN5326 = io_x[37] ? _GEN5325 : _GEN4879;
wire  _GEN5327 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5328 = io_x[37] ? _GEN5327 : _GEN4879;
wire  _GEN5329 = io_x[39] ? _GEN5328 : _GEN5326;
wire  _GEN5330 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5331 = io_x[37] ? _GEN4879 : _GEN5330;
wire  _GEN5332 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5333 = io_x[25] ? _GEN2288 : _GEN5332;
wire  _GEN5334 = io_x[37] ? _GEN5333 : _GEN4879;
wire  _GEN5335 = io_x[39] ? _GEN5334 : _GEN5331;
wire  _GEN5336 = io_x[72] ? _GEN5335 : _GEN5329;
wire  _GEN5337 = io_x[29] ? _GEN5005 : _GEN5336;
wire  _GEN5338 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5339 = io_x[75] ? _GEN5338 : _GEN1899;
wire  _GEN5340 = io_x[25] ? _GEN2288 : _GEN5339;
wire  _GEN5341 = io_x[37] ? _GEN5340 : _GEN4879;
wire  _GEN5342 = io_x[39] ? _GEN4883 : _GEN5341;
wire  _GEN5343 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5344 = io_x[75] ? _GEN1899 : _GEN5343;
wire  _GEN5345 = io_x[25] ? _GEN2288 : _GEN5344;
wire  _GEN5346 = io_x[37] ? _GEN5345 : _GEN4879;
wire  _GEN5347 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN5348 = io_x[39] ? _GEN5347 : _GEN5346;
wire  _GEN5349 = io_x[72] ? _GEN5348 : _GEN5342;
wire  _GEN5350 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN5351 = io_x[39] ? _GEN5350 : _GEN4883;
wire  _GEN5352 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5353 = io_x[25] ? _GEN2288 : _GEN5352;
wire  _GEN5354 = io_x[37] ? _GEN5353 : _GEN4879;
wire  _GEN5355 = io_x[39] ? _GEN4883 : _GEN5354;
wire  _GEN5356 = io_x[72] ? _GEN5355 : _GEN5351;
wire  _GEN5357 = io_x[29] ? _GEN5356 : _GEN5349;
wire  _GEN5358 = io_x[18] ? _GEN5357 : _GEN5337;
wire  _GEN5359 = io_x[19] ? _GEN5358 : _GEN5323;
wire  _GEN5360 = 1'b1;
wire  _GEN5361 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5362 = io_x[75] ? _GEN5361 : _GEN1899;
wire  _GEN5363 = io_x[25] ? _GEN2239 : _GEN5362;
wire  _GEN5364 = io_x[37] ? _GEN4879 : _GEN5363;
wire  _GEN5365 = io_x[39] ? _GEN5364 : _GEN4883;
wire  _GEN5366 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5367 = io_x[75] ? _GEN5366 : _GEN1903;
wire  _GEN5368 = io_x[25] ? _GEN2239 : _GEN5367;
wire  _GEN5369 = io_x[37] ? _GEN5368 : _GEN4885;
wire  _GEN5370 = io_x[39] ? _GEN4883 : _GEN5369;
wire  _GEN5371 = io_x[72] ? _GEN5370 : _GEN5365;
wire  _GEN5372 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5373 = io_x[75] ? _GEN1899 : _GEN5372;
wire  _GEN5374 = io_x[25] ? _GEN5373 : _GEN2288;
wire  _GEN5375 = io_x[37] ? _GEN5374 : _GEN4879;
wire  _GEN5376 = io_x[39] ? _GEN4887 : _GEN5375;
wire  _GEN5377 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5378 = io_x[75] ? _GEN1903 : _GEN5377;
wire  _GEN5379 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5380 = io_x[75] ? _GEN1899 : _GEN5379;
wire  _GEN5381 = io_x[25] ? _GEN5380 : _GEN5378;
wire  _GEN5382 = io_x[37] ? _GEN5381 : _GEN4885;
wire  _GEN5383 = io_x[39] ? _GEN4883 : _GEN5382;
wire  _GEN5384 = io_x[72] ? _GEN5383 : _GEN5376;
wire  _GEN5385 = io_x[29] ? _GEN5384 : _GEN5371;
wire  _GEN5386 = io_x[18] ? _GEN5385 : _GEN5360;
wire  _GEN5387 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5388 = io_x[17] ? _GEN1731 : _GEN5387;
wire  _GEN5389 = io_x[75] ? _GEN1899 : _GEN5388;
wire  _GEN5390 = io_x[25] ? _GEN5389 : _GEN2288;
wire  _GEN5391 = io_x[37] ? _GEN4879 : _GEN5390;
wire  _GEN5392 = io_x[39] ? _GEN5391 : _GEN4883;
wire  _GEN5393 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5394 = io_x[37] ? _GEN4879 : _GEN5393;
wire  _GEN5395 = io_x[39] ? _GEN4883 : _GEN5394;
wire  _GEN5396 = io_x[72] ? _GEN5395 : _GEN5392;
wire  _GEN5397 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5398 = io_x[17] ? _GEN1731 : _GEN5397;
wire  _GEN5399 = io_x[75] ? _GEN5398 : _GEN1899;
wire  _GEN5400 = io_x[25] ? _GEN5399 : _GEN2288;
wire  _GEN5401 = io_x[37] ? _GEN5400 : _GEN4885;
wire  _GEN5402 = io_x[39] ? _GEN4883 : _GEN5401;
wire  _GEN5403 = io_x[72] ? _GEN5402 : _GEN4890;
wire  _GEN5404 = io_x[29] ? _GEN5403 : _GEN5396;
wire  _GEN5405 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5406 = io_x[17] ? _GEN5405 : _GEN1731;
wire  _GEN5407 = io_x[75] ? _GEN1899 : _GEN5406;
wire  _GEN5408 = io_x[25] ? _GEN5407 : _GEN2239;
wire  _GEN5409 = io_x[37] ? _GEN5408 : _GEN4879;
wire  _GEN5410 = io_x[39] ? _GEN4887 : _GEN5409;
wire  _GEN5411 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5412 = io_x[17] ? _GEN5411 : _GEN1711;
wire  _GEN5413 = io_x[75] ? _GEN1899 : _GEN5412;
wire  _GEN5414 = io_x[25] ? _GEN2239 : _GEN5413;
wire  _GEN5415 = io_x[37] ? _GEN5414 : _GEN4885;
wire  _GEN5416 = io_x[39] ? _GEN4883 : _GEN5415;
wire  _GEN5417 = io_x[72] ? _GEN5416 : _GEN5410;
wire  _GEN5418 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5419 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5420 = io_x[17] ? _GEN5419 : _GEN5418;
wire  _GEN5421 = io_x[75] ? _GEN1899 : _GEN5420;
wire  _GEN5422 = io_x[25] ? _GEN5421 : _GEN2288;
wire  _GEN5423 = io_x[37] ? _GEN5422 : _GEN4879;
wire  _GEN5424 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5425 = io_x[75] ? _GEN5424 : _GEN1899;
wire  _GEN5426 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5427 = io_x[75] ? _GEN5426 : _GEN1899;
wire  _GEN5428 = io_x[25] ? _GEN5427 : _GEN5425;
wire  _GEN5429 = io_x[37] ? _GEN4885 : _GEN5428;
wire  _GEN5430 = io_x[39] ? _GEN5429 : _GEN5423;
wire  _GEN5431 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5432 = io_x[75] ? _GEN5431 : _GEN1899;
wire  _GEN5433 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5434 = io_x[75] ? _GEN1903 : _GEN5433;
wire  _GEN5435 = io_x[25] ? _GEN5434 : _GEN5432;
wire  _GEN5436 = io_x[37] ? _GEN5435 : _GEN4885;
wire  _GEN5437 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5438 = io_x[17] ? _GEN5437 : _GEN1731;
wire  _GEN5439 = io_x[75] ? _GEN1899 : _GEN5438;
wire  _GEN5440 = io_x[25] ? _GEN5439 : _GEN2239;
wire  _GEN5441 = io_x[37] ? _GEN4879 : _GEN5440;
wire  _GEN5442 = io_x[39] ? _GEN5441 : _GEN5436;
wire  _GEN5443 = io_x[72] ? _GEN5442 : _GEN5430;
wire  _GEN5444 = io_x[29] ? _GEN5443 : _GEN5417;
wire  _GEN5445 = io_x[18] ? _GEN5444 : _GEN5404;
wire  _GEN5446 = io_x[19] ? _GEN5445 : _GEN5386;
wire  _GEN5447 = io_x[24] ? _GEN5446 : _GEN5359;
wire  _GEN5448 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5449 = io_x[17] ? _GEN1731 : _GEN5448;
wire  _GEN5450 = io_x[75] ? _GEN1899 : _GEN5449;
wire  _GEN5451 = io_x[25] ? _GEN5450 : _GEN2288;
wire  _GEN5452 = io_x[37] ? _GEN4885 : _GEN5451;
wire  _GEN5453 = io_x[39] ? _GEN4883 : _GEN5452;
wire  _GEN5454 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN5455 = io_x[39] ? _GEN4883 : _GEN5454;
wire  _GEN5456 = io_x[72] ? _GEN5455 : _GEN5453;
wire  _GEN5457 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5458 = io_x[37] ? _GEN5457 : _GEN4879;
wire  _GEN5459 = io_x[39] ? _GEN5458 : _GEN4883;
wire  _GEN5460 = io_x[72] ? _GEN5459 : _GEN4979;
wire  _GEN5461 = io_x[29] ? _GEN5460 : _GEN5456;
wire  _GEN5462 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5463 = io_x[25] ? _GEN5462 : _GEN2288;
wire  _GEN5464 = io_x[37] ? _GEN5463 : _GEN4879;
wire  _GEN5465 = io_x[39] ? _GEN5464 : _GEN4887;
wire  _GEN5466 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5467 = io_x[25] ? _GEN5466 : _GEN2288;
wire  _GEN5468 = io_x[37] ? _GEN4879 : _GEN5467;
wire  _GEN5469 = io_x[39] ? _GEN5468 : _GEN4887;
wire  _GEN5470 = io_x[72] ? _GEN5469 : _GEN5465;
wire  _GEN5471 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5472 = io_x[75] ? _GEN1903 : _GEN5471;
wire  _GEN5473 = io_x[25] ? _GEN5472 : _GEN2288;
wire  _GEN5474 = io_x[37] ? _GEN5473 : _GEN4879;
wire  _GEN5475 = io_x[39] ? _GEN4883 : _GEN5474;
wire  _GEN5476 = io_x[72] ? _GEN4890 : _GEN5475;
wire  _GEN5477 = io_x[29] ? _GEN5476 : _GEN5470;
wire  _GEN5478 = io_x[18] ? _GEN5477 : _GEN5461;
wire  _GEN5479 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5480 = io_x[75] ? _GEN5479 : _GEN1899;
wire  _GEN5481 = io_x[25] ? _GEN5480 : _GEN2288;
wire  _GEN5482 = io_x[37] ? _GEN4879 : _GEN5481;
wire  _GEN5483 = io_x[39] ? _GEN4883 : _GEN5482;
wire  _GEN5484 = io_x[72] ? _GEN4890 : _GEN5483;
wire  _GEN5485 = io_x[29] ? _GEN5484 : _GEN4925;
wire  _GEN5486 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5487 = io_x[17] ? _GEN5486 : _GEN1731;
wire  _GEN5488 = io_x[75] ? _GEN1899 : _GEN5487;
wire  _GEN5489 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5490 = io_x[17] ? _GEN5489 : _GEN1731;
wire  _GEN5491 = io_x[75] ? _GEN1899 : _GEN5490;
wire  _GEN5492 = io_x[25] ? _GEN5491 : _GEN5488;
wire  _GEN5493 = io_x[37] ? _GEN5492 : _GEN4885;
wire  _GEN5494 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5495 = io_x[25] ? _GEN5494 : _GEN2288;
wire  _GEN5496 = io_x[37] ? _GEN4879 : _GEN5495;
wire  _GEN5497 = io_x[39] ? _GEN5496 : _GEN5493;
wire  _GEN5498 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN5499 = io_x[37] ? _GEN4879 : _GEN5498;
wire  _GEN5500 = io_x[39] ? _GEN5499 : _GEN4887;
wire  _GEN5501 = io_x[72] ? _GEN5500 : _GEN5497;
wire  _GEN5502 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5503 = io_x[17] ? _GEN5502 : _GEN1711;
wire  _GEN5504 = io_x[75] ? _GEN1899 : _GEN5503;
wire  _GEN5505 = io_x[25] ? _GEN5504 : _GEN2288;
wire  _GEN5506 = io_x[37] ? _GEN5505 : _GEN4885;
wire  _GEN5507 = io_x[39] ? _GEN4887 : _GEN5506;
wire  _GEN5508 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5509 = io_x[25] ? _GEN5508 : _GEN2288;
wire  _GEN5510 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5511 = io_x[25] ? _GEN2239 : _GEN5510;
wire  _GEN5512 = io_x[37] ? _GEN5511 : _GEN5509;
wire  _GEN5513 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5514 = io_x[37] ? _GEN5513 : _GEN4885;
wire  _GEN5515 = io_x[39] ? _GEN5514 : _GEN5512;
wire  _GEN5516 = io_x[72] ? _GEN5515 : _GEN5507;
wire  _GEN5517 = io_x[29] ? _GEN5516 : _GEN5501;
wire  _GEN5518 = io_x[18] ? _GEN5517 : _GEN5485;
wire  _GEN5519 = io_x[19] ? _GEN5518 : _GEN5478;
wire  _GEN5520 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN5521 = io_x[39] ? _GEN4883 : _GEN5520;
wire  _GEN5522 = io_x[72] ? _GEN4979 : _GEN5521;
wire  _GEN5523 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5524 = io_x[17] ? _GEN1731 : _GEN5523;
wire  _GEN5525 = io_x[75] ? _GEN1899 : _GEN5524;
wire  _GEN5526 = io_x[25] ? _GEN5525 : _GEN2239;
wire  _GEN5527 = io_x[37] ? _GEN5526 : _GEN4885;
wire  _GEN5528 = io_x[39] ? _GEN4887 : _GEN5527;
wire  _GEN5529 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5530 = io_x[37] ? _GEN4885 : _GEN5529;
wire  _GEN5531 = io_x[39] ? _GEN4883 : _GEN5530;
wire  _GEN5532 = io_x[72] ? _GEN5531 : _GEN5528;
wire  _GEN5533 = io_x[29] ? _GEN5532 : _GEN5522;
wire  _GEN5534 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5535 = io_x[17] ? _GEN5534 : _GEN1711;
wire  _GEN5536 = io_x[75] ? _GEN1899 : _GEN5535;
wire  _GEN5537 = io_x[25] ? _GEN5536 : _GEN2288;
wire  _GEN5538 = io_x[37] ? _GEN5537 : _GEN4879;
wire  _GEN5539 = io_x[39] ? _GEN4883 : _GEN5538;
wire  _GEN5540 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5541 = io_x[17] ? _GEN5540 : _GEN1731;
wire  _GEN5542 = io_x[75] ? _GEN1899 : _GEN5541;
wire  _GEN5543 = io_x[25] ? _GEN5542 : _GEN2288;
wire  _GEN5544 = io_x[37] ? _GEN5543 : _GEN4879;
wire  _GEN5545 = io_x[39] ? _GEN4887 : _GEN5544;
wire  _GEN5546 = io_x[72] ? _GEN5545 : _GEN5539;
wire  _GEN5547 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5548 = io_x[75] ? _GEN1899 : _GEN5547;
wire  _GEN5549 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5550 = io_x[17] ? _GEN5549 : _GEN1731;
wire  _GEN5551 = io_x[75] ? _GEN1899 : _GEN5550;
wire  _GEN5552 = io_x[25] ? _GEN5551 : _GEN5548;
wire  _GEN5553 = io_x[37] ? _GEN5552 : _GEN4879;
wire  _GEN5554 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN5555 = io_x[37] ? _GEN4879 : _GEN5554;
wire  _GEN5556 = io_x[39] ? _GEN5555 : _GEN5553;
wire  _GEN5557 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5558 = io_x[75] ? _GEN1899 : _GEN5557;
wire  _GEN5559 = io_x[25] ? _GEN5558 : _GEN2239;
wire  _GEN5560 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5561 = io_x[17] ? _GEN5560 : _GEN1731;
wire  _GEN5562 = io_x[75] ? _GEN1899 : _GEN5561;
wire  _GEN5563 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5564 = io_x[75] ? _GEN1899 : _GEN5563;
wire  _GEN5565 = io_x[25] ? _GEN5564 : _GEN5562;
wire  _GEN5566 = io_x[37] ? _GEN5565 : _GEN5559;
wire  _GEN5567 = io_x[39] ? _GEN4883 : _GEN5566;
wire  _GEN5568 = io_x[72] ? _GEN5567 : _GEN5556;
wire  _GEN5569 = io_x[29] ? _GEN5568 : _GEN5546;
wire  _GEN5570 = io_x[18] ? _GEN5569 : _GEN5533;
wire  _GEN5571 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5572 = io_x[17] ? _GEN1731 : _GEN5571;
wire  _GEN5573 = io_x[75] ? _GEN5572 : _GEN1903;
wire  _GEN5574 = io_x[25] ? _GEN5573 : _GEN2288;
wire  _GEN5575 = io_x[37] ? _GEN5574 : _GEN4879;
wire  _GEN5576 = io_x[39] ? _GEN4883 : _GEN5575;
wire  _GEN5577 = io_x[72] ? _GEN5576 : _GEN4979;
wire  _GEN5578 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5579 = io_x[25] ? _GEN5578 : _GEN2288;
wire  _GEN5580 = io_x[37] ? _GEN5579 : _GEN4879;
wire  _GEN5581 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5582 = io_x[17] ? _GEN1731 : _GEN5581;
wire  _GEN5583 = io_x[75] ? _GEN5582 : _GEN1899;
wire  _GEN5584 = io_x[25] ? _GEN5583 : _GEN2288;
wire  _GEN5585 = io_x[37] ? _GEN5584 : _GEN4885;
wire  _GEN5586 = io_x[39] ? _GEN5585 : _GEN5580;
wire  _GEN5587 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5588 = io_x[17] ? _GEN1731 : _GEN5587;
wire  _GEN5589 = io_x[75] ? _GEN5588 : _GEN1903;
wire  _GEN5590 = io_x[25] ? _GEN5589 : _GEN2288;
wire  _GEN5591 = io_x[37] ? _GEN5590 : _GEN4885;
wire  _GEN5592 = io_x[39] ? _GEN4883 : _GEN5591;
wire  _GEN5593 = io_x[72] ? _GEN5592 : _GEN5586;
wire  _GEN5594 = io_x[29] ? _GEN5593 : _GEN5577;
wire  _GEN5595 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5596 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5597 = io_x[75] ? _GEN1899 : _GEN5596;
wire  _GEN5598 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5599 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5600 = io_x[17] ? _GEN5599 : _GEN5598;
wire  _GEN5601 = io_x[75] ? _GEN1899 : _GEN5600;
wire  _GEN5602 = io_x[25] ? _GEN5601 : _GEN5597;
wire  _GEN5603 = io_x[37] ? _GEN5602 : _GEN5595;
wire  _GEN5604 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5605 = io_x[75] ? _GEN5604 : _GEN1899;
wire  _GEN5606 = io_x[25] ? _GEN5605 : _GEN2288;
wire  _GEN5607 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN5608 = io_x[37] ? _GEN5607 : _GEN5606;
wire  _GEN5609 = io_x[39] ? _GEN5608 : _GEN5603;
wire  _GEN5610 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5611 = io_x[25] ? _GEN5610 : _GEN2239;
wire  _GEN5612 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5613 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5614 = io_x[17] ? _GEN5613 : _GEN1731;
wire  _GEN5615 = io_x[75] ? _GEN1899 : _GEN5614;
wire  _GEN5616 = io_x[25] ? _GEN5615 : _GEN5612;
wire  _GEN5617 = io_x[37] ? _GEN5616 : _GEN5611;
wire  _GEN5618 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5619 = io_x[37] ? _GEN4885 : _GEN5618;
wire  _GEN5620 = io_x[39] ? _GEN5619 : _GEN5617;
wire  _GEN5621 = io_x[72] ? _GEN5620 : _GEN5609;
wire  _GEN5622 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5623 = io_x[75] ? _GEN1899 : _GEN5622;
wire  _GEN5624 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5625 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5626 = io_x[17] ? _GEN5625 : _GEN5624;
wire  _GEN5627 = io_x[75] ? _GEN1899 : _GEN5626;
wire  _GEN5628 = io_x[25] ? _GEN5627 : _GEN5623;
wire  _GEN5629 = io_x[37] ? _GEN5628 : _GEN4879;
wire  _GEN5630 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5631 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5632 = io_x[75] ? _GEN5631 : _GEN5630;
wire  _GEN5633 = io_x[25] ? _GEN5632 : _GEN2239;
wire  _GEN5634 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5635 = io_x[17] ? _GEN5634 : _GEN1731;
wire  _GEN5636 = io_x[75] ? _GEN1899 : _GEN5635;
wire  _GEN5637 = io_x[25] ? _GEN5636 : _GEN2288;
wire  _GEN5638 = io_x[37] ? _GEN5637 : _GEN5633;
wire  _GEN5639 = io_x[39] ? _GEN5638 : _GEN5629;
wire  _GEN5640 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5641 = io_x[17] ? _GEN5640 : _GEN1731;
wire  _GEN5642 = io_x[75] ? _GEN5641 : _GEN1899;
wire  _GEN5643 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5644 = io_x[17] ? _GEN5643 : _GEN1731;
wire  _GEN5645 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5646 = io_x[17] ? _GEN1731 : _GEN5645;
wire  _GEN5647 = io_x[75] ? _GEN5646 : _GEN5644;
wire  _GEN5648 = io_x[25] ? _GEN5647 : _GEN5642;
wire  _GEN5649 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5650 = io_x[17] ? _GEN5649 : _GEN1731;
wire  _GEN5651 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5652 = io_x[17] ? _GEN1711 : _GEN5651;
wire  _GEN5653 = io_x[75] ? _GEN5652 : _GEN5650;
wire  _GEN5654 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5655 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5656 = io_x[17] ? _GEN5655 : _GEN5654;
wire  _GEN5657 = io_x[75] ? _GEN5656 : _GEN1903;
wire  _GEN5658 = io_x[25] ? _GEN5657 : _GEN5653;
wire  _GEN5659 = io_x[37] ? _GEN5658 : _GEN5648;
wire  _GEN5660 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5661 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5662 = io_x[17] ? _GEN5661 : _GEN5660;
wire  _GEN5663 = io_x[75] ? _GEN1899 : _GEN5662;
wire  _GEN5664 = io_x[25] ? _GEN5663 : _GEN2239;
wire  _GEN5665 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5666 = io_x[75] ? _GEN5665 : _GEN1903;
wire  _GEN5667 = io_x[25] ? _GEN5666 : _GEN2288;
wire  _GEN5668 = io_x[37] ? _GEN5667 : _GEN5664;
wire  _GEN5669 = io_x[39] ? _GEN5668 : _GEN5659;
wire  _GEN5670 = io_x[72] ? _GEN5669 : _GEN5639;
wire  _GEN5671 = io_x[29] ? _GEN5670 : _GEN5621;
wire  _GEN5672 = io_x[18] ? _GEN5671 : _GEN5594;
wire  _GEN5673 = io_x[19] ? _GEN5672 : _GEN5570;
wire  _GEN5674 = io_x[24] ? _GEN5673 : _GEN5519;
wire  _GEN5675 = io_x[23] ? _GEN5674 : _GEN5447;
wire  _GEN5676 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5677 = io_x[75] ? _GEN1903 : _GEN5676;
wire  _GEN5678 = io_x[25] ? _GEN2288 : _GEN5677;
wire  _GEN5679 = io_x[37] ? _GEN5678 : _GEN4885;
wire  _GEN5680 = io_x[39] ? _GEN4883 : _GEN5679;
wire  _GEN5681 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5682 = io_x[17] ? _GEN5681 : _GEN1711;
wire  _GEN5683 = io_x[75] ? _GEN5682 : _GEN1903;
wire  _GEN5684 = io_x[25] ? _GEN2288 : _GEN5683;
wire  _GEN5685 = io_x[37] ? _GEN4879 : _GEN5684;
wire  _GEN5686 = io_x[39] ? _GEN4887 : _GEN5685;
wire  _GEN5687 = io_x[72] ? _GEN5686 : _GEN5680;
wire  _GEN5688 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5689 = io_x[37] ? _GEN5688 : _GEN4879;
wire  _GEN5690 = io_x[39] ? _GEN4887 : _GEN5689;
wire  _GEN5691 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5692 = io_x[17] ? _GEN1731 : _GEN5691;
wire  _GEN5693 = io_x[75] ? _GEN1899 : _GEN5692;
wire  _GEN5694 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5695 = io_x[25] ? _GEN5694 : _GEN5693;
wire  _GEN5696 = io_x[37] ? _GEN4885 : _GEN5695;
wire  _GEN5697 = io_x[39] ? _GEN4887 : _GEN5696;
wire  _GEN5698 = io_x[72] ? _GEN5697 : _GEN5690;
wire  _GEN5699 = io_x[29] ? _GEN5698 : _GEN5687;
wire  _GEN5700 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5701 = io_x[75] ? _GEN1899 : _GEN5700;
wire  _GEN5702 = io_x[25] ? _GEN2288 : _GEN5701;
wire  _GEN5703 = io_x[37] ? _GEN4885 : _GEN5702;
wire  _GEN5704 = io_x[39] ? _GEN4883 : _GEN5703;
wire  _GEN5705 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN5706 = io_x[39] ? _GEN5705 : _GEN4887;
wire  _GEN5707 = io_x[72] ? _GEN5706 : _GEN5704;
wire  _GEN5708 = io_x[72] ? _GEN4979 : _GEN4890;
wire  _GEN5709 = io_x[29] ? _GEN5708 : _GEN5707;
wire  _GEN5710 = io_x[18] ? _GEN5709 : _GEN5699;
wire  _GEN5711 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5712 = io_x[25] ? _GEN2288 : _GEN5711;
wire  _GEN5713 = io_x[37] ? _GEN5712 : _GEN4879;
wire  _GEN5714 = io_x[39] ? _GEN4887 : _GEN5713;
wire  _GEN5715 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5716 = io_x[25] ? _GEN2239 : _GEN5715;
wire  _GEN5717 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN5718 = io_x[37] ? _GEN5717 : _GEN5716;
wire  _GEN5719 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5720 = io_x[75] ? _GEN5719 : _GEN1903;
wire  _GEN5721 = io_x[25] ? _GEN2239 : _GEN5720;
wire  _GEN5722 = io_x[37] ? _GEN5721 : _GEN4879;
wire  _GEN5723 = io_x[39] ? _GEN5722 : _GEN5718;
wire  _GEN5724 = io_x[72] ? _GEN5723 : _GEN5714;
wire  _GEN5725 = io_x[39] ? _GEN4887 : _GEN4883;
wire  _GEN5726 = io_x[72] ? _GEN5725 : _GEN4890;
wire  _GEN5727 = io_x[29] ? _GEN5726 : _GEN5724;
wire  _GEN5728 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5729 = io_x[17] ? _GEN5728 : _GEN1731;
wire  _GEN5730 = io_x[75] ? _GEN1903 : _GEN5729;
wire  _GEN5731 = io_x[25] ? _GEN2288 : _GEN5730;
wire  _GEN5732 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5733 = io_x[75] ? _GEN1899 : _GEN5732;
wire  _GEN5734 = io_x[25] ? _GEN2288 : _GEN5733;
wire  _GEN5735 = io_x[37] ? _GEN5734 : _GEN5731;
wire  _GEN5736 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5737 = io_x[25] ? _GEN2288 : _GEN5736;
wire  _GEN5738 = io_x[37] ? _GEN5737 : _GEN4885;
wire  _GEN5739 = io_x[39] ? _GEN5738 : _GEN5735;
wire  _GEN5740 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5741 = io_x[17] ? _GEN5740 : _GEN1711;
wire  _GEN5742 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5743 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5744 = io_x[17] ? _GEN5743 : _GEN5742;
wire  _GEN5745 = io_x[75] ? _GEN5744 : _GEN5741;
wire  _GEN5746 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5747 = io_x[17] ? _GEN5746 : _GEN1731;
wire  _GEN5748 = io_x[75] ? _GEN5747 : _GEN1899;
wire  _GEN5749 = io_x[25] ? _GEN5748 : _GEN5745;
wire  _GEN5750 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5751 = io_x[17] ? _GEN1711 : _GEN5750;
wire  _GEN5752 = io_x[75] ? _GEN1903 : _GEN5751;
wire  _GEN5753 = io_x[25] ? _GEN2239 : _GEN5752;
wire  _GEN5754 = io_x[37] ? _GEN5753 : _GEN5749;
wire  _GEN5755 = io_x[39] ? _GEN4883 : _GEN5754;
wire  _GEN5756 = io_x[72] ? _GEN5755 : _GEN5739;
wire  _GEN5757 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5758 = io_x[75] ? _GEN1899 : _GEN5757;
wire  _GEN5759 = io_x[25] ? _GEN2288 : _GEN5758;
wire  _GEN5760 = io_x[37] ? _GEN5759 : _GEN4879;
wire  _GEN5761 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5762 = io_x[75] ? _GEN1899 : _GEN5761;
wire  _GEN5763 = io_x[25] ? _GEN2288 : _GEN5762;
wire  _GEN5764 = io_x[37] ? _GEN4885 : _GEN5763;
wire  _GEN5765 = io_x[39] ? _GEN5764 : _GEN5760;
wire  _GEN5766 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5767 = io_x[17] ? _GEN1711 : _GEN5766;
wire  _GEN5768 = io_x[75] ? _GEN5767 : _GEN1899;
wire  _GEN5769 = io_x[25] ? _GEN5768 : _GEN2288;
wire  _GEN5770 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5771 = io_x[75] ? _GEN1903 : _GEN5770;
wire  _GEN5772 = io_x[25] ? _GEN2288 : _GEN5771;
wire  _GEN5773 = io_x[37] ? _GEN5772 : _GEN5769;
wire  _GEN5774 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5775 = io_x[17] ? _GEN5774 : _GEN1731;
wire  _GEN5776 = io_x[75] ? _GEN1899 : _GEN5775;
wire  _GEN5777 = io_x[25] ? _GEN2239 : _GEN5776;
wire  _GEN5778 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN5779 = io_x[37] ? _GEN5778 : _GEN5777;
wire  _GEN5780 = io_x[39] ? _GEN5779 : _GEN5773;
wire  _GEN5781 = io_x[72] ? _GEN5780 : _GEN5765;
wire  _GEN5782 = io_x[29] ? _GEN5781 : _GEN5756;
wire  _GEN5783 = io_x[18] ? _GEN5782 : _GEN5727;
wire  _GEN5784 = io_x[19] ? _GEN5783 : _GEN5710;
wire  _GEN5785 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5786 = io_x[17] ? _GEN5785 : _GEN1731;
wire  _GEN5787 = io_x[75] ? _GEN1899 : _GEN5786;
wire  _GEN5788 = io_x[25] ? _GEN2288 : _GEN5787;
wire  _GEN5789 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5790 = io_x[37] ? _GEN5789 : _GEN5788;
wire  _GEN5791 = io_x[39] ? _GEN4887 : _GEN5790;
wire  _GEN5792 = io_x[72] ? _GEN4890 : _GEN5791;
wire  _GEN5793 = io_x[29] ? _GEN5005 : _GEN5792;
wire  _GEN5794 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5795 = io_x[17] ? _GEN5794 : _GEN1731;
wire  _GEN5796 = io_x[75] ? _GEN1899 : _GEN5795;
wire  _GEN5797 = io_x[25] ? _GEN5796 : _GEN2288;
wire  _GEN5798 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5799 = io_x[75] ? _GEN1899 : _GEN5798;
wire  _GEN5800 = io_x[25] ? _GEN2288 : _GEN5799;
wire  _GEN5801 = io_x[37] ? _GEN5800 : _GEN5797;
wire  _GEN5802 = io_x[39] ? _GEN4883 : _GEN5801;
wire  _GEN5803 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5804 = io_x[17] ? _GEN1731 : _GEN5803;
wire  _GEN5805 = io_x[75] ? _GEN1899 : _GEN5804;
wire  _GEN5806 = io_x[25] ? _GEN2288 : _GEN5805;
wire  _GEN5807 = io_x[37] ? _GEN5806 : _GEN4879;
wire  _GEN5808 = io_x[39] ? _GEN4887 : _GEN5807;
wire  _GEN5809 = io_x[72] ? _GEN5808 : _GEN5802;
wire  _GEN5810 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5811 = io_x[17] ? _GEN5810 : _GEN1731;
wire  _GEN5812 = io_x[75] ? _GEN1899 : _GEN5811;
wire  _GEN5813 = io_x[25] ? _GEN2239 : _GEN5812;
wire  _GEN5814 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5815 = io_x[75] ? _GEN1899 : _GEN5814;
wire  _GEN5816 = io_x[25] ? _GEN5815 : _GEN2239;
wire  _GEN5817 = io_x[37] ? _GEN5816 : _GEN5813;
wire  _GEN5818 = io_x[39] ? _GEN4887 : _GEN5817;
wire  _GEN5819 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN5820 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5821 = io_x[25] ? _GEN5820 : _GEN2288;
wire  _GEN5822 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN5823 = io_x[37] ? _GEN5822 : _GEN5821;
wire  _GEN5824 = io_x[39] ? _GEN5823 : _GEN5819;
wire  _GEN5825 = io_x[72] ? _GEN5824 : _GEN5818;
wire  _GEN5826 = io_x[29] ? _GEN5825 : _GEN5809;
wire  _GEN5827 = io_x[18] ? _GEN5826 : _GEN5793;
wire  _GEN5828 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN5829 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5830 = io_x[17] ? _GEN5829 : _GEN1731;
wire  _GEN5831 = io_x[75] ? _GEN1899 : _GEN5830;
wire  _GEN5832 = io_x[25] ? _GEN5831 : _GEN2288;
wire  _GEN5833 = io_x[37] ? _GEN5832 : _GEN4885;
wire  _GEN5834 = io_x[39] ? _GEN5833 : _GEN5828;
wire  _GEN5835 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5836 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5837 = io_x[75] ? _GEN5836 : _GEN5835;
wire  _GEN5838 = io_x[25] ? _GEN5837 : _GEN2239;
wire  _GEN5839 = io_x[37] ? _GEN4879 : _GEN5838;
wire  _GEN5840 = io_x[39] ? _GEN4887 : _GEN5839;
wire  _GEN5841 = io_x[72] ? _GEN5840 : _GEN5834;
wire  _GEN5842 = io_x[29] ? _GEN5841 : _GEN5005;
wire  _GEN5843 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5844 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN5845 = io_x[37] ? _GEN5844 : _GEN5843;
wire  _GEN5846 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5847 = io_x[37] ? _GEN5846 : _GEN4879;
wire  _GEN5848 = io_x[39] ? _GEN5847 : _GEN5845;
wire  _GEN5849 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5850 = io_x[17] ? _GEN5849 : _GEN1711;
wire  _GEN5851 = io_x[75] ? _GEN1899 : _GEN5850;
wire  _GEN5852 = io_x[25] ? _GEN5851 : _GEN2288;
wire  _GEN5853 = io_x[37] ? _GEN5852 : _GEN4879;
wire  _GEN5854 = io_x[39] ? _GEN4883 : _GEN5853;
wire  _GEN5855 = io_x[72] ? _GEN5854 : _GEN5848;
wire  _GEN5856 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5857 = io_x[17] ? _GEN5856 : _GEN1731;
wire  _GEN5858 = io_x[75] ? _GEN5857 : _GEN1903;
wire  _GEN5859 = io_x[25] ? _GEN5858 : _GEN2239;
wire  _GEN5860 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5861 = io_x[17] ? _GEN5860 : _GEN1731;
wire  _GEN5862 = io_x[75] ? _GEN1899 : _GEN5861;
wire  _GEN5863 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5864 = io_x[17] ? _GEN5863 : _GEN1731;
wire  _GEN5865 = io_x[75] ? _GEN1899 : _GEN5864;
wire  _GEN5866 = io_x[25] ? _GEN5865 : _GEN5862;
wire  _GEN5867 = io_x[37] ? _GEN5866 : _GEN5859;
wire  _GEN5868 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5869 = io_x[37] ? _GEN5868 : _GEN4885;
wire  _GEN5870 = io_x[39] ? _GEN5869 : _GEN5867;
wire  _GEN5871 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5872 = io_x[17] ? _GEN5871 : _GEN1731;
wire  _GEN5873 = io_x[75] ? _GEN1903 : _GEN5872;
wire  _GEN5874 = io_x[25] ? _GEN5873 : _GEN2239;
wire  _GEN5875 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5876 = io_x[17] ? _GEN5875 : _GEN1731;
wire  _GEN5877 = io_x[75] ? _GEN1903 : _GEN5876;
wire  _GEN5878 = io_x[25] ? _GEN5877 : _GEN2239;
wire  _GEN5879 = io_x[37] ? _GEN5878 : _GEN5874;
wire  _GEN5880 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5881 = io_x[75] ? _GEN1899 : _GEN5880;
wire  _GEN5882 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5883 = io_x[17] ? _GEN5882 : _GEN1731;
wire  _GEN5884 = io_x[75] ? _GEN1899 : _GEN5883;
wire  _GEN5885 = io_x[25] ? _GEN5884 : _GEN5881;
wire  _GEN5886 = io_x[37] ? _GEN4879 : _GEN5885;
wire  _GEN5887 = io_x[39] ? _GEN5886 : _GEN5879;
wire  _GEN5888 = io_x[72] ? _GEN5887 : _GEN5870;
wire  _GEN5889 = io_x[29] ? _GEN5888 : _GEN5855;
wire  _GEN5890 = io_x[18] ? _GEN5889 : _GEN5842;
wire  _GEN5891 = io_x[19] ? _GEN5890 : _GEN5827;
wire  _GEN5892 = io_x[24] ? _GEN5891 : _GEN5784;
wire  _GEN5893 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5894 = io_x[17] ? _GEN1731 : _GEN5893;
wire  _GEN5895 = io_x[75] ? _GEN1899 : _GEN5894;
wire  _GEN5896 = io_x[25] ? _GEN2288 : _GEN5895;
wire  _GEN5897 = io_x[37] ? _GEN5896 : _GEN4879;
wire  _GEN5898 = io_x[39] ? _GEN4883 : _GEN5897;
wire  _GEN5899 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5900 = io_x[25] ? _GEN2239 : _GEN5899;
wire  _GEN5901 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5902 = io_x[17] ? _GEN1731 : _GEN5901;
wire  _GEN5903 = io_x[75] ? _GEN1899 : _GEN5902;
wire  _GEN5904 = io_x[25] ? _GEN2288 : _GEN5903;
wire  _GEN5905 = io_x[37] ? _GEN5904 : _GEN5900;
wire  _GEN5906 = io_x[39] ? _GEN4883 : _GEN5905;
wire  _GEN5907 = io_x[72] ? _GEN5906 : _GEN5898;
wire  _GEN5908 = io_x[39] ? _GEN4887 : _GEN4883;
wire  _GEN5909 = io_x[72] ? _GEN4979 : _GEN5908;
wire  _GEN5910 = io_x[29] ? _GEN5909 : _GEN5907;
wire  _GEN5911 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN5912 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5913 = io_x[17] ? _GEN5912 : _GEN1731;
wire  _GEN5914 = io_x[75] ? _GEN1903 : _GEN5913;
wire  _GEN5915 = io_x[25] ? _GEN5914 : _GEN2288;
wire  _GEN5916 = io_x[37] ? _GEN5915 : _GEN4879;
wire  _GEN5917 = io_x[39] ? _GEN5916 : _GEN5911;
wire  _GEN5918 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5919 = io_x[25] ? _GEN2239 : _GEN5918;
wire  _GEN5920 = io_x[37] ? _GEN5919 : _GEN4879;
wire  _GEN5921 = io_x[39] ? _GEN4887 : _GEN5920;
wire  _GEN5922 = io_x[72] ? _GEN5921 : _GEN5917;
wire  _GEN5923 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN5924 = io_x[39] ? _GEN4887 : _GEN5923;
wire  _GEN5925 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5926 = io_x[25] ? _GEN2288 : _GEN5925;
wire  _GEN5927 = io_x[37] ? _GEN5926 : _GEN4879;
wire  _GEN5928 = io_x[39] ? _GEN5927 : _GEN4883;
wire  _GEN5929 = io_x[72] ? _GEN5928 : _GEN5924;
wire  _GEN5930 = io_x[29] ? _GEN5929 : _GEN5922;
wire  _GEN5931 = io_x[18] ? _GEN5930 : _GEN5910;
wire  _GEN5932 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN5933 = io_x[39] ? _GEN4883 : _GEN5932;
wire  _GEN5934 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5935 = io_x[75] ? _GEN1899 : _GEN5934;
wire  _GEN5936 = io_x[25] ? _GEN2288 : _GEN5935;
wire  _GEN5937 = io_x[37] ? _GEN4879 : _GEN5936;
wire  _GEN5938 = io_x[39] ? _GEN4883 : _GEN5937;
wire  _GEN5939 = io_x[72] ? _GEN5938 : _GEN5933;
wire  _GEN5940 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5941 = io_x[37] ? _GEN5940 : _GEN4879;
wire  _GEN5942 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5943 = io_x[17] ? _GEN5942 : _GEN1731;
wire  _GEN5944 = io_x[75] ? _GEN1903 : _GEN5943;
wire  _GEN5945 = io_x[25] ? _GEN5944 : _GEN2288;
wire  _GEN5946 = io_x[37] ? _GEN5945 : _GEN4879;
wire  _GEN5947 = io_x[39] ? _GEN5946 : _GEN5941;
wire  _GEN5948 = io_x[25] ? _GEN2239 : _GEN2288;
wire  _GEN5949 = io_x[37] ? _GEN4879 : _GEN5948;
wire  _GEN5950 = io_x[39] ? _GEN4883 : _GEN5949;
wire  _GEN5951 = io_x[72] ? _GEN5950 : _GEN5947;
wire  _GEN5952 = io_x[29] ? _GEN5951 : _GEN5939;
wire  _GEN5953 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5954 = io_x[17] ? _GEN1731 : _GEN5953;
wire  _GEN5955 = io_x[75] ? _GEN1899 : _GEN5954;
wire  _GEN5956 = io_x[25] ? _GEN2239 : _GEN5955;
wire  _GEN5957 = io_x[37] ? _GEN5956 : _GEN4885;
wire  _GEN5958 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN5959 = io_x[75] ? _GEN1899 : _GEN5958;
wire  _GEN5960 = io_x[25] ? _GEN5959 : _GEN2288;
wire  _GEN5961 = io_x[37] ? _GEN5960 : _GEN4885;
wire  _GEN5962 = io_x[39] ? _GEN5961 : _GEN5957;
wire  _GEN5963 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5964 = io_x[25] ? _GEN5963 : _GEN2288;
wire  _GEN5965 = io_x[37] ? _GEN4879 : _GEN5964;
wire  _GEN5966 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5967 = io_x[25] ? _GEN2288 : _GEN5966;
wire  _GEN5968 = io_x[37] ? _GEN4879 : _GEN5967;
wire  _GEN5969 = io_x[39] ? _GEN5968 : _GEN5965;
wire  _GEN5970 = io_x[72] ? _GEN5969 : _GEN5962;
wire  _GEN5971 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5972 = io_x[17] ? _GEN5971 : _GEN1731;
wire  _GEN5973 = io_x[75] ? _GEN1899 : _GEN5972;
wire  _GEN5974 = io_x[25] ? _GEN5973 : _GEN2288;
wire  _GEN5975 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5976 = io_x[17] ? _GEN1731 : _GEN5975;
wire  _GEN5977 = io_x[75] ? _GEN1899 : _GEN5976;
wire  _GEN5978 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN5979 = io_x[75] ? _GEN1899 : _GEN5978;
wire  _GEN5980 = io_x[25] ? _GEN5979 : _GEN5977;
wire  _GEN5981 = io_x[37] ? _GEN5980 : _GEN5974;
wire  _GEN5982 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN5983 = io_x[37] ? _GEN4879 : _GEN5982;
wire  _GEN5984 = io_x[39] ? _GEN5983 : _GEN5981;
wire  _GEN5985 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN5986 = io_x[17] ? _GEN5985 : _GEN1731;
wire  _GEN5987 = io_x[75] ? _GEN1899 : _GEN5986;
wire  _GEN5988 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN5989 = io_x[17] ? _GEN5988 : _GEN1731;
wire  _GEN5990 = io_x[75] ? _GEN1899 : _GEN5989;
wire  _GEN5991 = io_x[25] ? _GEN5990 : _GEN5987;
wire  _GEN5992 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN5993 = io_x[25] ? _GEN2239 : _GEN5992;
wire  _GEN5994 = io_x[37] ? _GEN5993 : _GEN5991;
wire  _GEN5995 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN5996 = io_x[25] ? _GEN5995 : _GEN2288;
wire  _GEN5997 = io_x[37] ? _GEN4885 : _GEN5996;
wire  _GEN5998 = io_x[39] ? _GEN5997 : _GEN5994;
wire  _GEN5999 = io_x[72] ? _GEN5998 : _GEN5984;
wire  _GEN6000 = io_x[29] ? _GEN5999 : _GEN5970;
wire  _GEN6001 = io_x[18] ? _GEN6000 : _GEN5952;
wire  _GEN6002 = io_x[19] ? _GEN6001 : _GEN5931;
wire  _GEN6003 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6004 = io_x[17] ? _GEN1731 : _GEN6003;
wire  _GEN6005 = io_x[75] ? _GEN6004 : _GEN1899;
wire  _GEN6006 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6007 = io_x[17] ? _GEN6006 : _GEN1731;
wire  _GEN6008 = io_x[75] ? _GEN6007 : _GEN1899;
wire  _GEN6009 = io_x[25] ? _GEN6008 : _GEN6005;
wire  _GEN6010 = io_x[37] ? _GEN4879 : _GEN6009;
wire  _GEN6011 = io_x[39] ? _GEN4883 : _GEN6010;
wire  _GEN6012 = io_x[72] ? _GEN6011 : _GEN4979;
wire  _GEN6013 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN6014 = io_x[75] ? _GEN1899 : _GEN6013;
wire  _GEN6015 = io_x[25] ? _GEN2288 : _GEN6014;
wire  _GEN6016 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6017 = io_x[17] ? _GEN1731 : _GEN6016;
wire  _GEN6018 = io_x[75] ? _GEN1899 : _GEN6017;
wire  _GEN6019 = io_x[25] ? _GEN2288 : _GEN6018;
wire  _GEN6020 = io_x[37] ? _GEN6019 : _GEN6015;
wire  _GEN6021 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN6022 = io_x[39] ? _GEN6021 : _GEN6020;
wire  _GEN6023 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN6024 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN6025 = io_x[39] ? _GEN6024 : _GEN6023;
wire  _GEN6026 = io_x[72] ? _GEN6025 : _GEN6022;
wire  _GEN6027 = io_x[29] ? _GEN6026 : _GEN6012;
wire  _GEN6028 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6029 = io_x[17] ? _GEN6028 : _GEN1731;
wire  _GEN6030 = io_x[75] ? _GEN1899 : _GEN6029;
wire  _GEN6031 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN6032 = io_x[75] ? _GEN1899 : _GEN6031;
wire  _GEN6033 = io_x[25] ? _GEN6032 : _GEN6030;
wire  _GEN6034 = io_x[37] ? _GEN6033 : _GEN4885;
wire  _GEN6035 = io_x[39] ? _GEN4883 : _GEN6034;
wire  _GEN6036 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6037 = io_x[17] ? _GEN6036 : _GEN1731;
wire  _GEN6038 = io_x[75] ? _GEN1903 : _GEN6037;
wire  _GEN6039 = io_x[25] ? _GEN6038 : _GEN2288;
wire  _GEN6040 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6041 = io_x[17] ? _GEN6040 : _GEN1731;
wire  _GEN6042 = io_x[75] ? _GEN1903 : _GEN6041;
wire  _GEN6043 = io_x[25] ? _GEN6042 : _GEN2288;
wire  _GEN6044 = io_x[37] ? _GEN6043 : _GEN6039;
wire  _GEN6045 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6046 = io_x[17] ? _GEN6045 : _GEN1731;
wire  _GEN6047 = io_x[75] ? _GEN6046 : _GEN1899;
wire  _GEN6048 = io_x[25] ? _GEN6047 : _GEN2288;
wire  _GEN6049 = io_x[37] ? _GEN6048 : _GEN4879;
wire  _GEN6050 = io_x[39] ? _GEN6049 : _GEN6044;
wire  _GEN6051 = io_x[72] ? _GEN6050 : _GEN6035;
wire  _GEN6052 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6053 = io_x[17] ? _GEN6052 : _GEN1731;
wire  _GEN6054 = io_x[75] ? _GEN1899 : _GEN6053;
wire  _GEN6055 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6056 = io_x[17] ? _GEN6055 : _GEN1731;
wire  _GEN6057 = io_x[75] ? _GEN1899 : _GEN6056;
wire  _GEN6058 = io_x[25] ? _GEN6057 : _GEN6054;
wire  _GEN6059 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6060 = io_x[17] ? _GEN6059 : _GEN1731;
wire  _GEN6061 = io_x[75] ? _GEN1899 : _GEN6060;
wire  _GEN6062 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6063 = io_x[17] ? _GEN6062 : _GEN1731;
wire  _GEN6064 = io_x[75] ? _GEN1899 : _GEN6063;
wire  _GEN6065 = io_x[25] ? _GEN6064 : _GEN6061;
wire  _GEN6066 = io_x[37] ? _GEN6065 : _GEN6058;
wire  _GEN6067 = io_x[39] ? _GEN4887 : _GEN6066;
wire  _GEN6068 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN6069 = io_x[25] ? _GEN6068 : _GEN2239;
wire  _GEN6070 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6071 = io_x[17] ? _GEN6070 : _GEN1731;
wire  _GEN6072 = io_x[75] ? _GEN1899 : _GEN6071;
wire  _GEN6073 = io_x[25] ? _GEN6072 : _GEN2239;
wire  _GEN6074 = io_x[37] ? _GEN6073 : _GEN6069;
wire  _GEN6075 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN6076 = io_x[25] ? _GEN6075 : _GEN2288;
wire  _GEN6077 = io_x[37] ? _GEN4879 : _GEN6076;
wire  _GEN6078 = io_x[39] ? _GEN6077 : _GEN6074;
wire  _GEN6079 = io_x[72] ? _GEN6078 : _GEN6067;
wire  _GEN6080 = io_x[29] ? _GEN6079 : _GEN6051;
wire  _GEN6081 = io_x[18] ? _GEN6080 : _GEN6027;
wire  _GEN6082 = io_x[37] ? _GEN4879 : _GEN4885;
wire  _GEN6083 = io_x[25] ? _GEN2288 : _GEN2239;
wire  _GEN6084 = io_x[37] ? _GEN6083 : _GEN4879;
wire  _GEN6085 = io_x[39] ? _GEN6084 : _GEN6082;
wire  _GEN6086 = io_x[72] ? _GEN4979 : _GEN6085;
wire  _GEN6087 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN6088 = io_x[75] ? _GEN1899 : _GEN6087;
wire  _GEN6089 = io_x[25] ? _GEN6088 : _GEN2288;
wire  _GEN6090 = io_x[37] ? _GEN6089 : _GEN4879;
wire  _GEN6091 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN6092 = io_x[75] ? _GEN6091 : _GEN1903;
wire  _GEN6093 = io_x[25] ? _GEN6092 : _GEN2288;
wire  _GEN6094 = io_x[37] ? _GEN6093 : _GEN4879;
wire  _GEN6095 = io_x[39] ? _GEN6094 : _GEN6090;
wire  _GEN6096 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN6097 = io_x[75] ? _GEN1899 : _GEN6096;
wire  _GEN6098 = io_x[25] ? _GEN6097 : _GEN2288;
wire  _GEN6099 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6100 = io_x[17] ? _GEN1731 : _GEN6099;
wire  _GEN6101 = io_x[75] ? _GEN6100 : _GEN1899;
wire  _GEN6102 = io_x[25] ? _GEN6101 : _GEN2288;
wire  _GEN6103 = io_x[37] ? _GEN6102 : _GEN6098;
wire  _GEN6104 = io_x[37] ? _GEN4885 : _GEN4879;
wire  _GEN6105 = io_x[39] ? _GEN6104 : _GEN6103;
wire  _GEN6106 = io_x[72] ? _GEN6105 : _GEN6095;
wire  _GEN6107 = io_x[29] ? _GEN6106 : _GEN6086;
wire  _GEN6108 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6109 = io_x[17] ? _GEN6108 : _GEN1731;
wire  _GEN6110 = io_x[75] ? _GEN1899 : _GEN6109;
wire  _GEN6111 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN6112 = io_x[75] ? _GEN1903 : _GEN6111;
wire  _GEN6113 = io_x[25] ? _GEN6112 : _GEN6110;
wire  _GEN6114 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6115 = io_x[17] ? _GEN6114 : _GEN1731;
wire  _GEN6116 = io_x[75] ? _GEN1899 : _GEN6115;
wire  _GEN6117 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6118 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6119 = io_x[17] ? _GEN6118 : _GEN6117;
wire  _GEN6120 = io_x[75] ? _GEN1903 : _GEN6119;
wire  _GEN6121 = io_x[25] ? _GEN6120 : _GEN6116;
wire  _GEN6122 = io_x[37] ? _GEN6121 : _GEN6113;
wire  _GEN6123 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN6124 = io_x[75] ? _GEN1899 : _GEN6123;
wire  _GEN6125 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN6126 = io_x[25] ? _GEN6125 : _GEN6124;
wire  _GEN6127 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6128 = io_x[17] ? _GEN1711 : _GEN6127;
wire  _GEN6129 = io_x[75] ? _GEN1899 : _GEN6128;
wire  _GEN6130 = io_x[25] ? _GEN6129 : _GEN2288;
wire  _GEN6131 = io_x[37] ? _GEN6130 : _GEN6126;
wire  _GEN6132 = io_x[39] ? _GEN6131 : _GEN6122;
wire  _GEN6133 = io_x[75] ? _GEN1903 : _GEN1899;
wire  _GEN6134 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6135 = io_x[17] ? _GEN6134 : _GEN1731;
wire  _GEN6136 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6137 = io_x[17] ? _GEN6136 : _GEN1731;
wire  _GEN6138 = io_x[75] ? _GEN6137 : _GEN6135;
wire  _GEN6139 = io_x[25] ? _GEN6138 : _GEN6133;
wire  _GEN6140 = io_x[75] ? _GEN1899 : _GEN1903;
wire  _GEN6141 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6142 = io_x[17] ? _GEN6141 : _GEN1711;
wire  _GEN6143 = io_x[75] ? _GEN6142 : _GEN1899;
wire  _GEN6144 = io_x[25] ? _GEN6143 : _GEN6140;
wire  _GEN6145 = io_x[37] ? _GEN6144 : _GEN6139;
wire  _GEN6146 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6147 = io_x[17] ? _GEN6146 : _GEN1731;
wire  _GEN6148 = io_x[75] ? _GEN1899 : _GEN6147;
wire  _GEN6149 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6150 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6151 = io_x[17] ? _GEN6150 : _GEN6149;
wire  _GEN6152 = io_x[75] ? _GEN1899 : _GEN6151;
wire  _GEN6153 = io_x[25] ? _GEN6152 : _GEN6148;
wire  _GEN6154 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6155 = io_x[17] ? _GEN6154 : _GEN1731;
wire  _GEN6156 = io_x[75] ? _GEN6155 : _GEN1899;
wire  _GEN6157 = io_x[25] ? _GEN6156 : _GEN2239;
wire  _GEN6158 = io_x[37] ? _GEN6157 : _GEN6153;
wire  _GEN6159 = io_x[39] ? _GEN6158 : _GEN6145;
wire  _GEN6160 = io_x[72] ? _GEN6159 : _GEN6132;
wire  _GEN6161 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6162 = io_x[17] ? _GEN6161 : _GEN1731;
wire  _GEN6163 = io_x[75] ? _GEN1903 : _GEN6162;
wire  _GEN6164 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6165 = io_x[17] ? _GEN6164 : _GEN1731;
wire  _GEN6166 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6167 = io_x[17] ? _GEN6166 : _GEN1731;
wire  _GEN6168 = io_x[75] ? _GEN6167 : _GEN6165;
wire  _GEN6169 = io_x[25] ? _GEN6168 : _GEN6163;
wire  _GEN6170 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6171 = io_x[17] ? _GEN6170 : _GEN1731;
wire  _GEN6172 = io_x[75] ? _GEN1903 : _GEN6171;
wire  _GEN6173 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6174 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6175 = io_x[17] ? _GEN6174 : _GEN6173;
wire  _GEN6176 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6177 = io_x[17] ? _GEN6176 : _GEN1711;
wire  _GEN6178 = io_x[75] ? _GEN6177 : _GEN6175;
wire  _GEN6179 = io_x[25] ? _GEN6178 : _GEN6172;
wire  _GEN6180 = io_x[37] ? _GEN6179 : _GEN6169;
wire  _GEN6181 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN6182 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN6183 = io_x[75] ? _GEN6182 : _GEN6181;
wire  _GEN6184 = io_x[25] ? _GEN6183 : _GEN2239;
wire  _GEN6185 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN6186 = io_x[75] ? _GEN1899 : _GEN6185;
wire  _GEN6187 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6188 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6189 = io_x[17] ? _GEN6188 : _GEN6187;
wire  _GEN6190 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6191 = io_x[17] ? _GEN6190 : _GEN1711;
wire  _GEN6192 = io_x[75] ? _GEN6191 : _GEN6189;
wire  _GEN6193 = io_x[25] ? _GEN6192 : _GEN6186;
wire  _GEN6194 = io_x[37] ? _GEN6193 : _GEN6184;
wire  _GEN6195 = io_x[39] ? _GEN6194 : _GEN6180;
wire  _GEN6196 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6197 = io_x[17] ? _GEN6196 : _GEN1731;
wire  _GEN6198 = io_x[75] ? _GEN1899 : _GEN6197;
wire  _GEN6199 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6200 = io_x[17] ? _GEN6199 : _GEN1731;
wire  _GEN6201 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6202 = io_x[17] ? _GEN6201 : _GEN1731;
wire  _GEN6203 = io_x[75] ? _GEN6202 : _GEN6200;
wire  _GEN6204 = io_x[25] ? _GEN6203 : _GEN6198;
wire  _GEN6205 = io_x[17] ? _GEN1731 : _GEN1711;
wire  _GEN6206 = io_x[75] ? _GEN1903 : _GEN6205;
wire  _GEN6207 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6208 = io_x[17] ? _GEN6207 : _GEN1711;
wire  _GEN6209 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6210 = io_x[17] ? _GEN6209 : _GEN1711;
wire  _GEN6211 = io_x[75] ? _GEN6210 : _GEN6208;
wire  _GEN6212 = io_x[25] ? _GEN6211 : _GEN6206;
wire  _GEN6213 = io_x[37] ? _GEN6212 : _GEN6204;
wire  _GEN6214 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6215 = io_x[17] ? _GEN6214 : _GEN1711;
wire  _GEN6216 = io_x[75] ? _GEN1899 : _GEN6215;
wire  _GEN6217 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6218 = io_x[17] ? _GEN6217 : _GEN1731;
wire  _GEN6219 = io_x[75] ? _GEN1903 : _GEN6218;
wire  _GEN6220 = io_x[25] ? _GEN6219 : _GEN6216;
wire  _GEN6221 = io_x[21] ? _GEN1698 : _GEN1699;
wire  _GEN6222 = io_x[17] ? _GEN6221 : _GEN1731;
wire  _GEN6223 = io_x[75] ? _GEN6222 : _GEN1899;
wire  _GEN6224 = io_x[17] ? _GEN1711 : _GEN1731;
wire  _GEN6225 = io_x[21] ? _GEN1699 : _GEN1698;
wire  _GEN6226 = io_x[17] ? _GEN6225 : _GEN1731;
wire  _GEN6227 = io_x[75] ? _GEN6226 : _GEN6224;
wire  _GEN6228 = io_x[25] ? _GEN6227 : _GEN6223;
wire  _GEN6229 = io_x[37] ? _GEN6228 : _GEN6220;
wire  _GEN6230 = io_x[39] ? _GEN6229 : _GEN6213;
wire  _GEN6231 = io_x[72] ? _GEN6230 : _GEN6195;
wire  _GEN6232 = io_x[29] ? _GEN6231 : _GEN6160;
wire  _GEN6233 = io_x[18] ? _GEN6232 : _GEN6107;
wire  _GEN6234 = io_x[19] ? _GEN6233 : _GEN6081;
wire  _GEN6235 = io_x[24] ? _GEN6234 : _GEN6002;
wire  _GEN6236 = io_x[23] ? _GEN6235 : _GEN5892;
wire  _GEN6237 = io_x[33] ? _GEN6236 : _GEN5675;
wire  _GEN6238 = io_x[32] ? _GEN6237 : _GEN5293;
assign io_y[16] = _GEN6238;
wire  _GEN6239 = 1'b0;
wire  _GEN6240 = 1'b1;
wire  _GEN6241 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6242 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6243 = io_x[20] ? _GEN6242 : _GEN6241;
wire  _GEN6244 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6245 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6246 = io_x[20] ? _GEN6245 : _GEN6244;
wire  _GEN6247 = io_x[28] ? _GEN6246 : _GEN6243;
wire  _GEN6248 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6249 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6250 = io_x[20] ? _GEN6249 : _GEN6248;
wire  _GEN6251 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6252 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6253 = io_x[20] ? _GEN6252 : _GEN6251;
wire  _GEN6254 = io_x[28] ? _GEN6253 : _GEN6250;
wire  _GEN6255 = io_x[24] ? _GEN6254 : _GEN6247;
wire  _GEN6256 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6257 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6258 = io_x[20] ? _GEN6257 : _GEN6256;
wire  _GEN6259 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6260 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6261 = io_x[20] ? _GEN6260 : _GEN6259;
wire  _GEN6262 = io_x[28] ? _GEN6261 : _GEN6258;
wire  _GEN6263 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6264 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6265 = io_x[20] ? _GEN6264 : _GEN6263;
wire  _GEN6266 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6267 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6268 = io_x[20] ? _GEN6267 : _GEN6266;
wire  _GEN6269 = io_x[28] ? _GEN6268 : _GEN6265;
wire  _GEN6270 = io_x[24] ? _GEN6269 : _GEN6262;
wire  _GEN6271 = io_x[18] ? _GEN6270 : _GEN6255;
wire  _GEN6272 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6273 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6274 = io_x[20] ? _GEN6273 : _GEN6272;
wire  _GEN6275 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6276 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6277 = io_x[20] ? _GEN6276 : _GEN6275;
wire  _GEN6278 = io_x[28] ? _GEN6277 : _GEN6274;
wire  _GEN6279 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6280 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6281 = io_x[20] ? _GEN6280 : _GEN6279;
wire  _GEN6282 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6283 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6284 = io_x[20] ? _GEN6283 : _GEN6282;
wire  _GEN6285 = io_x[28] ? _GEN6284 : _GEN6281;
wire  _GEN6286 = io_x[24] ? _GEN6285 : _GEN6278;
wire  _GEN6287 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6288 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6289 = io_x[20] ? _GEN6288 : _GEN6287;
wire  _GEN6290 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6291 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6292 = io_x[20] ? _GEN6291 : _GEN6290;
wire  _GEN6293 = io_x[28] ? _GEN6292 : _GEN6289;
wire  _GEN6294 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6295 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6296 = io_x[20] ? _GEN6295 : _GEN6294;
wire  _GEN6297 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6298 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6299 = io_x[20] ? _GEN6298 : _GEN6297;
wire  _GEN6300 = io_x[28] ? _GEN6299 : _GEN6296;
wire  _GEN6301 = io_x[24] ? _GEN6300 : _GEN6293;
wire  _GEN6302 = io_x[18] ? _GEN6301 : _GEN6286;
wire  _GEN6303 = io_x[74] ? _GEN6302 : _GEN6271;
wire  _GEN6304 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6305 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6306 = io_x[20] ? _GEN6305 : _GEN6304;
wire  _GEN6307 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6308 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6309 = io_x[20] ? _GEN6308 : _GEN6307;
wire  _GEN6310 = io_x[28] ? _GEN6309 : _GEN6306;
wire  _GEN6311 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6312 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6313 = io_x[20] ? _GEN6312 : _GEN6311;
wire  _GEN6314 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6315 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6316 = io_x[20] ? _GEN6315 : _GEN6314;
wire  _GEN6317 = io_x[28] ? _GEN6316 : _GEN6313;
wire  _GEN6318 = io_x[24] ? _GEN6317 : _GEN6310;
wire  _GEN6319 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6320 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6321 = io_x[20] ? _GEN6320 : _GEN6319;
wire  _GEN6322 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6323 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6324 = io_x[20] ? _GEN6323 : _GEN6322;
wire  _GEN6325 = io_x[28] ? _GEN6324 : _GEN6321;
wire  _GEN6326 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6327 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6328 = io_x[20] ? _GEN6327 : _GEN6326;
wire  _GEN6329 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6330 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6331 = io_x[20] ? _GEN6330 : _GEN6329;
wire  _GEN6332 = io_x[28] ? _GEN6331 : _GEN6328;
wire  _GEN6333 = io_x[24] ? _GEN6332 : _GEN6325;
wire  _GEN6334 = io_x[18] ? _GEN6333 : _GEN6318;
wire  _GEN6335 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6336 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6337 = io_x[20] ? _GEN6336 : _GEN6335;
wire  _GEN6338 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6339 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6340 = io_x[20] ? _GEN6339 : _GEN6338;
wire  _GEN6341 = io_x[28] ? _GEN6340 : _GEN6337;
wire  _GEN6342 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6343 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6344 = io_x[20] ? _GEN6343 : _GEN6342;
wire  _GEN6345 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6346 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6347 = io_x[20] ? _GEN6346 : _GEN6345;
wire  _GEN6348 = io_x[28] ? _GEN6347 : _GEN6344;
wire  _GEN6349 = io_x[24] ? _GEN6348 : _GEN6341;
wire  _GEN6350 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6351 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6352 = io_x[20] ? _GEN6351 : _GEN6350;
wire  _GEN6353 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6354 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6355 = io_x[20] ? _GEN6354 : _GEN6353;
wire  _GEN6356 = io_x[28] ? _GEN6355 : _GEN6352;
wire  _GEN6357 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6358 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6359 = io_x[20] ? _GEN6358 : _GEN6357;
wire  _GEN6360 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6361 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6362 = io_x[20] ? _GEN6361 : _GEN6360;
wire  _GEN6363 = io_x[28] ? _GEN6362 : _GEN6359;
wire  _GEN6364 = io_x[24] ? _GEN6363 : _GEN6356;
wire  _GEN6365 = io_x[18] ? _GEN6364 : _GEN6349;
wire  _GEN6366 = io_x[74] ? _GEN6365 : _GEN6334;
wire  _GEN6367 = io_x[75] ? _GEN6366 : _GEN6303;
wire  _GEN6368 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6369 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6370 = io_x[20] ? _GEN6369 : _GEN6368;
wire  _GEN6371 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6372 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6373 = io_x[20] ? _GEN6372 : _GEN6371;
wire  _GEN6374 = io_x[28] ? _GEN6373 : _GEN6370;
wire  _GEN6375 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6376 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6377 = io_x[20] ? _GEN6376 : _GEN6375;
wire  _GEN6378 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6379 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6380 = io_x[20] ? _GEN6379 : _GEN6378;
wire  _GEN6381 = io_x[28] ? _GEN6380 : _GEN6377;
wire  _GEN6382 = io_x[24] ? _GEN6381 : _GEN6374;
wire  _GEN6383 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6384 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6385 = io_x[20] ? _GEN6384 : _GEN6383;
wire  _GEN6386 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6387 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6388 = io_x[20] ? _GEN6387 : _GEN6386;
wire  _GEN6389 = io_x[28] ? _GEN6388 : _GEN6385;
wire  _GEN6390 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6391 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6392 = io_x[20] ? _GEN6391 : _GEN6390;
wire  _GEN6393 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6394 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6395 = io_x[20] ? _GEN6394 : _GEN6393;
wire  _GEN6396 = io_x[28] ? _GEN6395 : _GEN6392;
wire  _GEN6397 = io_x[24] ? _GEN6396 : _GEN6389;
wire  _GEN6398 = io_x[18] ? _GEN6397 : _GEN6382;
wire  _GEN6399 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6400 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6401 = io_x[20] ? _GEN6400 : _GEN6399;
wire  _GEN6402 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6403 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6404 = io_x[20] ? _GEN6403 : _GEN6402;
wire  _GEN6405 = io_x[28] ? _GEN6404 : _GEN6401;
wire  _GEN6406 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6407 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6408 = io_x[20] ? _GEN6407 : _GEN6406;
wire  _GEN6409 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6410 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6411 = io_x[20] ? _GEN6410 : _GEN6409;
wire  _GEN6412 = io_x[28] ? _GEN6411 : _GEN6408;
wire  _GEN6413 = io_x[24] ? _GEN6412 : _GEN6405;
wire  _GEN6414 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6415 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6416 = io_x[20] ? _GEN6415 : _GEN6414;
wire  _GEN6417 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6418 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6419 = io_x[20] ? _GEN6418 : _GEN6417;
wire  _GEN6420 = io_x[28] ? _GEN6419 : _GEN6416;
wire  _GEN6421 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6422 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6423 = io_x[20] ? _GEN6422 : _GEN6421;
wire  _GEN6424 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6425 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6426 = io_x[20] ? _GEN6425 : _GEN6424;
wire  _GEN6427 = io_x[28] ? _GEN6426 : _GEN6423;
wire  _GEN6428 = io_x[24] ? _GEN6427 : _GEN6420;
wire  _GEN6429 = io_x[18] ? _GEN6428 : _GEN6413;
wire  _GEN6430 = io_x[74] ? _GEN6429 : _GEN6398;
wire  _GEN6431 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6432 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6433 = io_x[20] ? _GEN6432 : _GEN6431;
wire  _GEN6434 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6435 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6436 = io_x[20] ? _GEN6435 : _GEN6434;
wire  _GEN6437 = io_x[28] ? _GEN6436 : _GEN6433;
wire  _GEN6438 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6439 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6440 = io_x[20] ? _GEN6439 : _GEN6438;
wire  _GEN6441 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6442 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6443 = io_x[20] ? _GEN6442 : _GEN6441;
wire  _GEN6444 = io_x[28] ? _GEN6443 : _GEN6440;
wire  _GEN6445 = io_x[24] ? _GEN6444 : _GEN6437;
wire  _GEN6446 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6447 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6448 = io_x[20] ? _GEN6447 : _GEN6446;
wire  _GEN6449 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6450 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6451 = io_x[20] ? _GEN6450 : _GEN6449;
wire  _GEN6452 = io_x[28] ? _GEN6451 : _GEN6448;
wire  _GEN6453 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6454 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6455 = io_x[20] ? _GEN6454 : _GEN6453;
wire  _GEN6456 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6457 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6458 = io_x[20] ? _GEN6457 : _GEN6456;
wire  _GEN6459 = io_x[28] ? _GEN6458 : _GEN6455;
wire  _GEN6460 = io_x[24] ? _GEN6459 : _GEN6452;
wire  _GEN6461 = io_x[18] ? _GEN6460 : _GEN6445;
wire  _GEN6462 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6463 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6464 = io_x[20] ? _GEN6463 : _GEN6462;
wire  _GEN6465 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6466 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6467 = io_x[20] ? _GEN6466 : _GEN6465;
wire  _GEN6468 = io_x[28] ? _GEN6467 : _GEN6464;
wire  _GEN6469 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6470 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6471 = io_x[20] ? _GEN6470 : _GEN6469;
wire  _GEN6472 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6473 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6474 = io_x[20] ? _GEN6473 : _GEN6472;
wire  _GEN6475 = io_x[28] ? _GEN6474 : _GEN6471;
wire  _GEN6476 = io_x[24] ? _GEN6475 : _GEN6468;
wire  _GEN6477 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6478 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6479 = io_x[20] ? _GEN6478 : _GEN6477;
wire  _GEN6480 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6481 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6482 = io_x[20] ? _GEN6481 : _GEN6480;
wire  _GEN6483 = io_x[28] ? _GEN6482 : _GEN6479;
wire  _GEN6484 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6485 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6486 = io_x[20] ? _GEN6485 : _GEN6484;
wire  _GEN6487 = io_x[16] ? _GEN6239 : _GEN6240;
wire  _GEN6488 = io_x[16] ? _GEN6240 : _GEN6239;
wire  _GEN6489 = io_x[20] ? _GEN6488 : _GEN6487;
wire  _GEN6490 = io_x[28] ? _GEN6489 : _GEN6486;
wire  _GEN6491 = io_x[24] ? _GEN6490 : _GEN6483;
wire  _GEN6492 = io_x[18] ? _GEN6491 : _GEN6476;
wire  _GEN6493 = io_x[74] ? _GEN6492 : _GEN6461;
wire  _GEN6494 = io_x[75] ? _GEN6493 : _GEN6430;
wire  _GEN6495 = io_x[72] ? _GEN6494 : _GEN6367;
assign io_y[15] = _GEN6495;
wire  _GEN6496 = 1'b0;
wire  _GEN6497 = 1'b1;
wire  _GEN6498 = io_x[73] ? _GEN6497 : _GEN6496;
assign io_y[14] = _GEN6498;
wire  _GEN6499 = 1'b0;
wire  _GEN6500 = 1'b1;
wire  _GEN6501 = io_x[72] ? _GEN6500 : _GEN6499;
wire  _GEN6502 = io_x[72] ? _GEN6500 : _GEN6499;
wire  _GEN6503 = io_x[39] ? _GEN6502 : _GEN6501;
wire  _GEN6504 = io_x[72] ? _GEN6500 : _GEN6499;
wire  _GEN6505 = io_x[72] ? _GEN6500 : _GEN6499;
wire  _GEN6506 = io_x[39] ? _GEN6505 : _GEN6504;
wire  _GEN6507 = io_x[69] ? _GEN6506 : _GEN6503;
assign io_y[13] = _GEN6507;
wire  _GEN6508 = 1'b0;
wire  _GEN6509 = 1'b1;
wire  _GEN6510 = io_x[71] ? _GEN6509 : _GEN6508;
wire  _GEN6511 = io_x[71] ? _GEN6509 : _GEN6508;
wire  _GEN6512 = io_x[69] ? _GEN6511 : _GEN6510;
assign io_y[12] = _GEN6512;
wire  _GEN6513 = 1'b0;
wire  _GEN6514 = 1'b1;
wire  _GEN6515 = io_x[70] ? _GEN6514 : _GEN6513;
assign io_y[11] = _GEN6515;
wire  _GEN6516 = 1'b0;
wire  _GEN6517 = 1'b1;
wire  _GEN6518 = io_x[69] ? _GEN6517 : _GEN6516;
wire  _GEN6519 = io_x[69] ? _GEN6517 : _GEN6516;
wire  _GEN6520 = io_x[70] ? _GEN6519 : _GEN6518;
wire  _GEN6521 = io_x[69] ? _GEN6517 : _GEN6516;
wire  _GEN6522 = io_x[69] ? _GEN6517 : _GEN6516;
wire  _GEN6523 = io_x[70] ? _GEN6522 : _GEN6521;
wire  _GEN6524 = io_x[39] ? _GEN6523 : _GEN6520;
wire  _GEN6525 = io_x[69] ? _GEN6517 : _GEN6516;
wire  _GEN6526 = io_x[69] ? _GEN6517 : _GEN6516;
wire  _GEN6527 = io_x[70] ? _GEN6526 : _GEN6525;
wire  _GEN6528 = io_x[69] ? _GEN6517 : _GEN6516;
wire  _GEN6529 = io_x[69] ? _GEN6517 : _GEN6516;
wire  _GEN6530 = io_x[70] ? _GEN6529 : _GEN6528;
wire  _GEN6531 = io_x[39] ? _GEN6530 : _GEN6527;
wire  _GEN6532 = io_x[72] ? _GEN6531 : _GEN6524;
assign io_y[10] = _GEN6532;
wire  _GEN6533 = 1'b1;
wire  _GEN6534 = 1'b0;
wire  _GEN6535 = 1'b1;
wire  _GEN6536 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6537 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6538 = io_x[11] ? _GEN6537 : _GEN6536;
wire  _GEN6539 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6540 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6541 = io_x[11] ? _GEN6540 : _GEN6539;
wire  _GEN6542 = io_x[15] ? _GEN6541 : _GEN6538;
wire  _GEN6543 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6544 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6545 = io_x[11] ? _GEN6544 : _GEN6543;
wire  _GEN6546 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6547 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6548 = io_x[11] ? _GEN6547 : _GEN6546;
wire  _GEN6549 = io_x[15] ? _GEN6548 : _GEN6545;
wire  _GEN6550 = io_x[3] ? _GEN6549 : _GEN6542;
wire  _GEN6551 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6552 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6553 = io_x[11] ? _GEN6552 : _GEN6551;
wire  _GEN6554 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6555 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6556 = io_x[11] ? _GEN6555 : _GEN6554;
wire  _GEN6557 = io_x[15] ? _GEN6556 : _GEN6553;
wire  _GEN6558 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6559 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6560 = io_x[11] ? _GEN6559 : _GEN6558;
wire  _GEN6561 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6562 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6563 = io_x[11] ? _GEN6562 : _GEN6561;
wire  _GEN6564 = io_x[15] ? _GEN6563 : _GEN6560;
wire  _GEN6565 = io_x[3] ? _GEN6564 : _GEN6557;
wire  _GEN6566 = io_x[24] ? _GEN6565 : _GEN6550;
wire  _GEN6567 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6568 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6569 = io_x[11] ? _GEN6568 : _GEN6567;
wire  _GEN6570 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6571 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6572 = io_x[11] ? _GEN6571 : _GEN6570;
wire  _GEN6573 = io_x[15] ? _GEN6572 : _GEN6569;
wire  _GEN6574 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6575 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6576 = io_x[11] ? _GEN6575 : _GEN6574;
wire  _GEN6577 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6578 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6579 = io_x[11] ? _GEN6578 : _GEN6577;
wire  _GEN6580 = io_x[15] ? _GEN6579 : _GEN6576;
wire  _GEN6581 = io_x[3] ? _GEN6580 : _GEN6573;
wire  _GEN6582 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6583 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6584 = io_x[11] ? _GEN6583 : _GEN6582;
wire  _GEN6585 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6586 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6587 = io_x[11] ? _GEN6586 : _GEN6585;
wire  _GEN6588 = io_x[15] ? _GEN6587 : _GEN6584;
wire  _GEN6589 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6590 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6591 = io_x[11] ? _GEN6590 : _GEN6589;
wire  _GEN6592 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6593 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6594 = io_x[11] ? _GEN6593 : _GEN6592;
wire  _GEN6595 = io_x[15] ? _GEN6594 : _GEN6591;
wire  _GEN6596 = io_x[3] ? _GEN6595 : _GEN6588;
wire  _GEN6597 = io_x[24] ? _GEN6596 : _GEN6581;
wire  _GEN6598 = io_x[33] ? _GEN6597 : _GEN6566;
wire  _GEN6599 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6600 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6601 = io_x[11] ? _GEN6600 : _GEN6599;
wire  _GEN6602 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6603 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6604 = io_x[11] ? _GEN6603 : _GEN6602;
wire  _GEN6605 = io_x[15] ? _GEN6604 : _GEN6601;
wire  _GEN6606 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6607 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6608 = io_x[11] ? _GEN6607 : _GEN6606;
wire  _GEN6609 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6610 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6611 = io_x[11] ? _GEN6610 : _GEN6609;
wire  _GEN6612 = io_x[15] ? _GEN6611 : _GEN6608;
wire  _GEN6613 = io_x[3] ? _GEN6612 : _GEN6605;
wire  _GEN6614 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6615 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6616 = io_x[11] ? _GEN6615 : _GEN6614;
wire  _GEN6617 = 1'b0;
wire  _GEN6618 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6619 = io_x[11] ? _GEN6618 : _GEN6617;
wire  _GEN6620 = io_x[15] ? _GEN6619 : _GEN6616;
wire  _GEN6621 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6622 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6623 = io_x[11] ? _GEN6622 : _GEN6621;
wire  _GEN6624 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6625 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6626 = io_x[11] ? _GEN6625 : _GEN6624;
wire  _GEN6627 = io_x[15] ? _GEN6626 : _GEN6623;
wire  _GEN6628 = io_x[3] ? _GEN6627 : _GEN6620;
wire  _GEN6629 = io_x[24] ? _GEN6628 : _GEN6613;
wire  _GEN6630 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6631 = io_x[11] ? _GEN6630 : _GEN6617;
wire  _GEN6632 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6633 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6634 = io_x[11] ? _GEN6633 : _GEN6632;
wire  _GEN6635 = io_x[15] ? _GEN6634 : _GEN6631;
wire  _GEN6636 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6637 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6638 = io_x[11] ? _GEN6637 : _GEN6636;
wire  _GEN6639 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6640 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6641 = io_x[11] ? _GEN6640 : _GEN6639;
wire  _GEN6642 = io_x[15] ? _GEN6641 : _GEN6638;
wire  _GEN6643 = io_x[3] ? _GEN6642 : _GEN6635;
wire  _GEN6644 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6645 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6646 = io_x[11] ? _GEN6645 : _GEN6644;
wire  _GEN6647 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6648 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6649 = io_x[11] ? _GEN6648 : _GEN6647;
wire  _GEN6650 = io_x[15] ? _GEN6649 : _GEN6646;
wire  _GEN6651 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6652 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6653 = io_x[11] ? _GEN6652 : _GEN6651;
wire  _GEN6654 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6655 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6656 = io_x[11] ? _GEN6655 : _GEN6654;
wire  _GEN6657 = io_x[15] ? _GEN6656 : _GEN6653;
wire  _GEN6658 = io_x[3] ? _GEN6657 : _GEN6650;
wire  _GEN6659 = io_x[24] ? _GEN6658 : _GEN6643;
wire  _GEN6660 = io_x[33] ? _GEN6659 : _GEN6629;
wire  _GEN6661 = io_x[81] ? _GEN6660 : _GEN6598;
wire  _GEN6662 = 1'b1;
wire  _GEN6663 = io_x[82] ? _GEN6662 : _GEN6661;
wire  _GEN6664 = 1'b1;
wire  _GEN6665 = io_x[83] ? _GEN6664 : _GEN6663;
wire  _GEN6666 = 1'b1;
wire  _GEN6667 = io_x[84] ? _GEN6666 : _GEN6665;
wire  _GEN6668 = 1'b1;
wire  _GEN6669 = io_x[85] ? _GEN6668 : _GEN6667;
wire  _GEN6670 = 1'b1;
wire  _GEN6671 = io_x[86] ? _GEN6670 : _GEN6669;
wire  _GEN6672 = 1'b1;
wire  _GEN6673 = io_x[87] ? _GEN6672 : _GEN6671;
wire  _GEN6674 = 1'b1;
wire  _GEN6675 = io_x[88] ? _GEN6674 : _GEN6673;
wire  _GEN6676 = 1'b1;
wire  _GEN6677 = io_x[89] ? _GEN6676 : _GEN6675;
wire  _GEN6678 = 1'b1;
wire  _GEN6679 = io_x[90] ? _GEN6678 : _GEN6677;
wire  _GEN6680 = 1'b1;
wire  _GEN6681 = io_x[91] ? _GEN6680 : _GEN6679;
wire  _GEN6682 = 1'b1;
wire  _GEN6683 = io_x[92] ? _GEN6682 : _GEN6681;
wire  _GEN6684 = 1'b1;
wire  _GEN6685 = io_x[93] ? _GEN6684 : _GEN6683;
wire  _GEN6686 = 1'b1;
wire  _GEN6687 = io_x[94] ? _GEN6686 : _GEN6685;
wire  _GEN6688 = 1'b1;
wire  _GEN6689 = io_x[95] ? _GEN6688 : _GEN6687;
wire  _GEN6690 = 1'b1;
wire  _GEN6691 = io_x[96] ? _GEN6690 : _GEN6689;
wire  _GEN6692 = 1'b1;
wire  _GEN6693 = io_x[97] ? _GEN6692 : _GEN6691;
wire  _GEN6694 = io_x[98] ? _GEN6693 : _GEN6533;
wire  _GEN6695 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6696 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6697 = io_x[11] ? _GEN6696 : _GEN6695;
wire  _GEN6698 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6699 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6700 = io_x[11] ? _GEN6699 : _GEN6698;
wire  _GEN6701 = io_x[15] ? _GEN6700 : _GEN6697;
wire  _GEN6702 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6703 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6704 = io_x[11] ? _GEN6703 : _GEN6702;
wire  _GEN6705 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6706 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6707 = io_x[11] ? _GEN6706 : _GEN6705;
wire  _GEN6708 = io_x[15] ? _GEN6707 : _GEN6704;
wire  _GEN6709 = io_x[3] ? _GEN6708 : _GEN6701;
wire  _GEN6710 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6711 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6712 = io_x[11] ? _GEN6711 : _GEN6710;
wire  _GEN6713 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6714 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6715 = io_x[11] ? _GEN6714 : _GEN6713;
wire  _GEN6716 = io_x[15] ? _GEN6715 : _GEN6712;
wire  _GEN6717 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6718 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6719 = io_x[11] ? _GEN6718 : _GEN6717;
wire  _GEN6720 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6721 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6722 = io_x[11] ? _GEN6721 : _GEN6720;
wire  _GEN6723 = io_x[15] ? _GEN6722 : _GEN6719;
wire  _GEN6724 = io_x[3] ? _GEN6723 : _GEN6716;
wire  _GEN6725 = io_x[24] ? _GEN6724 : _GEN6709;
wire  _GEN6726 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6727 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6728 = io_x[11] ? _GEN6727 : _GEN6726;
wire  _GEN6729 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6730 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6731 = io_x[11] ? _GEN6730 : _GEN6729;
wire  _GEN6732 = io_x[15] ? _GEN6731 : _GEN6728;
wire  _GEN6733 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6734 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6735 = io_x[11] ? _GEN6734 : _GEN6733;
wire  _GEN6736 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6737 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6738 = io_x[11] ? _GEN6737 : _GEN6736;
wire  _GEN6739 = io_x[15] ? _GEN6738 : _GEN6735;
wire  _GEN6740 = io_x[3] ? _GEN6739 : _GEN6732;
wire  _GEN6741 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6742 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6743 = io_x[11] ? _GEN6742 : _GEN6741;
wire  _GEN6744 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6745 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6746 = io_x[11] ? _GEN6745 : _GEN6744;
wire  _GEN6747 = io_x[15] ? _GEN6746 : _GEN6743;
wire  _GEN6748 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6749 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6750 = io_x[11] ? _GEN6749 : _GEN6748;
wire  _GEN6751 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6752 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6753 = io_x[11] ? _GEN6752 : _GEN6751;
wire  _GEN6754 = io_x[15] ? _GEN6753 : _GEN6750;
wire  _GEN6755 = io_x[3] ? _GEN6754 : _GEN6747;
wire  _GEN6756 = io_x[24] ? _GEN6755 : _GEN6740;
wire  _GEN6757 = io_x[33] ? _GEN6756 : _GEN6725;
wire  _GEN6758 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6759 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6760 = io_x[11] ? _GEN6759 : _GEN6758;
wire  _GEN6761 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6762 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6763 = io_x[11] ? _GEN6762 : _GEN6761;
wire  _GEN6764 = io_x[15] ? _GEN6763 : _GEN6760;
wire  _GEN6765 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6766 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6767 = io_x[11] ? _GEN6766 : _GEN6765;
wire  _GEN6768 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6769 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6770 = io_x[11] ? _GEN6769 : _GEN6768;
wire  _GEN6771 = io_x[15] ? _GEN6770 : _GEN6767;
wire  _GEN6772 = io_x[3] ? _GEN6771 : _GEN6764;
wire  _GEN6773 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6774 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6775 = io_x[11] ? _GEN6774 : _GEN6773;
wire  _GEN6776 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6777 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6778 = io_x[11] ? _GEN6777 : _GEN6776;
wire  _GEN6779 = io_x[15] ? _GEN6778 : _GEN6775;
wire  _GEN6780 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6781 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6782 = io_x[11] ? _GEN6781 : _GEN6780;
wire  _GEN6783 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6784 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6785 = io_x[11] ? _GEN6784 : _GEN6783;
wire  _GEN6786 = io_x[15] ? _GEN6785 : _GEN6782;
wire  _GEN6787 = io_x[3] ? _GEN6786 : _GEN6779;
wire  _GEN6788 = io_x[24] ? _GEN6787 : _GEN6772;
wire  _GEN6789 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6790 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6791 = io_x[11] ? _GEN6790 : _GEN6789;
wire  _GEN6792 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6793 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6794 = io_x[11] ? _GEN6793 : _GEN6792;
wire  _GEN6795 = io_x[15] ? _GEN6794 : _GEN6791;
wire  _GEN6796 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6797 = 1'b1;
wire  _GEN6798 = io_x[11] ? _GEN6797 : _GEN6796;
wire  _GEN6799 = io_x[11] ? _GEN6617 : _GEN6797;
wire  _GEN6800 = io_x[15] ? _GEN6799 : _GEN6798;
wire  _GEN6801 = io_x[3] ? _GEN6800 : _GEN6795;
wire  _GEN6802 = io_x[7] ? _GEN6534 : _GEN6535;
wire  _GEN6803 = io_x[11] ? _GEN6797 : _GEN6802;
wire  _GEN6804 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6805 = io_x[11] ? _GEN6617 : _GEN6804;
wire  _GEN6806 = io_x[15] ? _GEN6805 : _GEN6803;
wire  _GEN6807 = io_x[7] ? _GEN6535 : _GEN6534;
wire  _GEN6808 = io_x[11] ? _GEN6617 : _GEN6807;
wire  _GEN6809 = io_x[11] ? _GEN6797 : _GEN6617;
wire  _GEN6810 = io_x[15] ? _GEN6809 : _GEN6808;
wire  _GEN6811 = io_x[3] ? _GEN6810 : _GEN6806;
wire  _GEN6812 = io_x[24] ? _GEN6811 : _GEN6801;
wire  _GEN6813 = io_x[33] ? _GEN6812 : _GEN6788;
wire  _GEN6814 = io_x[81] ? _GEN6813 : _GEN6757;
wire  _GEN6815 = io_x[82] ? _GEN6662 : _GEN6814;
wire  _GEN6816 = io_x[83] ? _GEN6664 : _GEN6815;
wire  _GEN6817 = io_x[84] ? _GEN6666 : _GEN6816;
wire  _GEN6818 = io_x[85] ? _GEN6668 : _GEN6817;
wire  _GEN6819 = io_x[86] ? _GEN6670 : _GEN6818;
wire  _GEN6820 = io_x[87] ? _GEN6672 : _GEN6819;
wire  _GEN6821 = io_x[88] ? _GEN6674 : _GEN6820;
wire  _GEN6822 = io_x[89] ? _GEN6676 : _GEN6821;
wire  _GEN6823 = io_x[90] ? _GEN6678 : _GEN6822;
wire  _GEN6824 = io_x[91] ? _GEN6680 : _GEN6823;
wire  _GEN6825 = io_x[92] ? _GEN6682 : _GEN6824;
wire  _GEN6826 = io_x[93] ? _GEN6684 : _GEN6825;
wire  _GEN6827 = io_x[94] ? _GEN6686 : _GEN6826;
wire  _GEN6828 = io_x[95] ? _GEN6688 : _GEN6827;
wire  _GEN6829 = io_x[96] ? _GEN6690 : _GEN6828;
wire  _GEN6830 = io_x[97] ? _GEN6692 : _GEN6829;
wire  _GEN6831 = io_x[98] ? _GEN6830 : _GEN6533;
wire  _GEN6832 = io_x[45] ? _GEN6831 : _GEN6694;
assign io_y[9] = _GEN6832;
wire  _GEN6833 = 1'b0;
wire  _GEN6834 = 1'b1;
wire  _GEN6835 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN6836 = 1'b1;
wire  _GEN6837 = 1'b1;
wire  _GEN6838 = 1'b0;
wire  _GEN6839 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN6840 = 1'b0;
wire  _GEN6841 = io_x[6] ? _GEN6840 : _GEN6839;
wire  _GEN6842 = io_x[41] ? _GEN6841 : _GEN6836;
wire  _GEN6843 = 1'b1;
wire  _GEN6844 = io_x[14] ? _GEN6843 : _GEN6842;
wire  _GEN6845 = 1'b1;
wire  _GEN6846 = io_x[0] ? _GEN6845 : _GEN6844;
wire  _GEN6847 = io_x[76] ? _GEN6833 : _GEN6846;
wire  _GEN6848 = io_x[42] ? _GEN6847 : _GEN6835;
wire  _GEN6849 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN6850 = 1'b1;
wire  _GEN6851 = io_x[6] ? _GEN6850 : _GEN6849;
wire  _GEN6852 = io_x[41] ? _GEN6851 : _GEN6836;
wire  _GEN6853 = io_x[14] ? _GEN6843 : _GEN6852;
wire  _GEN6854 = io_x[0] ? _GEN6845 : _GEN6853;
wire  _GEN6855 = io_x[76] ? _GEN6834 : _GEN6854;
wire  _GEN6856 = 1'b0;
wire  _GEN6857 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN6858 = 1'b0;
wire  _GEN6859 = io_x[0] ? _GEN6858 : _GEN6857;
wire  _GEN6860 = io_x[76] ? _GEN6834 : _GEN6859;
wire  _GEN6861 = io_x[42] ? _GEN6860 : _GEN6855;
wire  _GEN6862 = io_x[38] ? _GEN6861 : _GEN6848;
wire  _GEN6863 = 1'b0;
wire  _GEN6864 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN6865 = io_x[6] ? _GEN6864 : _GEN6850;
wire  _GEN6866 = io_x[41] ? _GEN6865 : _GEN6836;
wire  _GEN6867 = io_x[14] ? _GEN6843 : _GEN6866;
wire  _GEN6868 = io_x[0] ? _GEN6845 : _GEN6867;
wire  _GEN6869 = io_x[76] ? _GEN6834 : _GEN6868;
wire  _GEN6870 = io_x[42] ? _GEN6869 : _GEN6863;
wire  _GEN6871 = 1'b1;
wire  _GEN6872 = io_x[38] ? _GEN6871 : _GEN6870;
wire  _GEN6873 = io_x[10] ? _GEN6872 : _GEN6862;
wire  _GEN6874 = 1'b1;
wire  _GEN6875 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN6876 = io_x[6] ? _GEN6850 : _GEN6875;
wire  _GEN6877 = io_x[41] ? _GEN6876 : _GEN6836;
wire  _GEN6878 = io_x[14] ? _GEN6843 : _GEN6877;
wire  _GEN6879 = io_x[0] ? _GEN6878 : _GEN6845;
wire  _GEN6880 = io_x[76] ? _GEN6833 : _GEN6879;
wire  _GEN6881 = io_x[42] ? _GEN6880 : _GEN6874;
wire  _GEN6882 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN6883 = io_x[76] ? _GEN6882 : _GEN6834;
wire  _GEN6884 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN6885 = io_x[6] ? _GEN6850 : _GEN6884;
wire  _GEN6886 = io_x[41] ? _GEN6885 : _GEN6836;
wire  _GEN6887 = io_x[14] ? _GEN6843 : _GEN6886;
wire  _GEN6888 = io_x[0] ? _GEN6845 : _GEN6887;
wire  _GEN6889 = io_x[76] ? _GEN6888 : _GEN6833;
wire  _GEN6890 = io_x[42] ? _GEN6889 : _GEN6883;
wire  _GEN6891 = io_x[38] ? _GEN6890 : _GEN6881;
wire  _GEN6892 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN6893 = io_x[41] ? _GEN6892 : _GEN6836;
wire  _GEN6894 = io_x[14] ? _GEN6893 : _GEN6843;
wire  _GEN6895 = io_x[0] ? _GEN6894 : _GEN6845;
wire  _GEN6896 = io_x[76] ? _GEN6834 : _GEN6895;
wire  _GEN6897 = io_x[42] ? _GEN6896 : _GEN6874;
wire  _GEN6898 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN6899 = io_x[0] ? _GEN6845 : _GEN6898;
wire  _GEN6900 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN6901 = io_x[76] ? _GEN6900 : _GEN6899;
wire  _GEN6902 = io_x[42] ? _GEN6874 : _GEN6901;
wire  _GEN6903 = io_x[38] ? _GEN6902 : _GEN6897;
wire  _GEN6904 = io_x[10] ? _GEN6903 : _GEN6891;
wire  _GEN6905 = io_x[71] ? _GEN6904 : _GEN6873;
wire  _GEN6906 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN6907 = io_x[6] ? _GEN6850 : _GEN6906;
wire  _GEN6908 = io_x[41] ? _GEN6836 : _GEN6907;
wire  _GEN6909 = io_x[14] ? _GEN6908 : _GEN6856;
wire  _GEN6910 = io_x[0] ? _GEN6909 : _GEN6845;
wire  _GEN6911 = io_x[76] ? _GEN6910 : _GEN6834;
wire  _GEN6912 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN6913 = 1'b0;
wire  _GEN6914 = 1'b1;
wire  _GEN6915 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN6916 = io_x[2] ? _GEN6837 : _GEN6915;
wire  _GEN6917 = io_x[6] ? _GEN6850 : _GEN6916;
wire  _GEN6918 = io_x[41] ? _GEN6917 : _GEN6912;
wire  _GEN6919 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN6920 = io_x[41] ? _GEN6836 : _GEN6919;
wire  _GEN6921 = io_x[14] ? _GEN6920 : _GEN6918;
wire  _GEN6922 = io_x[0] ? _GEN6858 : _GEN6921;
wire  _GEN6923 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN6924 = 1'b0;
wire  _GEN6925 = io_x[41] ? _GEN6924 : _GEN6923;
wire  _GEN6926 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN6927 = io_x[41] ? _GEN6836 : _GEN6926;
wire  _GEN6928 = io_x[14] ? _GEN6927 : _GEN6925;
wire  _GEN6929 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN6930 = io_x[14] ? _GEN6843 : _GEN6929;
wire  _GEN6931 = io_x[0] ? _GEN6930 : _GEN6928;
wire  _GEN6932 = io_x[76] ? _GEN6931 : _GEN6922;
wire  _GEN6933 = io_x[42] ? _GEN6932 : _GEN6911;
wire  _GEN6934 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN6935 = io_x[14] ? _GEN6934 : _GEN6856;
wire  _GEN6936 = io_x[0] ? _GEN6845 : _GEN6935;
wire  _GEN6937 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN6938 = io_x[76] ? _GEN6937 : _GEN6936;
wire  _GEN6939 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN6940 = io_x[2] ? _GEN6837 : _GEN6939;
wire  _GEN6941 = io_x[6] ? _GEN6850 : _GEN6940;
wire  _GEN6942 = io_x[41] ? _GEN6941 : _GEN6836;
wire  _GEN6943 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN6944 = io_x[41] ? _GEN6836 : _GEN6943;
wire  _GEN6945 = io_x[14] ? _GEN6944 : _GEN6942;
wire  _GEN6946 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN6947 = io_x[0] ? _GEN6946 : _GEN6945;
wire  _GEN6948 = io_x[76] ? _GEN6834 : _GEN6947;
wire  _GEN6949 = io_x[42] ? _GEN6948 : _GEN6938;
wire  _GEN6950 = io_x[38] ? _GEN6949 : _GEN6933;
wire  _GEN6951 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN6952 = io_x[0] ? _GEN6845 : _GEN6951;
wire  _GEN6953 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN6954 = io_x[41] ? _GEN6836 : _GEN6953;
wire  _GEN6955 = io_x[14] ? _GEN6954 : _GEN6843;
wire  _GEN6956 = io_x[0] ? _GEN6845 : _GEN6955;
wire  _GEN6957 = io_x[76] ? _GEN6956 : _GEN6952;
wire  _GEN6958 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN6959 = io_x[6] ? _GEN6850 : _GEN6958;
wire  _GEN6960 = io_x[41] ? _GEN6836 : _GEN6959;
wire  _GEN6961 = io_x[14] ? _GEN6960 : _GEN6843;
wire  _GEN6962 = io_x[0] ? _GEN6961 : _GEN6845;
wire  _GEN6963 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN6964 = io_x[14] ? _GEN6856 : _GEN6963;
wire  _GEN6965 = io_x[0] ? _GEN6845 : _GEN6964;
wire  _GEN6966 = io_x[76] ? _GEN6965 : _GEN6962;
wire  _GEN6967 = io_x[42] ? _GEN6966 : _GEN6957;
wire  _GEN6968 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN6969 = io_x[0] ? _GEN6968 : _GEN6845;
wire  _GEN6970 = io_x[76] ? _GEN6833 : _GEN6969;
wire  _GEN6971 = io_x[42] ? _GEN6863 : _GEN6970;
wire  _GEN6972 = io_x[38] ? _GEN6971 : _GEN6967;
wire  _GEN6973 = io_x[10] ? _GEN6972 : _GEN6950;
wire  _GEN6974 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN6975 = io_x[76] ? _GEN6833 : _GEN6974;
wire  _GEN6976 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN6977 = io_x[6] ? _GEN6850 : _GEN6976;
wire  _GEN6978 = io_x[41] ? _GEN6977 : _GEN6836;
wire  _GEN6979 = io_x[14] ? _GEN6843 : _GEN6978;
wire  _GEN6980 = io_x[0] ? _GEN6845 : _GEN6979;
wire  _GEN6981 = io_x[76] ? _GEN6980 : _GEN6833;
wire  _GEN6982 = io_x[42] ? _GEN6981 : _GEN6975;
wire  _GEN6983 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN6984 = io_x[41] ? _GEN6983 : _GEN6836;
wire  _GEN6985 = io_x[14] ? _GEN6843 : _GEN6984;
wire  _GEN6986 = io_x[0] ? _GEN6985 : _GEN6845;
wire  _GEN6987 = io_x[76] ? _GEN6833 : _GEN6986;
wire  _GEN6988 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN6989 = io_x[2] ? _GEN6837 : _GEN6988;
wire  _GEN6990 = io_x[6] ? _GEN6850 : _GEN6989;
wire  _GEN6991 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN6992 = io_x[2] ? _GEN6837 : _GEN6991;
wire  _GEN6993 = io_x[6] ? _GEN6850 : _GEN6992;
wire  _GEN6994 = io_x[41] ? _GEN6993 : _GEN6990;
wire  _GEN6995 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN6996 = io_x[2] ? _GEN6837 : _GEN6995;
wire  _GEN6997 = io_x[6] ? _GEN6840 : _GEN6996;
wire  _GEN6998 = io_x[41] ? _GEN6836 : _GEN6997;
wire  _GEN6999 = io_x[14] ? _GEN6998 : _GEN6994;
wire  _GEN7000 = io_x[0] ? _GEN6845 : _GEN6999;
wire  _GEN7001 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN7002 = io_x[14] ? _GEN6843 : _GEN7001;
wire  _GEN7003 = io_x[0] ? _GEN6845 : _GEN7002;
wire  _GEN7004 = io_x[76] ? _GEN7003 : _GEN7000;
wire  _GEN7005 = io_x[42] ? _GEN7004 : _GEN6987;
wire  _GEN7006 = io_x[38] ? _GEN7005 : _GEN6982;
wire  _GEN7007 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7008 = io_x[0] ? _GEN6858 : _GEN7007;
wire  _GEN7009 = io_x[76] ? _GEN7008 : _GEN6834;
wire  _GEN7010 = io_x[42] ? _GEN7009 : _GEN6874;
wire  _GEN7011 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN7012 = io_x[14] ? _GEN7011 : _GEN6856;
wire  _GEN7013 = io_x[0] ? _GEN7012 : _GEN6858;
wire  _GEN7014 = io_x[76] ? _GEN6834 : _GEN7013;
wire  _GEN7015 = io_x[42] ? _GEN6874 : _GEN7014;
wire  _GEN7016 = io_x[38] ? _GEN7015 : _GEN7010;
wire  _GEN7017 = io_x[10] ? _GEN7016 : _GEN7006;
wire  _GEN7018 = io_x[71] ? _GEN7017 : _GEN6973;
wire  _GEN7019 = io_x[70] ? _GEN7018 : _GEN6905;
wire  _GEN7020 = 1'b0;
wire  _GEN7021 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7022 = io_x[41] ? _GEN7021 : _GEN6836;
wire  _GEN7023 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7024 = io_x[41] ? _GEN7023 : _GEN6836;
wire  _GEN7025 = io_x[14] ? _GEN7024 : _GEN7022;
wire  _GEN7026 = io_x[0] ? _GEN7025 : _GEN6845;
wire  _GEN7027 = io_x[76] ? _GEN7026 : _GEN6833;
wire  _GEN7028 = io_x[42] ? _GEN6874 : _GEN7027;
wire  _GEN7029 = io_x[38] ? _GEN7028 : _GEN6871;
wire  _GEN7030 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7031 = io_x[0] ? _GEN7030 : _GEN6845;
wire  _GEN7032 = io_x[76] ? _GEN7031 : _GEN6833;
wire  _GEN7033 = io_x[42] ? _GEN6874 : _GEN7032;
wire  _GEN7034 = io_x[38] ? _GEN7033 : _GEN6871;
wire  _GEN7035 = io_x[10] ? _GEN7034 : _GEN7029;
wire  _GEN7036 = 1'b0;
wire  _GEN7037 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7038 = io_x[41] ? _GEN6836 : _GEN7037;
wire  _GEN7039 = io_x[14] ? _GEN7038 : _GEN6843;
wire  _GEN7040 = io_x[0] ? _GEN6845 : _GEN7039;
wire  _GEN7041 = io_x[76] ? _GEN6834 : _GEN7040;
wire  _GEN7042 = io_x[42] ? _GEN7041 : _GEN6874;
wire  _GEN7043 = io_x[38] ? _GEN7042 : _GEN7036;
wire  _GEN7044 = 1'b1;
wire  _GEN7045 = io_x[10] ? _GEN7044 : _GEN7043;
wire  _GEN7046 = io_x[71] ? _GEN7045 : _GEN7035;
wire  _GEN7047 = io_x[70] ? _GEN7046 : _GEN7020;
wire  _GEN7048 = io_x[33] ? _GEN7047 : _GEN7019;
wire  _GEN7049 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN7050 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7051 = io_x[6] ? _GEN6850 : _GEN7050;
wire  _GEN7052 = io_x[41] ? _GEN7051 : _GEN6836;
wire  _GEN7053 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN7054 = io_x[2] ? _GEN7053 : _GEN6837;
wire  _GEN7055 = io_x[6] ? _GEN6840 : _GEN7054;
wire  _GEN7056 = io_x[41] ? _GEN7055 : _GEN6836;
wire  _GEN7057 = io_x[14] ? _GEN7056 : _GEN7052;
wire  _GEN7058 = io_x[0] ? _GEN6845 : _GEN7057;
wire  _GEN7059 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7060 = io_x[0] ? _GEN6845 : _GEN7059;
wire  _GEN7061 = io_x[76] ? _GEN7060 : _GEN7058;
wire  _GEN7062 = io_x[42] ? _GEN7061 : _GEN7049;
wire  _GEN7063 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7064 = io_x[41] ? _GEN6836 : _GEN7063;
wire  _GEN7065 = io_x[14] ? _GEN7064 : _GEN6843;
wire  _GEN7066 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN7067 = io_x[14] ? _GEN6843 : _GEN7066;
wire  _GEN7068 = io_x[0] ? _GEN7067 : _GEN7065;
wire  _GEN7069 = io_x[76] ? _GEN6834 : _GEN7068;
wire  _GEN7070 = io_x[42] ? _GEN7069 : _GEN6863;
wire  _GEN7071 = io_x[38] ? _GEN7070 : _GEN7062;
wire  _GEN7072 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7073 = io_x[0] ? _GEN6845 : _GEN7072;
wire  _GEN7074 = io_x[76] ? _GEN7073 : _GEN6833;
wire  _GEN7075 = io_x[42] ? _GEN7074 : _GEN6874;
wire  _GEN7076 = io_x[38] ? _GEN7036 : _GEN7075;
wire  _GEN7077 = io_x[10] ? _GEN7076 : _GEN7071;
wire  _GEN7078 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7079 = io_x[0] ? _GEN6845 : _GEN7078;
wire  _GEN7080 = io_x[76] ? _GEN6834 : _GEN7079;
wire  _GEN7081 = io_x[42] ? _GEN7080 : _GEN6863;
wire  _GEN7082 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7083 = io_x[6] ? _GEN7082 : _GEN6840;
wire  _GEN7084 = io_x[41] ? _GEN6836 : _GEN7083;
wire  _GEN7085 = io_x[14] ? _GEN7084 : _GEN6856;
wire  _GEN7086 = io_x[0] ? _GEN6845 : _GEN7085;
wire  _GEN7087 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7088 = io_x[0] ? _GEN6845 : _GEN7087;
wire  _GEN7089 = io_x[76] ? _GEN7088 : _GEN7086;
wire  _GEN7090 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN7091 = io_x[76] ? _GEN7090 : _GEN6833;
wire  _GEN7092 = io_x[42] ? _GEN7091 : _GEN7089;
wire  _GEN7093 = io_x[38] ? _GEN7092 : _GEN7081;
wire  _GEN7094 = 1'b0;
wire  _GEN7095 = io_x[10] ? _GEN7094 : _GEN7093;
wire  _GEN7096 = io_x[71] ? _GEN7095 : _GEN7077;
wire  _GEN7097 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7098 = io_x[0] ? _GEN6845 : _GEN7097;
wire  _GEN7099 = io_x[76] ? _GEN6833 : _GEN7098;
wire  _GEN7100 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7101 = io_x[41] ? _GEN6924 : _GEN7100;
wire  _GEN7102 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7103 = io_x[41] ? _GEN6836 : _GEN7102;
wire  _GEN7104 = io_x[14] ? _GEN7103 : _GEN7101;
wire  _GEN7105 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7106 = io_x[6] ? _GEN7105 : _GEN6840;
wire  _GEN7107 = io_x[41] ? _GEN6836 : _GEN7106;
wire  _GEN7108 = io_x[14] ? _GEN7107 : _GEN6856;
wire  _GEN7109 = io_x[0] ? _GEN7108 : _GEN7104;
wire  _GEN7110 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN7111 = io_x[2] ? _GEN6837 : _GEN7110;
wire  _GEN7112 = io_x[6] ? _GEN6850 : _GEN7111;
wire  _GEN7113 = io_x[41] ? _GEN7112 : _GEN6924;
wire  _GEN7114 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN7115 = io_x[2] ? _GEN6837 : _GEN7114;
wire  _GEN7116 = io_x[6] ? _GEN6840 : _GEN7115;
wire  _GEN7117 = io_x[41] ? _GEN7116 : _GEN6836;
wire  _GEN7118 = io_x[14] ? _GEN7117 : _GEN7113;
wire  _GEN7119 = io_x[0] ? _GEN6858 : _GEN7118;
wire  _GEN7120 = io_x[76] ? _GEN7119 : _GEN7109;
wire  _GEN7121 = io_x[42] ? _GEN7120 : _GEN7099;
wire  _GEN7122 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7123 = io_x[41] ? _GEN6924 : _GEN7122;
wire  _GEN7124 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7125 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7126 = io_x[6] ? _GEN7125 : _GEN7124;
wire  _GEN7127 = io_x[41] ? _GEN6836 : _GEN7126;
wire  _GEN7128 = io_x[14] ? _GEN7127 : _GEN7123;
wire  _GEN7129 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7130 = io_x[41] ? _GEN6836 : _GEN7129;
wire  _GEN7131 = io_x[14] ? _GEN6856 : _GEN7130;
wire  _GEN7132 = io_x[0] ? _GEN7131 : _GEN7128;
wire  _GEN7133 = io_x[76] ? _GEN6834 : _GEN7132;
wire  _GEN7134 = io_x[42] ? _GEN7133 : _GEN6874;
wire  _GEN7135 = io_x[38] ? _GEN7134 : _GEN7121;
wire  _GEN7136 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7137 = io_x[0] ? _GEN6845 : _GEN7136;
wire  _GEN7138 = io_x[76] ? _GEN6833 : _GEN7137;
wire  _GEN7139 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7140 = io_x[6] ? _GEN7139 : _GEN6850;
wire  _GEN7141 = io_x[41] ? _GEN6836 : _GEN7140;
wire  _GEN7142 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7143 = io_x[41] ? _GEN6836 : _GEN7142;
wire  _GEN7144 = io_x[14] ? _GEN7143 : _GEN7141;
wire  _GEN7145 = io_x[0] ? _GEN7144 : _GEN6845;
wire  _GEN7146 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN7147 = io_x[2] ? _GEN6837 : _GEN7146;
wire  _GEN7148 = io_x[6] ? _GEN6840 : _GEN7147;
wire  _GEN7149 = io_x[41] ? _GEN7148 : _GEN6924;
wire  _GEN7150 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7151 = io_x[41] ? _GEN6836 : _GEN7150;
wire  _GEN7152 = io_x[14] ? _GEN7151 : _GEN7149;
wire  _GEN7153 = io_x[0] ? _GEN6845 : _GEN7152;
wire  _GEN7154 = io_x[76] ? _GEN7153 : _GEN7145;
wire  _GEN7155 = io_x[42] ? _GEN7154 : _GEN7138;
wire  _GEN7156 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7157 = io_x[0] ? _GEN7156 : _GEN6845;
wire  _GEN7158 = io_x[76] ? _GEN6834 : _GEN7157;
wire  _GEN7159 = io_x[42] ? _GEN7158 : _GEN6863;
wire  _GEN7160 = io_x[38] ? _GEN7159 : _GEN7155;
wire  _GEN7161 = io_x[10] ? _GEN7160 : _GEN7135;
wire  _GEN7162 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7163 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7164 = io_x[41] ? _GEN7163 : _GEN7162;
wire  _GEN7165 = io_x[14] ? _GEN7164 : _GEN6843;
wire  _GEN7166 = io_x[0] ? _GEN6858 : _GEN7165;
wire  _GEN7167 = io_x[76] ? _GEN6834 : _GEN7166;
wire  _GEN7168 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7169 = io_x[0] ? _GEN6845 : _GEN7168;
wire  _GEN7170 = io_x[76] ? _GEN7169 : _GEN6833;
wire  _GEN7171 = io_x[42] ? _GEN7170 : _GEN7167;
wire  _GEN7172 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN7173 = io_x[2] ? _GEN6837 : _GEN7172;
wire  _GEN7174 = io_x[6] ? _GEN6850 : _GEN7173;
wire  _GEN7175 = io_x[41] ? _GEN6924 : _GEN7174;
wire  _GEN7176 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7177 = io_x[41] ? _GEN6836 : _GEN7176;
wire  _GEN7178 = io_x[14] ? _GEN7177 : _GEN7175;
wire  _GEN7179 = io_x[0] ? _GEN6845 : _GEN7178;
wire  _GEN7180 = io_x[76] ? _GEN6834 : _GEN7179;
wire  _GEN7181 = io_x[42] ? _GEN7180 : _GEN6863;
wire  _GEN7182 = io_x[38] ? _GEN7181 : _GEN7171;
wire  _GEN7183 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7184 = io_x[0] ? _GEN6845 : _GEN7183;
wire  _GEN7185 = io_x[76] ? _GEN6834 : _GEN7184;
wire  _GEN7186 = io_x[42] ? _GEN6863 : _GEN7185;
wire  _GEN7187 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7188 = io_x[0] ? _GEN6845 : _GEN7187;
wire  _GEN7189 = io_x[76] ? _GEN6834 : _GEN7188;
wire  _GEN7190 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN7191 = io_x[42] ? _GEN7190 : _GEN7189;
wire  _GEN7192 = io_x[38] ? _GEN7191 : _GEN7186;
wire  _GEN7193 = io_x[10] ? _GEN7192 : _GEN7182;
wire  _GEN7194 = io_x[71] ? _GEN7193 : _GEN7161;
wire  _GEN7195 = io_x[70] ? _GEN7194 : _GEN7096;
wire  _GEN7196 = 1'b1;
wire  _GEN7197 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN7198 = io_x[76] ? _GEN6834 : _GEN7197;
wire  _GEN7199 = io_x[42] ? _GEN7198 : _GEN6874;
wire  _GEN7200 = io_x[38] ? _GEN7199 : _GEN6871;
wire  _GEN7201 = io_x[10] ? _GEN7044 : _GEN7200;
wire  _GEN7202 = io_x[71] ? _GEN7201 : _GEN7196;
wire  _GEN7203 = 1'b0;
wire  _GEN7204 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7205 = io_x[41] ? _GEN6836 : _GEN7204;
wire  _GEN7206 = io_x[14] ? _GEN7205 : _GEN6856;
wire  _GEN7207 = io_x[0] ? _GEN6845 : _GEN7206;
wire  _GEN7208 = io_x[76] ? _GEN6834 : _GEN7207;
wire  _GEN7209 = io_x[42] ? _GEN7208 : _GEN6863;
wire  _GEN7210 = io_x[38] ? _GEN7209 : _GEN7036;
wire  _GEN7211 = io_x[10] ? _GEN7094 : _GEN7210;
wire  _GEN7212 = io_x[71] ? _GEN7211 : _GEN7203;
wire  _GEN7213 = io_x[70] ? _GEN7212 : _GEN7202;
wire  _GEN7214 = io_x[33] ? _GEN7213 : _GEN7195;
wire  _GEN7215 = io_x[21] ? _GEN7214 : _GEN7048;
wire  _GEN7216 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7217 = io_x[6] ? _GEN6850 : _GEN7216;
wire  _GEN7218 = io_x[41] ? _GEN7217 : _GEN6836;
wire  _GEN7219 = io_x[14] ? _GEN6843 : _GEN7218;
wire  _GEN7220 = io_x[0] ? _GEN7219 : _GEN6845;
wire  _GEN7221 = io_x[76] ? _GEN6834 : _GEN7220;
wire  _GEN7222 = io_x[42] ? _GEN6874 : _GEN7221;
wire  _GEN7223 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7224 = io_x[6] ? _GEN6850 : _GEN7223;
wire  _GEN7225 = io_x[41] ? _GEN7224 : _GEN6836;
wire  _GEN7226 = io_x[14] ? _GEN6843 : _GEN7225;
wire  _GEN7227 = io_x[0] ? _GEN6845 : _GEN7226;
wire  _GEN7228 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN7229 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7230 = io_x[41] ? _GEN6836 : _GEN7229;
wire  _GEN7231 = io_x[14] ? _GEN7230 : _GEN7228;
wire  _GEN7232 = io_x[0] ? _GEN7231 : _GEN6845;
wire  _GEN7233 = io_x[76] ? _GEN7232 : _GEN7227;
wire  _GEN7234 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7235 = io_x[6] ? _GEN6850 : _GEN7234;
wire  _GEN7236 = io_x[41] ? _GEN6836 : _GEN7235;
wire  _GEN7237 = io_x[14] ? _GEN6856 : _GEN7236;
wire  _GEN7238 = io_x[0] ? _GEN7237 : _GEN6845;
wire  _GEN7239 = io_x[76] ? _GEN6833 : _GEN7238;
wire  _GEN7240 = io_x[42] ? _GEN7239 : _GEN7233;
wire  _GEN7241 = io_x[38] ? _GEN7240 : _GEN7222;
wire  _GEN7242 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7243 = io_x[0] ? _GEN7242 : _GEN6845;
wire  _GEN7244 = io_x[76] ? _GEN6834 : _GEN7243;
wire  _GEN7245 = io_x[42] ? _GEN7244 : _GEN6874;
wire  _GEN7246 = io_x[38] ? _GEN7245 : _GEN6871;
wire  _GEN7247 = io_x[10] ? _GEN7246 : _GEN7241;
wire  _GEN7248 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN7249 = io_x[42] ? _GEN7248 : _GEN6863;
wire  _GEN7250 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7251 = io_x[6] ? _GEN6850 : _GEN7250;
wire  _GEN7252 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN7253 = io_x[2] ? _GEN6837 : _GEN7252;
wire  _GEN7254 = io_x[6] ? _GEN6850 : _GEN7253;
wire  _GEN7255 = io_x[41] ? _GEN7254 : _GEN7251;
wire  _GEN7256 = io_x[14] ? _GEN6843 : _GEN7255;
wire  _GEN7257 = io_x[0] ? _GEN6858 : _GEN7256;
wire  _GEN7258 = io_x[76] ? _GEN7257 : _GEN6833;
wire  _GEN7259 = io_x[42] ? _GEN7258 : _GEN6863;
wire  _GEN7260 = io_x[38] ? _GEN7259 : _GEN7249;
wire  _GEN7261 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7262 = io_x[0] ? _GEN6845 : _GEN7261;
wire  _GEN7263 = io_x[76] ? _GEN6834 : _GEN7262;
wire  _GEN7264 = io_x[42] ? _GEN7263 : _GEN6874;
wire  _GEN7265 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN7266 = io_x[42] ? _GEN6874 : _GEN7265;
wire  _GEN7267 = io_x[38] ? _GEN7266 : _GEN7264;
wire  _GEN7268 = io_x[10] ? _GEN7267 : _GEN7260;
wire  _GEN7269 = io_x[71] ? _GEN7268 : _GEN7247;
wire  _GEN7270 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN7271 = io_x[14] ? _GEN6843 : _GEN7270;
wire  _GEN7272 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN7273 = io_x[14] ? _GEN6856 : _GEN7272;
wire  _GEN7274 = io_x[0] ? _GEN7273 : _GEN7271;
wire  _GEN7275 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7276 = io_x[41] ? _GEN6836 : _GEN7275;
wire  _GEN7277 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7278 = io_x[41] ? _GEN6836 : _GEN7277;
wire  _GEN7279 = io_x[14] ? _GEN7278 : _GEN7276;
wire  _GEN7280 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN7281 = io_x[2] ? _GEN6837 : _GEN7280;
wire  _GEN7282 = io_x[6] ? _GEN6850 : _GEN7281;
wire  _GEN7283 = io_x[41] ? _GEN7282 : _GEN6836;
wire  _GEN7284 = io_x[14] ? _GEN6843 : _GEN7283;
wire  _GEN7285 = io_x[0] ? _GEN7284 : _GEN7279;
wire  _GEN7286 = io_x[76] ? _GEN7285 : _GEN7274;
wire  _GEN7287 = io_x[42] ? _GEN7286 : _GEN6863;
wire  _GEN7288 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7289 = io_x[6] ? _GEN6850 : _GEN7288;
wire  _GEN7290 = io_x[41] ? _GEN7289 : _GEN6836;
wire  _GEN7291 = io_x[14] ? _GEN6843 : _GEN7290;
wire  _GEN7292 = io_x[0] ? _GEN6845 : _GEN7291;
wire  _GEN7293 = io_x[76] ? _GEN6833 : _GEN7292;
wire  _GEN7294 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN7295 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN7296 = io_x[2] ? _GEN6837 : _GEN7295;
wire  _GEN7297 = io_x[6] ? _GEN6850 : _GEN7296;
wire  _GEN7298 = io_x[41] ? _GEN7297 : _GEN6836;
wire  _GEN7299 = io_x[14] ? _GEN6843 : _GEN7298;
wire  _GEN7300 = io_x[0] ? _GEN6858 : _GEN7299;
wire  _GEN7301 = io_x[76] ? _GEN7300 : _GEN7294;
wire  _GEN7302 = io_x[42] ? _GEN7301 : _GEN7293;
wire  _GEN7303 = io_x[38] ? _GEN7302 : _GEN7287;
wire  _GEN7304 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN7305 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7306 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7307 = io_x[6] ? _GEN6850 : _GEN7306;
wire  _GEN7308 = io_x[41] ? _GEN6836 : _GEN7307;
wire  _GEN7309 = io_x[14] ? _GEN7308 : _GEN6856;
wire  _GEN7310 = io_x[0] ? _GEN7309 : _GEN7305;
wire  _GEN7311 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7312 = io_x[0] ? _GEN6845 : _GEN7311;
wire  _GEN7313 = io_x[76] ? _GEN7312 : _GEN7310;
wire  _GEN7314 = io_x[42] ? _GEN7313 : _GEN7304;
wire  _GEN7315 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7316 = io_x[0] ? _GEN6845 : _GEN7315;
wire  _GEN7317 = io_x[76] ? _GEN6833 : _GEN7316;
wire  _GEN7318 = io_x[42] ? _GEN6874 : _GEN7317;
wire  _GEN7319 = io_x[38] ? _GEN7318 : _GEN7314;
wire  _GEN7320 = io_x[10] ? _GEN7319 : _GEN7303;
wire  _GEN7321 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN7322 = io_x[2] ? _GEN6837 : _GEN7321;
wire  _GEN7323 = io_x[6] ? _GEN6850 : _GEN7322;
wire  _GEN7324 = io_x[41] ? _GEN7323 : _GEN6836;
wire  _GEN7325 = io_x[14] ? _GEN6843 : _GEN7324;
wire  _GEN7326 = io_x[0] ? _GEN7325 : _GEN6845;
wire  _GEN7327 = io_x[76] ? _GEN6833 : _GEN7326;
wire  _GEN7328 = io_x[42] ? _GEN7327 : _GEN6874;
wire  _GEN7329 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7330 = io_x[6] ? _GEN6850 : _GEN7329;
wire  _GEN7331 = io_x[41] ? _GEN6836 : _GEN7330;
wire  _GEN7332 = io_x[14] ? _GEN6843 : _GEN7331;
wire  _GEN7333 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7334 = io_x[41] ? _GEN6836 : _GEN7333;
wire  _GEN7335 = io_x[14] ? _GEN7334 : _GEN6856;
wire  _GEN7336 = io_x[0] ? _GEN7335 : _GEN7332;
wire  _GEN7337 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN7338 = io_x[76] ? _GEN7337 : _GEN7336;
wire  _GEN7339 = io_x[42] ? _GEN7338 : _GEN6874;
wire  _GEN7340 = io_x[38] ? _GEN7339 : _GEN7328;
wire  _GEN7341 = io_x[10] ? _GEN7044 : _GEN7340;
wire  _GEN7342 = io_x[71] ? _GEN7341 : _GEN7320;
wire  _GEN7343 = io_x[70] ? _GEN7342 : _GEN7269;
wire  _GEN7344 = io_x[71] ? _GEN7196 : _GEN7203;
wire  _GEN7345 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7346 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7347 = io_x[6] ? _GEN7346 : _GEN7345;
wire  _GEN7348 = io_x[41] ? _GEN7347 : _GEN6836;
wire  _GEN7349 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7350 = io_x[41] ? _GEN7349 : _GEN6836;
wire  _GEN7351 = io_x[14] ? _GEN7350 : _GEN7348;
wire  _GEN7352 = io_x[0] ? _GEN7351 : _GEN6845;
wire  _GEN7353 = io_x[76] ? _GEN7352 : _GEN6834;
wire  _GEN7354 = io_x[42] ? _GEN6874 : _GEN7353;
wire  _GEN7355 = io_x[38] ? _GEN7354 : _GEN6871;
wire  _GEN7356 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7357 = io_x[41] ? _GEN7356 : _GEN6836;
wire  _GEN7358 = io_x[14] ? _GEN7357 : _GEN6856;
wire  _GEN7359 = io_x[0] ? _GEN7358 : _GEN6845;
wire  _GEN7360 = io_x[76] ? _GEN7359 : _GEN6834;
wire  _GEN7361 = io_x[42] ? _GEN6874 : _GEN7360;
wire  _GEN7362 = io_x[38] ? _GEN7361 : _GEN7036;
wire  _GEN7363 = io_x[10] ? _GEN7362 : _GEN7355;
wire  _GEN7364 = io_x[71] ? _GEN7203 : _GEN7363;
wire  _GEN7365 = io_x[70] ? _GEN7364 : _GEN7344;
wire  _GEN7366 = io_x[33] ? _GEN7365 : _GEN7343;
wire  _GEN7367 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN7368 = io_x[76] ? _GEN6834 : _GEN7367;
wire  _GEN7369 = io_x[42] ? _GEN7368 : _GEN6874;
wire  _GEN7370 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7371 = io_x[6] ? _GEN7370 : _GEN6850;
wire  _GEN7372 = io_x[41] ? _GEN6836 : _GEN7371;
wire  _GEN7373 = io_x[14] ? _GEN7372 : _GEN6843;
wire  _GEN7374 = io_x[0] ? _GEN7373 : _GEN6845;
wire  _GEN7375 = io_x[76] ? _GEN7374 : _GEN6834;
wire  _GEN7376 = io_x[42] ? _GEN6863 : _GEN7375;
wire  _GEN7377 = io_x[38] ? _GEN7376 : _GEN7369;
wire  _GEN7378 = io_x[10] ? _GEN7044 : _GEN7377;
wire  _GEN7379 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7380 = io_x[6] ? _GEN6850 : _GEN7379;
wire  _GEN7381 = io_x[41] ? _GEN7380 : _GEN6836;
wire  _GEN7382 = io_x[14] ? _GEN6843 : _GEN7381;
wire  _GEN7383 = io_x[0] ? _GEN7382 : _GEN6845;
wire  _GEN7384 = io_x[76] ? _GEN6834 : _GEN7383;
wire  _GEN7385 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7386 = io_x[6] ? _GEN6850 : _GEN7385;
wire  _GEN7387 = io_x[41] ? _GEN7386 : _GEN6836;
wire  _GEN7388 = io_x[14] ? _GEN6843 : _GEN7387;
wire  _GEN7389 = io_x[0] ? _GEN6858 : _GEN7388;
wire  _GEN7390 = io_x[76] ? _GEN6834 : _GEN7389;
wire  _GEN7391 = io_x[42] ? _GEN7390 : _GEN7384;
wire  _GEN7392 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN7393 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7394 = io_x[6] ? _GEN6850 : _GEN7393;
wire  _GEN7395 = io_x[41] ? _GEN6924 : _GEN7394;
wire  _GEN7396 = io_x[14] ? _GEN6843 : _GEN7395;
wire  _GEN7397 = io_x[0] ? _GEN6845 : _GEN7396;
wire  _GEN7398 = io_x[76] ? _GEN7397 : _GEN6833;
wire  _GEN7399 = io_x[42] ? _GEN7398 : _GEN7392;
wire  _GEN7400 = io_x[38] ? _GEN7399 : _GEN7391;
wire  _GEN7401 = io_x[10] ? _GEN7094 : _GEN7400;
wire  _GEN7402 = io_x[71] ? _GEN7401 : _GEN7378;
wire  _GEN7403 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7404 = io_x[41] ? _GEN6836 : _GEN7403;
wire  _GEN7405 = io_x[14] ? _GEN7404 : _GEN6856;
wire  _GEN7406 = io_x[0] ? _GEN7405 : _GEN6845;
wire  _GEN7407 = io_x[76] ? _GEN6833 : _GEN7406;
wire  _GEN7408 = io_x[42] ? _GEN7407 : _GEN6863;
wire  _GEN7409 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN7410 = io_x[14] ? _GEN6843 : _GEN7409;
wire  _GEN7411 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7412 = io_x[6] ? _GEN7411 : _GEN6850;
wire  _GEN7413 = io_x[41] ? _GEN6836 : _GEN7412;
wire  _GEN7414 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7415 = io_x[6] ? _GEN6850 : _GEN7414;
wire  _GEN7416 = io_x[41] ? _GEN6836 : _GEN7415;
wire  _GEN7417 = io_x[14] ? _GEN7416 : _GEN7413;
wire  _GEN7418 = io_x[0] ? _GEN7417 : _GEN7410;
wire  _GEN7419 = io_x[76] ? _GEN6834 : _GEN7418;
wire  _GEN7420 = io_x[42] ? _GEN7419 : _GEN6874;
wire  _GEN7421 = io_x[38] ? _GEN7420 : _GEN7408;
wire  _GEN7422 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7423 = io_x[41] ? _GEN6836 : _GEN7422;
wire  _GEN7424 = io_x[14] ? _GEN7423 : _GEN6843;
wire  _GEN7425 = io_x[0] ? _GEN6845 : _GEN7424;
wire  _GEN7426 = io_x[76] ? _GEN7425 : _GEN6834;
wire  _GEN7427 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7428 = io_x[41] ? _GEN6836 : _GEN7427;
wire  _GEN7429 = io_x[14] ? _GEN7428 : _GEN6856;
wire  _GEN7430 = io_x[0] ? _GEN7429 : _GEN6845;
wire  _GEN7431 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN7432 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7433 = io_x[41] ? _GEN6836 : _GEN7432;
wire  _GEN7434 = io_x[14] ? _GEN7433 : _GEN7431;
wire  _GEN7435 = io_x[0] ? _GEN6845 : _GEN7434;
wire  _GEN7436 = io_x[76] ? _GEN7435 : _GEN7430;
wire  _GEN7437 = io_x[42] ? _GEN7436 : _GEN7426;
wire  _GEN7438 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7439 = io_x[41] ? _GEN6836 : _GEN7438;
wire  _GEN7440 = io_x[14] ? _GEN6856 : _GEN7439;
wire  _GEN7441 = io_x[0] ? _GEN7440 : _GEN6845;
wire  _GEN7442 = io_x[76] ? _GEN6834 : _GEN7441;
wire  _GEN7443 = io_x[42] ? _GEN7442 : _GEN6863;
wire  _GEN7444 = io_x[38] ? _GEN7443 : _GEN7437;
wire  _GEN7445 = io_x[10] ? _GEN7444 : _GEN7421;
wire  _GEN7446 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN7447 = io_x[42] ? _GEN7446 : _GEN6874;
wire  _GEN7448 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN7449 = io_x[2] ? _GEN6837 : _GEN7448;
wire  _GEN7450 = io_x[6] ? _GEN6850 : _GEN7449;
wire  _GEN7451 = io_x[41] ? _GEN7450 : _GEN6836;
wire  _GEN7452 = io_x[14] ? _GEN6843 : _GEN7451;
wire  _GEN7453 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7454 = io_x[41] ? _GEN6836 : _GEN7453;
wire  _GEN7455 = io_x[14] ? _GEN7454 : _GEN6843;
wire  _GEN7456 = io_x[0] ? _GEN7455 : _GEN7452;
wire  _GEN7457 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN7458 = io_x[14] ? _GEN6843 : _GEN7457;
wire  _GEN7459 = io_x[0] ? _GEN6845 : _GEN7458;
wire  _GEN7460 = io_x[76] ? _GEN7459 : _GEN7456;
wire  _GEN7461 = io_x[42] ? _GEN7460 : _GEN6863;
wire  _GEN7462 = io_x[38] ? _GEN7461 : _GEN7447;
wire  _GEN7463 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN7464 = io_x[76] ? _GEN6834 : _GEN7463;
wire  _GEN7465 = io_x[42] ? _GEN6874 : _GEN7464;
wire  _GEN7466 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN7467 = io_x[38] ? _GEN7466 : _GEN7465;
wire  _GEN7468 = io_x[10] ? _GEN7467 : _GEN7462;
wire  _GEN7469 = io_x[71] ? _GEN7468 : _GEN7445;
wire  _GEN7470 = io_x[70] ? _GEN7469 : _GEN7402;
wire  _GEN7471 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN7472 = io_x[10] ? _GEN7094 : _GEN7471;
wire  _GEN7473 = io_x[71] ? _GEN7472 : _GEN7196;
wire  _GEN7474 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7475 = io_x[0] ? _GEN7474 : _GEN6845;
wire  _GEN7476 = io_x[76] ? _GEN6833 : _GEN7475;
wire  _GEN7477 = io_x[42] ? _GEN7476 : _GEN6874;
wire  _GEN7478 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7479 = io_x[41] ? _GEN7478 : _GEN6836;
wire  _GEN7480 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7481 = io_x[41] ? _GEN7480 : _GEN6924;
wire  _GEN7482 = io_x[14] ? _GEN7481 : _GEN7479;
wire  _GEN7483 = io_x[0] ? _GEN7482 : _GEN6845;
wire  _GEN7484 = io_x[76] ? _GEN6834 : _GEN7483;
wire  _GEN7485 = io_x[42] ? _GEN6874 : _GEN7484;
wire  _GEN7486 = io_x[38] ? _GEN7485 : _GEN7477;
wire  _GEN7487 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7488 = io_x[41] ? _GEN6836 : _GEN7487;
wire  _GEN7489 = io_x[14] ? _GEN7488 : _GEN6843;
wire  _GEN7490 = io_x[0] ? _GEN7489 : _GEN6845;
wire  _GEN7491 = io_x[76] ? _GEN6834 : _GEN7490;
wire  _GEN7492 = io_x[42] ? _GEN7491 : _GEN6874;
wire  _GEN7493 = io_x[38] ? _GEN6871 : _GEN7492;
wire  _GEN7494 = io_x[10] ? _GEN7493 : _GEN7486;
wire  _GEN7495 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7496 = io_x[41] ? _GEN6836 : _GEN7495;
wire  _GEN7497 = io_x[14] ? _GEN6856 : _GEN7496;
wire  _GEN7498 = io_x[0] ? _GEN7497 : _GEN6858;
wire  _GEN7499 = io_x[76] ? _GEN6834 : _GEN7498;
wire  _GEN7500 = io_x[42] ? _GEN7499 : _GEN6863;
wire  _GEN7501 = io_x[38] ? _GEN7500 : _GEN6871;
wire  _GEN7502 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN7503 = io_x[38] ? _GEN7502 : _GEN6871;
wire  _GEN7504 = io_x[10] ? _GEN7503 : _GEN7501;
wire  _GEN7505 = io_x[71] ? _GEN7504 : _GEN7494;
wire  _GEN7506 = io_x[70] ? _GEN7505 : _GEN7473;
wire  _GEN7507 = io_x[33] ? _GEN7506 : _GEN7470;
wire  _GEN7508 = io_x[21] ? _GEN7507 : _GEN7366;
wire  _GEN7509 = io_x[18] ? _GEN7508 : _GEN7215;
wire  _GEN7510 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN7511 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN7512 = io_x[38] ? _GEN7511 : _GEN7510;
wire  _GEN7513 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN7514 = io_x[10] ? _GEN7513 : _GEN7512;
wire  _GEN7515 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN7516 = io_x[76] ? _GEN7515 : _GEN6834;
wire  _GEN7517 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7518 = io_x[0] ? _GEN6845 : _GEN7517;
wire  _GEN7519 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7520 = io_x[0] ? _GEN6845 : _GEN7519;
wire  _GEN7521 = io_x[76] ? _GEN7520 : _GEN7518;
wire  _GEN7522 = io_x[42] ? _GEN7521 : _GEN7516;
wire  _GEN7523 = io_x[38] ? _GEN7522 : _GEN7036;
wire  _GEN7524 = io_x[10] ? _GEN7094 : _GEN7523;
wire  _GEN7525 = io_x[71] ? _GEN7524 : _GEN7514;
wire  _GEN7526 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7527 = io_x[6] ? _GEN7526 : _GEN6840;
wire  _GEN7528 = io_x[41] ? _GEN6836 : _GEN7527;
wire  _GEN7529 = io_x[14] ? _GEN7528 : _GEN6843;
wire  _GEN7530 = io_x[0] ? _GEN6845 : _GEN7529;
wire  _GEN7531 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7532 = io_x[0] ? _GEN6845 : _GEN7531;
wire  _GEN7533 = io_x[76] ? _GEN7532 : _GEN7530;
wire  _GEN7534 = io_x[42] ? _GEN7533 : _GEN6874;
wire  _GEN7535 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7536 = io_x[0] ? _GEN6845 : _GEN7535;
wire  _GEN7537 = io_x[76] ? _GEN6834 : _GEN7536;
wire  _GEN7538 = io_x[42] ? _GEN6874 : _GEN7537;
wire  _GEN7539 = io_x[38] ? _GEN7538 : _GEN7534;
wire  _GEN7540 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7541 = io_x[0] ? _GEN6858 : _GEN7540;
wire  _GEN7542 = io_x[76] ? _GEN6834 : _GEN7541;
wire  _GEN7543 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7544 = io_x[41] ? _GEN6836 : _GEN7543;
wire  _GEN7545 = io_x[14] ? _GEN6843 : _GEN7544;
wire  _GEN7546 = io_x[0] ? _GEN6845 : _GEN7545;
wire  _GEN7547 = io_x[76] ? _GEN7546 : _GEN6834;
wire  _GEN7548 = io_x[42] ? _GEN7547 : _GEN7542;
wire  _GEN7549 = io_x[38] ? _GEN7036 : _GEN7548;
wire  _GEN7550 = io_x[10] ? _GEN7549 : _GEN7539;
wire  _GEN7551 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7552 = io_x[6] ? _GEN6850 : _GEN7551;
wire  _GEN7553 = io_x[41] ? _GEN7552 : _GEN6836;
wire  _GEN7554 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN7555 = io_x[14] ? _GEN7554 : _GEN7553;
wire  _GEN7556 = io_x[0] ? _GEN6845 : _GEN7555;
wire  _GEN7557 = io_x[76] ? _GEN6834 : _GEN7556;
wire  _GEN7558 = io_x[42] ? _GEN6863 : _GEN7557;
wire  _GEN7559 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7560 = io_x[41] ? _GEN6836 : _GEN7559;
wire  _GEN7561 = io_x[14] ? _GEN6856 : _GEN7560;
wire  _GEN7562 = io_x[0] ? _GEN6845 : _GEN7561;
wire  _GEN7563 = io_x[76] ? _GEN6834 : _GEN7562;
wire  _GEN7564 = io_x[42] ? _GEN7563 : _GEN6874;
wire  _GEN7565 = io_x[38] ? _GEN7564 : _GEN7558;
wire  _GEN7566 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7567 = io_x[6] ? _GEN7566 : _GEN6850;
wire  _GEN7568 = io_x[41] ? _GEN7567 : _GEN6836;
wire  _GEN7569 = io_x[14] ? _GEN7568 : _GEN6843;
wire  _GEN7570 = io_x[0] ? _GEN6845 : _GEN7569;
wire  _GEN7571 = io_x[76] ? _GEN6834 : _GEN7570;
wire  _GEN7572 = io_x[42] ? _GEN6874 : _GEN7571;
wire  _GEN7573 = io_x[38] ? _GEN7036 : _GEN7572;
wire  _GEN7574 = io_x[10] ? _GEN7573 : _GEN7565;
wire  _GEN7575 = io_x[71] ? _GEN7574 : _GEN7550;
wire  _GEN7576 = io_x[70] ? _GEN7575 : _GEN7525;
wire  _GEN7577 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7578 = io_x[41] ? _GEN7577 : _GEN6836;
wire  _GEN7579 = io_x[14] ? _GEN6843 : _GEN7578;
wire  _GEN7580 = io_x[0] ? _GEN7579 : _GEN6845;
wire  _GEN7581 = io_x[76] ? _GEN7580 : _GEN6834;
wire  _GEN7582 = io_x[42] ? _GEN6874 : _GEN7581;
wire  _GEN7583 = io_x[38] ? _GEN7582 : _GEN6871;
wire  _GEN7584 = io_x[10] ? _GEN7044 : _GEN7583;
wire  _GEN7585 = io_x[71] ? _GEN7196 : _GEN7584;
wire  _GEN7586 = io_x[70] ? _GEN7585 : _GEN7020;
wire  _GEN7587 = io_x[33] ? _GEN7586 : _GEN7576;
wire  _GEN7588 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7589 = io_x[41] ? _GEN7588 : _GEN6836;
wire  _GEN7590 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7591 = io_x[41] ? _GEN7590 : _GEN6836;
wire  _GEN7592 = io_x[14] ? _GEN7591 : _GEN7589;
wire  _GEN7593 = io_x[0] ? _GEN6858 : _GEN7592;
wire  _GEN7594 = io_x[76] ? _GEN6833 : _GEN7593;
wire  _GEN7595 = io_x[42] ? _GEN7594 : _GEN6874;
wire  _GEN7596 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN7597 = io_x[42] ? _GEN6863 : _GEN7596;
wire  _GEN7598 = io_x[38] ? _GEN7597 : _GEN7595;
wire  _GEN7599 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7600 = io_x[0] ? _GEN7599 : _GEN6845;
wire  _GEN7601 = io_x[76] ? _GEN6834 : _GEN7600;
wire  _GEN7602 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7603 = io_x[41] ? _GEN7602 : _GEN6836;
wire  _GEN7604 = io_x[14] ? _GEN7603 : _GEN6843;
wire  _GEN7605 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7606 = io_x[0] ? _GEN7605 : _GEN7604;
wire  _GEN7607 = io_x[76] ? _GEN6834 : _GEN7606;
wire  _GEN7608 = io_x[42] ? _GEN7607 : _GEN7601;
wire  _GEN7609 = io_x[38] ? _GEN6871 : _GEN7608;
wire  _GEN7610 = io_x[10] ? _GEN7609 : _GEN7598;
wire  _GEN7611 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7612 = io_x[6] ? _GEN7611 : _GEN6850;
wire  _GEN7613 = io_x[41] ? _GEN7612 : _GEN6836;
wire  _GEN7614 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7615 = io_x[6] ? _GEN7614 : _GEN6850;
wire  _GEN7616 = io_x[41] ? _GEN7615 : _GEN6836;
wire  _GEN7617 = io_x[14] ? _GEN7616 : _GEN7613;
wire  _GEN7618 = io_x[0] ? _GEN6845 : _GEN7617;
wire  _GEN7619 = io_x[76] ? _GEN6834 : _GEN7618;
wire  _GEN7620 = io_x[42] ? _GEN7619 : _GEN6874;
wire  _GEN7621 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7622 = io_x[6] ? _GEN6850 : _GEN7621;
wire  _GEN7623 = io_x[41] ? _GEN6836 : _GEN7622;
wire  _GEN7624 = io_x[14] ? _GEN6843 : _GEN7623;
wire  _GEN7625 = io_x[0] ? _GEN6845 : _GEN7624;
wire  _GEN7626 = io_x[76] ? _GEN7625 : _GEN6834;
wire  _GEN7627 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN7628 = io_x[2] ? _GEN6837 : _GEN7627;
wire  _GEN7629 = io_x[6] ? _GEN6850 : _GEN7628;
wire  _GEN7630 = io_x[41] ? _GEN7629 : _GEN6836;
wire  _GEN7631 = io_x[14] ? _GEN6843 : _GEN7630;
wire  _GEN7632 = io_x[0] ? _GEN6845 : _GEN7631;
wire  _GEN7633 = io_x[76] ? _GEN7632 : _GEN6834;
wire  _GEN7634 = io_x[42] ? _GEN7633 : _GEN7626;
wire  _GEN7635 = io_x[38] ? _GEN7634 : _GEN7620;
wire  _GEN7636 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN7637 = io_x[76] ? _GEN6834 : _GEN7636;
wire  _GEN7638 = io_x[42] ? _GEN6863 : _GEN7637;
wire  _GEN7639 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN7640 = io_x[42] ? _GEN6874 : _GEN7639;
wire  _GEN7641 = io_x[38] ? _GEN7640 : _GEN7638;
wire  _GEN7642 = io_x[10] ? _GEN7641 : _GEN7635;
wire  _GEN7643 = io_x[71] ? _GEN7642 : _GEN7610;
wire  _GEN7644 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN7645 = io_x[14] ? _GEN7644 : _GEN6843;
wire  _GEN7646 = io_x[0] ? _GEN6845 : _GEN7645;
wire  _GEN7647 = io_x[76] ? _GEN6833 : _GEN7646;
wire  _GEN7648 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7649 = io_x[6] ? _GEN7648 : _GEN6850;
wire  _GEN7650 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7651 = io_x[6] ? _GEN6850 : _GEN7650;
wire  _GEN7652 = io_x[41] ? _GEN7651 : _GEN7649;
wire  _GEN7653 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7654 = io_x[41] ? _GEN6836 : _GEN7653;
wire  _GEN7655 = io_x[14] ? _GEN7654 : _GEN7652;
wire  _GEN7656 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7657 = io_x[6] ? _GEN7656 : _GEN6850;
wire  _GEN7658 = io_x[41] ? _GEN6836 : _GEN7657;
wire  _GEN7659 = io_x[14] ? _GEN7658 : _GEN6856;
wire  _GEN7660 = io_x[0] ? _GEN7659 : _GEN7655;
wire  _GEN7661 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7662 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7663 = io_x[41] ? _GEN7662 : _GEN7661;
wire  _GEN7664 = io_x[14] ? _GEN6843 : _GEN7663;
wire  _GEN7665 = io_x[0] ? _GEN6845 : _GEN7664;
wire  _GEN7666 = io_x[76] ? _GEN7665 : _GEN7660;
wire  _GEN7667 = io_x[42] ? _GEN7666 : _GEN7647;
wire  _GEN7668 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7669 = io_x[6] ? _GEN7668 : _GEN6850;
wire  _GEN7670 = io_x[41] ? _GEN6836 : _GEN7669;
wire  _GEN7671 = io_x[14] ? _GEN7670 : _GEN6843;
wire  _GEN7672 = io_x[0] ? _GEN6858 : _GEN7671;
wire  _GEN7673 = io_x[76] ? _GEN6833 : _GEN7672;
wire  _GEN7674 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7675 = io_x[0] ? _GEN6858 : _GEN7674;
wire  _GEN7676 = io_x[76] ? _GEN6834 : _GEN7675;
wire  _GEN7677 = io_x[42] ? _GEN7676 : _GEN7673;
wire  _GEN7678 = io_x[38] ? _GEN7677 : _GEN7667;
wire  _GEN7679 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7680 = io_x[41] ? _GEN6836 : _GEN7679;
wire  _GEN7681 = io_x[14] ? _GEN7680 : _GEN6856;
wire  _GEN7682 = io_x[0] ? _GEN7681 : _GEN6858;
wire  _GEN7683 = io_x[76] ? _GEN7682 : _GEN6833;
wire  _GEN7684 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7685 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7686 = io_x[6] ? _GEN7685 : _GEN6850;
wire  _GEN7687 = io_x[41] ? _GEN6836 : _GEN7686;
wire  _GEN7688 = io_x[14] ? _GEN6856 : _GEN7687;
wire  _GEN7689 = io_x[0] ? _GEN7688 : _GEN7684;
wire  _GEN7690 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7691 = io_x[0] ? _GEN6845 : _GEN7690;
wire  _GEN7692 = io_x[76] ? _GEN7691 : _GEN7689;
wire  _GEN7693 = io_x[42] ? _GEN7692 : _GEN7683;
wire  _GEN7694 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7695 = io_x[6] ? _GEN7694 : _GEN6850;
wire  _GEN7696 = io_x[41] ? _GEN7695 : _GEN6836;
wire  _GEN7697 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN7698 = io_x[14] ? _GEN7697 : _GEN7696;
wire  _GEN7699 = io_x[0] ? _GEN6845 : _GEN7698;
wire  _GEN7700 = io_x[76] ? _GEN6834 : _GEN7699;
wire  _GEN7701 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7702 = io_x[6] ? _GEN7701 : _GEN6850;
wire  _GEN7703 = io_x[41] ? _GEN6836 : _GEN7702;
wire  _GEN7704 = io_x[14] ? _GEN6843 : _GEN7703;
wire  _GEN7705 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7706 = io_x[41] ? _GEN6836 : _GEN7705;
wire  _GEN7707 = io_x[14] ? _GEN7706 : _GEN6843;
wire  _GEN7708 = io_x[0] ? _GEN7707 : _GEN7704;
wire  _GEN7709 = io_x[76] ? _GEN6834 : _GEN7708;
wire  _GEN7710 = io_x[42] ? _GEN7709 : _GEN7700;
wire  _GEN7711 = io_x[38] ? _GEN7710 : _GEN7693;
wire  _GEN7712 = io_x[10] ? _GEN7711 : _GEN7678;
wire  _GEN7713 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7714 = io_x[6] ? _GEN6850 : _GEN7713;
wire  _GEN7715 = io_x[41] ? _GEN7714 : _GEN6836;
wire  _GEN7716 = io_x[14] ? _GEN6843 : _GEN7715;
wire  _GEN7717 = io_x[0] ? _GEN6858 : _GEN7716;
wire  _GEN7718 = io_x[76] ? _GEN6834 : _GEN7717;
wire  _GEN7719 = io_x[42] ? _GEN6863 : _GEN7718;
wire  _GEN7720 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7721 = io_x[41] ? _GEN7720 : _GEN6836;
wire  _GEN7722 = io_x[14] ? _GEN7721 : _GEN6856;
wire  _GEN7723 = io_x[0] ? _GEN7722 : _GEN6845;
wire  _GEN7724 = io_x[76] ? _GEN6834 : _GEN7723;
wire  _GEN7725 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7726 = io_x[41] ? _GEN6836 : _GEN7725;
wire  _GEN7727 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7728 = io_x[41] ? _GEN6836 : _GEN7727;
wire  _GEN7729 = io_x[14] ? _GEN7728 : _GEN7726;
wire  _GEN7730 = io_x[0] ? _GEN6845 : _GEN7729;
wire  _GEN7731 = io_x[76] ? _GEN6834 : _GEN7730;
wire  _GEN7732 = io_x[42] ? _GEN7731 : _GEN7724;
wire  _GEN7733 = io_x[38] ? _GEN7732 : _GEN7719;
wire  _GEN7734 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7735 = io_x[41] ? _GEN7734 : _GEN6836;
wire  _GEN7736 = io_x[14] ? _GEN6856 : _GEN7735;
wire  _GEN7737 = io_x[0] ? _GEN7736 : _GEN6845;
wire  _GEN7738 = io_x[76] ? _GEN6834 : _GEN7737;
wire  _GEN7739 = io_x[42] ? _GEN6874 : _GEN7738;
wire  _GEN7740 = io_x[38] ? _GEN7739 : _GEN6871;
wire  _GEN7741 = io_x[10] ? _GEN7740 : _GEN7733;
wire  _GEN7742 = io_x[71] ? _GEN7741 : _GEN7712;
wire  _GEN7743 = io_x[70] ? _GEN7742 : _GEN7643;
wire  _GEN7744 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN7745 = io_x[76] ? _GEN6834 : _GEN7744;
wire  _GEN7746 = io_x[42] ? _GEN7745 : _GEN6874;
wire  _GEN7747 = io_x[38] ? _GEN7746 : _GEN6871;
wire  _GEN7748 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7749 = io_x[0] ? _GEN7748 : _GEN6845;
wire  _GEN7750 = io_x[76] ? _GEN7749 : _GEN6834;
wire  _GEN7751 = io_x[42] ? _GEN6874 : _GEN7750;
wire  _GEN7752 = io_x[38] ? _GEN7751 : _GEN6871;
wire  _GEN7753 = io_x[10] ? _GEN7752 : _GEN7747;
wire  _GEN7754 = io_x[71] ? _GEN7753 : _GEN7196;
wire  _GEN7755 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7756 = io_x[41] ? _GEN6836 : _GEN7755;
wire  _GEN7757 = io_x[14] ? _GEN6843 : _GEN7756;
wire  _GEN7758 = io_x[0] ? _GEN6845 : _GEN7757;
wire  _GEN7759 = io_x[76] ? _GEN6834 : _GEN7758;
wire  _GEN7760 = io_x[42] ? _GEN7759 : _GEN6874;
wire  _GEN7761 = io_x[38] ? _GEN7760 : _GEN6871;
wire  _GEN7762 = io_x[10] ? _GEN7044 : _GEN7761;
wire  _GEN7763 = io_x[71] ? _GEN7762 : _GEN7203;
wire  _GEN7764 = io_x[70] ? _GEN7763 : _GEN7754;
wire  _GEN7765 = io_x[33] ? _GEN7764 : _GEN7743;
wire  _GEN7766 = io_x[21] ? _GEN7765 : _GEN7587;
wire  _GEN7767 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN7768 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7769 = io_x[41] ? _GEN7768 : _GEN6836;
wire  _GEN7770 = io_x[14] ? _GEN6856 : _GEN7769;
wire  _GEN7771 = io_x[0] ? _GEN7770 : _GEN6845;
wire  _GEN7772 = io_x[76] ? _GEN7771 : _GEN6834;
wire  _GEN7773 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7774 = io_x[41] ? _GEN6836 : _GEN7773;
wire  _GEN7775 = io_x[14] ? _GEN7774 : _GEN6843;
wire  _GEN7776 = io_x[0] ? _GEN7775 : _GEN6845;
wire  _GEN7777 = io_x[76] ? _GEN6834 : _GEN7776;
wire  _GEN7778 = io_x[42] ? _GEN7777 : _GEN7772;
wire  _GEN7779 = io_x[38] ? _GEN7778 : _GEN7767;
wire  _GEN7780 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN7781 = io_x[10] ? _GEN7780 : _GEN7779;
wire  _GEN7782 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN7783 = io_x[76] ? _GEN6834 : _GEN7782;
wire  _GEN7784 = io_x[42] ? _GEN7783 : _GEN6874;
wire  _GEN7785 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN7786 = io_x[14] ? _GEN6843 : _GEN7785;
wire  _GEN7787 = io_x[0] ? _GEN7786 : _GEN6845;
wire  _GEN7788 = io_x[76] ? _GEN6834 : _GEN7787;
wire  _GEN7789 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN7790 = io_x[14] ? _GEN6843 : _GEN7789;
wire  _GEN7791 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7792 = io_x[0] ? _GEN7791 : _GEN7790;
wire  _GEN7793 = io_x[76] ? _GEN6834 : _GEN7792;
wire  _GEN7794 = io_x[42] ? _GEN7793 : _GEN7788;
wire  _GEN7795 = io_x[38] ? _GEN7794 : _GEN7784;
wire  _GEN7796 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7797 = io_x[0] ? _GEN7796 : _GEN6858;
wire  _GEN7798 = io_x[76] ? _GEN6834 : _GEN7797;
wire  _GEN7799 = io_x[42] ? _GEN7798 : _GEN6874;
wire  _GEN7800 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN7801 = io_x[2] ? _GEN7800 : _GEN6837;
wire  _GEN7802 = io_x[6] ? _GEN6850 : _GEN7801;
wire  _GEN7803 = io_x[41] ? _GEN6836 : _GEN7802;
wire  _GEN7804 = io_x[14] ? _GEN7803 : _GEN6856;
wire  _GEN7805 = io_x[0] ? _GEN7804 : _GEN6858;
wire  _GEN7806 = io_x[76] ? _GEN6834 : _GEN7805;
wire  _GEN7807 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN7808 = io_x[42] ? _GEN7807 : _GEN7806;
wire  _GEN7809 = io_x[38] ? _GEN7808 : _GEN7799;
wire  _GEN7810 = io_x[10] ? _GEN7809 : _GEN7795;
wire  _GEN7811 = io_x[71] ? _GEN7810 : _GEN7781;
wire  _GEN7812 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7813 = io_x[41] ? _GEN7812 : _GEN6836;
wire  _GEN7814 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7815 = io_x[41] ? _GEN7814 : _GEN6836;
wire  _GEN7816 = io_x[14] ? _GEN7815 : _GEN7813;
wire  _GEN7817 = io_x[0] ? _GEN7816 : _GEN6845;
wire  _GEN7818 = io_x[76] ? _GEN6833 : _GEN7817;
wire  _GEN7819 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7820 = io_x[0] ? _GEN7819 : _GEN6858;
wire  _GEN7821 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7822 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7823 = io_x[41] ? _GEN7822 : _GEN7821;
wire  _GEN7824 = io_x[14] ? _GEN6843 : _GEN7823;
wire  _GEN7825 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7826 = io_x[41] ? _GEN6836 : _GEN7825;
wire  _GEN7827 = io_x[14] ? _GEN6843 : _GEN7826;
wire  _GEN7828 = io_x[0] ? _GEN7827 : _GEN7824;
wire  _GEN7829 = io_x[76] ? _GEN7828 : _GEN7820;
wire  _GEN7830 = io_x[42] ? _GEN7829 : _GEN7818;
wire  _GEN7831 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN7832 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7833 = io_x[41] ? _GEN7832 : _GEN6836;
wire  _GEN7834 = io_x[14] ? _GEN6843 : _GEN7833;
wire  _GEN7835 = io_x[0] ? _GEN7834 : _GEN6845;
wire  _GEN7836 = io_x[76] ? _GEN7835 : _GEN7831;
wire  _GEN7837 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7838 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7839 = io_x[6] ? _GEN7838 : _GEN7837;
wire  _GEN7840 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN7841 = io_x[2] ? _GEN6837 : _GEN7840;
wire  _GEN7842 = io_x[6] ? _GEN6850 : _GEN7841;
wire  _GEN7843 = io_x[41] ? _GEN7842 : _GEN7839;
wire  _GEN7844 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7845 = io_x[6] ? _GEN6840 : _GEN7844;
wire  _GEN7846 = io_x[41] ? _GEN6836 : _GEN7845;
wire  _GEN7847 = io_x[14] ? _GEN7846 : _GEN7843;
wire  _GEN7848 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7849 = io_x[41] ? _GEN6836 : _GEN7848;
wire  _GEN7850 = io_x[14] ? _GEN6843 : _GEN7849;
wire  _GEN7851 = io_x[0] ? _GEN7850 : _GEN7847;
wire  _GEN7852 = io_x[76] ? _GEN6834 : _GEN7851;
wire  _GEN7853 = io_x[42] ? _GEN7852 : _GEN7836;
wire  _GEN7854 = io_x[38] ? _GEN7853 : _GEN7830;
wire  _GEN7855 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7856 = io_x[41] ? _GEN6924 : _GEN7855;
wire  _GEN7857 = io_x[14] ? _GEN6843 : _GEN7856;
wire  _GEN7858 = io_x[0] ? _GEN7857 : _GEN6845;
wire  _GEN7859 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN7860 = io_x[14] ? _GEN6843 : _GEN7859;
wire  _GEN7861 = io_x[0] ? _GEN6845 : _GEN7860;
wire  _GEN7862 = io_x[76] ? _GEN7861 : _GEN7858;
wire  _GEN7863 = io_x[42] ? _GEN7862 : _GEN6863;
wire  _GEN7864 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7865 = io_x[0] ? _GEN6845 : _GEN7864;
wire  _GEN7866 = io_x[76] ? _GEN6834 : _GEN7865;
wire  _GEN7867 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7868 = io_x[6] ? _GEN6840 : _GEN7867;
wire  _GEN7869 = io_x[41] ? _GEN6836 : _GEN7868;
wire  _GEN7870 = io_x[14] ? _GEN7869 : _GEN6843;
wire  _GEN7871 = io_x[0] ? _GEN6845 : _GEN7870;
wire  _GEN7872 = io_x[76] ? _GEN6834 : _GEN7871;
wire  _GEN7873 = io_x[42] ? _GEN7872 : _GEN7866;
wire  _GEN7874 = io_x[38] ? _GEN7873 : _GEN7863;
wire  _GEN7875 = io_x[10] ? _GEN7874 : _GEN7854;
wire  _GEN7876 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN7877 = io_x[14] ? _GEN6843 : _GEN7876;
wire  _GEN7878 = io_x[0] ? _GEN6845 : _GEN7877;
wire  _GEN7879 = io_x[76] ? _GEN6834 : _GEN7878;
wire  _GEN7880 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7881 = io_x[6] ? _GEN6850 : _GEN7880;
wire  _GEN7882 = io_x[41] ? _GEN7881 : _GEN6836;
wire  _GEN7883 = io_x[14] ? _GEN6843 : _GEN7882;
wire  _GEN7884 = io_x[0] ? _GEN6845 : _GEN7883;
wire  _GEN7885 = io_x[76] ? _GEN7884 : _GEN6833;
wire  _GEN7886 = io_x[42] ? _GEN7885 : _GEN7879;
wire  _GEN7887 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN7888 = io_x[6] ? _GEN6850 : _GEN7887;
wire  _GEN7889 = io_x[41] ? _GEN6836 : _GEN7888;
wire  _GEN7890 = io_x[14] ? _GEN6843 : _GEN7889;
wire  _GEN7891 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN7892 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7893 = io_x[41] ? _GEN6836 : _GEN7892;
wire  _GEN7894 = io_x[14] ? _GEN7893 : _GEN7891;
wire  _GEN7895 = io_x[0] ? _GEN7894 : _GEN7890;
wire  _GEN7896 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN7897 = io_x[14] ? _GEN6843 : _GEN7896;
wire  _GEN7898 = io_x[0] ? _GEN6845 : _GEN7897;
wire  _GEN7899 = io_x[76] ? _GEN7898 : _GEN7895;
wire  _GEN7900 = io_x[42] ? _GEN7899 : _GEN6874;
wire  _GEN7901 = io_x[38] ? _GEN7900 : _GEN7886;
wire  _GEN7902 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7903 = io_x[0] ? _GEN6845 : _GEN7902;
wire  _GEN7904 = io_x[76] ? _GEN6834 : _GEN7903;
wire  _GEN7905 = io_x[42] ? _GEN6874 : _GEN7904;
wire  _GEN7906 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7907 = io_x[0] ? _GEN6845 : _GEN7906;
wire  _GEN7908 = io_x[76] ? _GEN6833 : _GEN7907;
wire  _GEN7909 = io_x[42] ? _GEN7908 : _GEN6874;
wire  _GEN7910 = io_x[38] ? _GEN7909 : _GEN7905;
wire  _GEN7911 = io_x[10] ? _GEN7910 : _GEN7901;
wire  _GEN7912 = io_x[71] ? _GEN7911 : _GEN7875;
wire  _GEN7913 = io_x[70] ? _GEN7912 : _GEN7811;
wire  _GEN7914 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7915 = io_x[0] ? _GEN7914 : _GEN6845;
wire  _GEN7916 = io_x[76] ? _GEN7915 : _GEN6834;
wire  _GEN7917 = io_x[42] ? _GEN6874 : _GEN7916;
wire  _GEN7918 = io_x[38] ? _GEN7917 : _GEN6871;
wire  _GEN7919 = io_x[10] ? _GEN7918 : _GEN7044;
wire  _GEN7920 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7921 = io_x[0] ? _GEN7920 : _GEN6845;
wire  _GEN7922 = io_x[76] ? _GEN6834 : _GEN7921;
wire  _GEN7923 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7924 = io_x[0] ? _GEN7923 : _GEN6845;
wire  _GEN7925 = io_x[76] ? _GEN6834 : _GEN7924;
wire  _GEN7926 = io_x[42] ? _GEN7925 : _GEN7922;
wire  _GEN7927 = io_x[38] ? _GEN7926 : _GEN6871;
wire  _GEN7928 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7929 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN7930 = io_x[0] ? _GEN7929 : _GEN7928;
wire  _GEN7931 = io_x[76] ? _GEN6834 : _GEN7930;
wire  _GEN7932 = io_x[42] ? _GEN7931 : _GEN6874;
wire  _GEN7933 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN7934 = io_x[0] ? _GEN7933 : _GEN6845;
wire  _GEN7935 = io_x[76] ? _GEN6834 : _GEN7934;
wire  _GEN7936 = io_x[42] ? _GEN7935 : _GEN6874;
wire  _GEN7937 = io_x[38] ? _GEN7936 : _GEN7932;
wire  _GEN7938 = io_x[10] ? _GEN7937 : _GEN7927;
wire  _GEN7939 = io_x[71] ? _GEN7938 : _GEN7919;
wire  _GEN7940 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN7941 = io_x[76] ? _GEN6834 : _GEN7940;
wire  _GEN7942 = io_x[42] ? _GEN7941 : _GEN6874;
wire  _GEN7943 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7944 = io_x[41] ? _GEN7943 : _GEN6836;
wire  _GEN7945 = io_x[14] ? _GEN6843 : _GEN7944;
wire  _GEN7946 = io_x[0] ? _GEN7945 : _GEN6845;
wire  _GEN7947 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7948 = io_x[41] ? _GEN7947 : _GEN6836;
wire  _GEN7949 = io_x[14] ? _GEN6843 : _GEN7948;
wire  _GEN7950 = io_x[0] ? _GEN7949 : _GEN6845;
wire  _GEN7951 = io_x[76] ? _GEN7950 : _GEN7946;
wire  _GEN7952 = io_x[42] ? _GEN6874 : _GEN7951;
wire  _GEN7953 = io_x[38] ? _GEN7952 : _GEN7942;
wire  _GEN7954 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN7955 = io_x[10] ? _GEN7954 : _GEN7953;
wire  _GEN7956 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN7957 = io_x[71] ? _GEN7956 : _GEN7955;
wire  _GEN7958 = io_x[70] ? _GEN7957 : _GEN7939;
wire  _GEN7959 = io_x[33] ? _GEN7958 : _GEN7913;
wire  _GEN7960 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7961 = io_x[41] ? _GEN7960 : _GEN6836;
wire  _GEN7962 = io_x[14] ? _GEN6843 : _GEN7961;
wire  _GEN7963 = io_x[0] ? _GEN6845 : _GEN7962;
wire  _GEN7964 = io_x[76] ? _GEN6834 : _GEN7963;
wire  _GEN7965 = io_x[42] ? _GEN7964 : _GEN6874;
wire  _GEN7966 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN7967 = io_x[6] ? _GEN6850 : _GEN7966;
wire  _GEN7968 = io_x[41] ? _GEN7967 : _GEN6836;
wire  _GEN7969 = io_x[14] ? _GEN6843 : _GEN7968;
wire  _GEN7970 = io_x[0] ? _GEN6845 : _GEN7969;
wire  _GEN7971 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7972 = io_x[41] ? _GEN6836 : _GEN7971;
wire  _GEN7973 = io_x[14] ? _GEN7972 : _GEN6856;
wire  _GEN7974 = io_x[0] ? _GEN7973 : _GEN6845;
wire  _GEN7975 = io_x[76] ? _GEN7974 : _GEN7970;
wire  _GEN7976 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7977 = io_x[41] ? _GEN6836 : _GEN7976;
wire  _GEN7978 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN7979 = io_x[41] ? _GEN6836 : _GEN7978;
wire  _GEN7980 = io_x[14] ? _GEN7979 : _GEN7977;
wire  _GEN7981 = io_x[0] ? _GEN7980 : _GEN6858;
wire  _GEN7982 = io_x[76] ? _GEN6833 : _GEN7981;
wire  _GEN7983 = io_x[42] ? _GEN7982 : _GEN7975;
wire  _GEN7984 = io_x[38] ? _GEN7983 : _GEN7965;
wire  _GEN7985 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7986 = io_x[41] ? _GEN7985 : _GEN6836;
wire  _GEN7987 = io_x[14] ? _GEN6856 : _GEN7986;
wire  _GEN7988 = io_x[0] ? _GEN7987 : _GEN6845;
wire  _GEN7989 = io_x[76] ? _GEN6834 : _GEN7988;
wire  _GEN7990 = io_x[42] ? _GEN7989 : _GEN6874;
wire  _GEN7991 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7992 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN7993 = io_x[41] ? _GEN7992 : _GEN7991;
wire  _GEN7994 = io_x[14] ? _GEN7993 : _GEN6843;
wire  _GEN7995 = io_x[0] ? _GEN7994 : _GEN6858;
wire  _GEN7996 = io_x[76] ? _GEN6833 : _GEN7995;
wire  _GEN7997 = io_x[42] ? _GEN7996 : _GEN6863;
wire  _GEN7998 = io_x[38] ? _GEN7997 : _GEN7990;
wire  _GEN7999 = io_x[10] ? _GEN7998 : _GEN7984;
wire  _GEN8000 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN8001 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8002 = io_x[41] ? _GEN8001 : _GEN6836;
wire  _GEN8003 = io_x[14] ? _GEN8002 : _GEN6843;
wire  _GEN8004 = io_x[0] ? _GEN8003 : _GEN6845;
wire  _GEN8005 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8006 = io_x[0] ? _GEN6858 : _GEN8005;
wire  _GEN8007 = io_x[76] ? _GEN8006 : _GEN8004;
wire  _GEN8008 = io_x[42] ? _GEN8007 : _GEN8000;
wire  _GEN8009 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8010 = io_x[2] ? _GEN8009 : _GEN6837;
wire  _GEN8011 = io_x[6] ? _GEN6850 : _GEN8010;
wire  _GEN8012 = io_x[41] ? _GEN6836 : _GEN8011;
wire  _GEN8013 = io_x[14] ? _GEN8012 : _GEN6843;
wire  _GEN8014 = io_x[0] ? _GEN8013 : _GEN6845;
wire  _GEN8015 = io_x[76] ? _GEN6834 : _GEN8014;
wire  _GEN8016 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8017 = io_x[41] ? _GEN6924 : _GEN8016;
wire  _GEN8018 = io_x[14] ? _GEN6843 : _GEN8017;
wire  _GEN8019 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8020 = io_x[6] ? _GEN6850 : _GEN8019;
wire  _GEN8021 = io_x[41] ? _GEN6836 : _GEN8020;
wire  _GEN8022 = io_x[14] ? _GEN8021 : _GEN6843;
wire  _GEN8023 = io_x[0] ? _GEN8022 : _GEN8018;
wire  _GEN8024 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8025 = io_x[2] ? _GEN6837 : _GEN8024;
wire  _GEN8026 = io_x[6] ? _GEN6850 : _GEN8025;
wire  _GEN8027 = io_x[41] ? _GEN8026 : _GEN6836;
wire  _GEN8028 = io_x[14] ? _GEN6843 : _GEN8027;
wire  _GEN8029 = io_x[0] ? _GEN6845 : _GEN8028;
wire  _GEN8030 = io_x[76] ? _GEN8029 : _GEN8023;
wire  _GEN8031 = io_x[42] ? _GEN8030 : _GEN8015;
wire  _GEN8032 = io_x[38] ? _GEN8031 : _GEN8008;
wire  _GEN8033 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8034 = io_x[6] ? _GEN8033 : _GEN6850;
wire  _GEN8035 = io_x[41] ? _GEN8034 : _GEN6836;
wire  _GEN8036 = io_x[14] ? _GEN8035 : _GEN6843;
wire  _GEN8037 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8038 = io_x[41] ? _GEN8037 : _GEN6836;
wire  _GEN8039 = io_x[14] ? _GEN8038 : _GEN6856;
wire  _GEN8040 = io_x[0] ? _GEN8039 : _GEN8036;
wire  _GEN8041 = io_x[76] ? _GEN6834 : _GEN8040;
wire  _GEN8042 = io_x[42] ? _GEN8041 : _GEN6863;
wire  _GEN8043 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8044 = io_x[2] ? _GEN6838 : _GEN8043;
wire  _GEN8045 = io_x[6] ? _GEN6840 : _GEN8044;
wire  _GEN8046 = io_x[41] ? _GEN6924 : _GEN8045;
wire  _GEN8047 = io_x[14] ? _GEN8046 : _GEN6843;
wire  _GEN8048 = io_x[0] ? _GEN8047 : _GEN6858;
wire  _GEN8049 = io_x[76] ? _GEN6834 : _GEN8048;
wire  _GEN8050 = io_x[42] ? _GEN6874 : _GEN8049;
wire  _GEN8051 = io_x[38] ? _GEN8050 : _GEN8042;
wire  _GEN8052 = io_x[10] ? _GEN8051 : _GEN8032;
wire  _GEN8053 = io_x[71] ? _GEN8052 : _GEN7999;
wire  _GEN8054 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8055 = io_x[41] ? _GEN8054 : _GEN6836;
wire  _GEN8056 = io_x[14] ? _GEN6843 : _GEN8055;
wire  _GEN8057 = io_x[0] ? _GEN8056 : _GEN6858;
wire  _GEN8058 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8059 = io_x[6] ? _GEN8058 : _GEN6850;
wire  _GEN8060 = io_x[41] ? _GEN6836 : _GEN8059;
wire  _GEN8061 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8062 = io_x[6] ? _GEN8061 : _GEN6850;
wire  _GEN8063 = io_x[41] ? _GEN6836 : _GEN8062;
wire  _GEN8064 = io_x[14] ? _GEN8063 : _GEN8060;
wire  _GEN8065 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8066 = io_x[6] ? _GEN6850 : _GEN8065;
wire  _GEN8067 = io_x[41] ? _GEN6836 : _GEN8066;
wire  _GEN8068 = io_x[14] ? _GEN8067 : _GEN6843;
wire  _GEN8069 = io_x[0] ? _GEN8068 : _GEN8064;
wire  _GEN8070 = io_x[76] ? _GEN8069 : _GEN8057;
wire  _GEN8071 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8072 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8073 = io_x[6] ? _GEN8072 : _GEN6840;
wire  _GEN8074 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8075 = io_x[41] ? _GEN8074 : _GEN8073;
wire  _GEN8076 = io_x[14] ? _GEN8075 : _GEN6856;
wire  _GEN8077 = io_x[0] ? _GEN8076 : _GEN8071;
wire  _GEN8078 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8079 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8080 = io_x[6] ? _GEN6850 : _GEN8079;
wire  _GEN8081 = io_x[41] ? _GEN8080 : _GEN8078;
wire  _GEN8082 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8083 = io_x[41] ? _GEN8082 : _GEN6836;
wire  _GEN8084 = io_x[14] ? _GEN8083 : _GEN8081;
wire  _GEN8085 = io_x[0] ? _GEN6858 : _GEN8084;
wire  _GEN8086 = io_x[76] ? _GEN8085 : _GEN8077;
wire  _GEN8087 = io_x[42] ? _GEN8086 : _GEN8070;
wire  _GEN8088 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8089 = io_x[6] ? _GEN8088 : _GEN6850;
wire  _GEN8090 = io_x[41] ? _GEN6836 : _GEN8089;
wire  _GEN8091 = io_x[14] ? _GEN8090 : _GEN6856;
wire  _GEN8092 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8093 = io_x[41] ? _GEN6836 : _GEN8092;
wire  _GEN8094 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8095 = io_x[41] ? _GEN6836 : _GEN8094;
wire  _GEN8096 = io_x[14] ? _GEN8095 : _GEN8093;
wire  _GEN8097 = io_x[0] ? _GEN8096 : _GEN8091;
wire  _GEN8098 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8099 = io_x[2] ? _GEN6838 : _GEN8098;
wire  _GEN8100 = io_x[6] ? _GEN6850 : _GEN8099;
wire  _GEN8101 = io_x[41] ? _GEN8100 : _GEN6836;
wire  _GEN8102 = io_x[14] ? _GEN6843 : _GEN8101;
wire  _GEN8103 = io_x[0] ? _GEN6845 : _GEN8102;
wire  _GEN8104 = io_x[76] ? _GEN8103 : _GEN8097;
wire  _GEN8105 = io_x[42] ? _GEN8104 : _GEN6874;
wire  _GEN8106 = io_x[38] ? _GEN8105 : _GEN8087;
wire  _GEN8107 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN8108 = io_x[14] ? _GEN8107 : _GEN6843;
wire  _GEN8109 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN8110 = io_x[0] ? _GEN8109 : _GEN8108;
wire  _GEN8111 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8112 = io_x[0] ? _GEN6858 : _GEN8111;
wire  _GEN8113 = io_x[76] ? _GEN8112 : _GEN8110;
wire  _GEN8114 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8115 = io_x[41] ? _GEN6924 : _GEN8114;
wire  _GEN8116 = io_x[14] ? _GEN8115 : _GEN6843;
wire  _GEN8117 = io_x[0] ? _GEN8116 : _GEN6845;
wire  _GEN8118 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8119 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8120 = io_x[41] ? _GEN8119 : _GEN6836;
wire  _GEN8121 = io_x[14] ? _GEN8120 : _GEN6856;
wire  _GEN8122 = io_x[0] ? _GEN8121 : _GEN8118;
wire  _GEN8123 = io_x[76] ? _GEN8122 : _GEN8117;
wire  _GEN8124 = io_x[42] ? _GEN8123 : _GEN8113;
wire  _GEN8125 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8126 = io_x[6] ? _GEN8125 : _GEN6850;
wire  _GEN8127 = io_x[41] ? _GEN6836 : _GEN8126;
wire  _GEN8128 = io_x[14] ? _GEN8127 : _GEN6843;
wire  _GEN8129 = io_x[0] ? _GEN6845 : _GEN8128;
wire  _GEN8130 = io_x[76] ? _GEN6834 : _GEN8129;
wire  _GEN8131 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8132 = io_x[41] ? _GEN6836 : _GEN8131;
wire  _GEN8133 = io_x[14] ? _GEN8132 : _GEN6843;
wire  _GEN8134 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8135 = io_x[41] ? _GEN6836 : _GEN8134;
wire  _GEN8136 = io_x[14] ? _GEN8135 : _GEN6856;
wire  _GEN8137 = io_x[0] ? _GEN8136 : _GEN8133;
wire  _GEN8138 = io_x[76] ? _GEN6834 : _GEN8137;
wire  _GEN8139 = io_x[42] ? _GEN8138 : _GEN8130;
wire  _GEN8140 = io_x[38] ? _GEN8139 : _GEN8124;
wire  _GEN8141 = io_x[10] ? _GEN8140 : _GEN8106;
wire  _GEN8142 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN8143 = io_x[76] ? _GEN6833 : _GEN8142;
wire  _GEN8144 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN8145 = io_x[76] ? _GEN8144 : _GEN6833;
wire  _GEN8146 = io_x[42] ? _GEN8145 : _GEN8143;
wire  _GEN8147 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8148 = io_x[6] ? _GEN8147 : _GEN6850;
wire  _GEN8149 = io_x[41] ? _GEN8148 : _GEN6836;
wire  _GEN8150 = io_x[14] ? _GEN8149 : _GEN6856;
wire  _GEN8151 = io_x[0] ? _GEN8150 : _GEN6845;
wire  _GEN8152 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8153 = io_x[41] ? _GEN6924 : _GEN8152;
wire  _GEN8154 = io_x[14] ? _GEN8153 : _GEN6856;
wire  _GEN8155 = io_x[0] ? _GEN8154 : _GEN6845;
wire  _GEN8156 = io_x[76] ? _GEN8155 : _GEN8151;
wire  _GEN8157 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8158 = io_x[41] ? _GEN6836 : _GEN8157;
wire  _GEN8159 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8160 = io_x[41] ? _GEN6836 : _GEN8159;
wire  _GEN8161 = io_x[14] ? _GEN8160 : _GEN8158;
wire  _GEN8162 = io_x[0] ? _GEN8161 : _GEN6845;
wire  _GEN8163 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN8164 = io_x[14] ? _GEN6856 : _GEN8163;
wire  _GEN8165 = io_x[0] ? _GEN6845 : _GEN8164;
wire  _GEN8166 = io_x[76] ? _GEN8165 : _GEN8162;
wire  _GEN8167 = io_x[42] ? _GEN8166 : _GEN8156;
wire  _GEN8168 = io_x[38] ? _GEN8167 : _GEN8146;
wire  _GEN8169 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN8170 = io_x[14] ? _GEN8169 : _GEN6843;
wire  _GEN8171 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8172 = io_x[6] ? _GEN8171 : _GEN6850;
wire  _GEN8173 = io_x[41] ? _GEN6836 : _GEN8172;
wire  _GEN8174 = io_x[14] ? _GEN8173 : _GEN6856;
wire  _GEN8175 = io_x[0] ? _GEN8174 : _GEN8170;
wire  _GEN8176 = io_x[76] ? _GEN6833 : _GEN8175;
wire  _GEN8177 = io_x[42] ? _GEN6863 : _GEN8176;
wire  _GEN8178 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN8179 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN8180 = io_x[42] ? _GEN8179 : _GEN8178;
wire  _GEN8181 = io_x[38] ? _GEN8180 : _GEN8177;
wire  _GEN8182 = io_x[10] ? _GEN8181 : _GEN8168;
wire  _GEN8183 = io_x[71] ? _GEN8182 : _GEN8141;
wire  _GEN8184 = io_x[70] ? _GEN8183 : _GEN8053;
wire  _GEN8185 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN8186 = io_x[0] ? _GEN8185 : _GEN6845;
wire  _GEN8187 = io_x[76] ? _GEN6834 : _GEN8186;
wire  _GEN8188 = io_x[42] ? _GEN6874 : _GEN8187;
wire  _GEN8189 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN8190 = io_x[38] ? _GEN8189 : _GEN8188;
wire  _GEN8191 = io_x[10] ? _GEN7044 : _GEN8190;
wire  _GEN8192 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN8193 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN8194 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8195 = io_x[6] ? _GEN8194 : _GEN6850;
wire  _GEN8196 = io_x[41] ? _GEN6836 : _GEN8195;
wire  _GEN8197 = io_x[14] ? _GEN8196 : _GEN6843;
wire  _GEN8198 = io_x[0] ? _GEN8197 : _GEN6845;
wire  _GEN8199 = io_x[76] ? _GEN6834 : _GEN8198;
wire  _GEN8200 = io_x[42] ? _GEN8199 : _GEN8193;
wire  _GEN8201 = io_x[38] ? _GEN8200 : _GEN6871;
wire  _GEN8202 = io_x[10] ? _GEN8201 : _GEN8192;
wire  _GEN8203 = io_x[71] ? _GEN8202 : _GEN8191;
wire  _GEN8204 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8205 = io_x[0] ? _GEN6845 : _GEN8204;
wire  _GEN8206 = io_x[76] ? _GEN8205 : _GEN6833;
wire  _GEN8207 = io_x[42] ? _GEN8206 : _GEN6874;
wire  _GEN8208 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8209 = io_x[41] ? _GEN8208 : _GEN6836;
wire  _GEN8210 = io_x[14] ? _GEN6843 : _GEN8209;
wire  _GEN8211 = io_x[0] ? _GEN8210 : _GEN6845;
wire  _GEN8212 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8213 = io_x[6] ? _GEN6840 : _GEN8212;
wire  _GEN8214 = io_x[41] ? _GEN8213 : _GEN6836;
wire  _GEN8215 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8216 = io_x[41] ? _GEN8215 : _GEN6836;
wire  _GEN8217 = io_x[14] ? _GEN8216 : _GEN8214;
wire  _GEN8218 = io_x[0] ? _GEN8217 : _GEN6845;
wire  _GEN8219 = io_x[76] ? _GEN8218 : _GEN8211;
wire  _GEN8220 = io_x[42] ? _GEN6874 : _GEN8219;
wire  _GEN8221 = io_x[38] ? _GEN8220 : _GEN8207;
wire  _GEN8222 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8223 = io_x[41] ? _GEN6836 : _GEN8222;
wire  _GEN8224 = io_x[14] ? _GEN8223 : _GEN6843;
wire  _GEN8225 = io_x[0] ? _GEN8224 : _GEN6845;
wire  _GEN8226 = io_x[76] ? _GEN6834 : _GEN8225;
wire  _GEN8227 = io_x[42] ? _GEN8226 : _GEN6874;
wire  _GEN8228 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8229 = io_x[6] ? _GEN8228 : _GEN6850;
wire  _GEN8230 = io_x[41] ? _GEN8229 : _GEN6836;
wire  _GEN8231 = io_x[14] ? _GEN6856 : _GEN8230;
wire  _GEN8232 = io_x[0] ? _GEN8231 : _GEN6845;
wire  _GEN8233 = io_x[76] ? _GEN8232 : _GEN6834;
wire  _GEN8234 = io_x[42] ? _GEN6874 : _GEN8233;
wire  _GEN8235 = io_x[38] ? _GEN8234 : _GEN8227;
wire  _GEN8236 = io_x[10] ? _GEN8235 : _GEN8221;
wire  _GEN8237 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8238 = io_x[41] ? _GEN6836 : _GEN8237;
wire  _GEN8239 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8240 = io_x[41] ? _GEN6836 : _GEN8239;
wire  _GEN8241 = io_x[14] ? _GEN8240 : _GEN8238;
wire  _GEN8242 = io_x[0] ? _GEN8241 : _GEN6845;
wire  _GEN8243 = io_x[76] ? _GEN6834 : _GEN8242;
wire  _GEN8244 = io_x[42] ? _GEN8243 : _GEN6874;
wire  _GEN8245 = io_x[38] ? _GEN8244 : _GEN6871;
wire  _GEN8246 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8247 = io_x[6] ? _GEN6840 : _GEN8246;
wire  _GEN8248 = io_x[41] ? _GEN6836 : _GEN8247;
wire  _GEN8249 = io_x[14] ? _GEN8248 : _GEN6843;
wire  _GEN8250 = io_x[0] ? _GEN8249 : _GEN6845;
wire  _GEN8251 = io_x[76] ? _GEN6834 : _GEN8250;
wire  _GEN8252 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8253 = io_x[0] ? _GEN8252 : _GEN6845;
wire  _GEN8254 = io_x[76] ? _GEN6834 : _GEN8253;
wire  _GEN8255 = io_x[42] ? _GEN8254 : _GEN8251;
wire  _GEN8256 = io_x[38] ? _GEN8255 : _GEN6871;
wire  _GEN8257 = io_x[10] ? _GEN8256 : _GEN8245;
wire  _GEN8258 = io_x[71] ? _GEN8257 : _GEN8236;
wire  _GEN8259 = io_x[70] ? _GEN8258 : _GEN8203;
wire  _GEN8260 = io_x[33] ? _GEN8259 : _GEN8184;
wire  _GEN8261 = io_x[21] ? _GEN8260 : _GEN7959;
wire  _GEN8262 = io_x[18] ? _GEN8261 : _GEN7766;
wire  _GEN8263 = io_x[20] ? _GEN8262 : _GEN7509;
wire  _GEN8264 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8265 = io_x[6] ? _GEN6850 : _GEN8264;
wire  _GEN8266 = io_x[41] ? _GEN8265 : _GEN6836;
wire  _GEN8267 = io_x[14] ? _GEN6843 : _GEN8266;
wire  _GEN8268 = io_x[0] ? _GEN8267 : _GEN6858;
wire  _GEN8269 = io_x[76] ? _GEN6833 : _GEN8268;
wire  _GEN8270 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8271 = io_x[0] ? _GEN8270 : _GEN6845;
wire  _GEN8272 = io_x[76] ? _GEN6834 : _GEN8271;
wire  _GEN8273 = io_x[42] ? _GEN8272 : _GEN8269;
wire  _GEN8274 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN8275 = io_x[0] ? _GEN6858 : _GEN8274;
wire  _GEN8276 = io_x[76] ? _GEN6834 : _GEN8275;
wire  _GEN8277 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8278 = io_x[6] ? _GEN6850 : _GEN8277;
wire  _GEN8279 = io_x[41] ? _GEN8278 : _GEN6836;
wire  _GEN8280 = io_x[14] ? _GEN6856 : _GEN8279;
wire  _GEN8281 = io_x[0] ? _GEN8280 : _GEN6858;
wire  _GEN8282 = io_x[76] ? _GEN6834 : _GEN8281;
wire  _GEN8283 = io_x[42] ? _GEN8282 : _GEN8276;
wire  _GEN8284 = io_x[38] ? _GEN8283 : _GEN8273;
wire  _GEN8285 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN8286 = io_x[42] ? _GEN6874 : _GEN8285;
wire  _GEN8287 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8288 = io_x[0] ? _GEN6845 : _GEN8287;
wire  _GEN8289 = io_x[76] ? _GEN8288 : _GEN6834;
wire  _GEN8290 = io_x[42] ? _GEN8289 : _GEN6874;
wire  _GEN8291 = io_x[38] ? _GEN8290 : _GEN8286;
wire  _GEN8292 = io_x[10] ? _GEN8291 : _GEN8284;
wire  _GEN8293 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8294 = io_x[6] ? _GEN6850 : _GEN8293;
wire  _GEN8295 = io_x[41] ? _GEN6836 : _GEN8294;
wire  _GEN8296 = io_x[14] ? _GEN6856 : _GEN8295;
wire  _GEN8297 = io_x[0] ? _GEN6845 : _GEN8296;
wire  _GEN8298 = io_x[76] ? _GEN8297 : _GEN6834;
wire  _GEN8299 = io_x[42] ? _GEN8298 : _GEN6874;
wire  _GEN8300 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8301 = io_x[0] ? _GEN8300 : _GEN6858;
wire  _GEN8302 = io_x[76] ? _GEN6833 : _GEN8301;
wire  _GEN8303 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN8304 = io_x[14] ? _GEN6843 : _GEN8303;
wire  _GEN8305 = io_x[0] ? _GEN6845 : _GEN8304;
wire  _GEN8306 = io_x[76] ? _GEN8305 : _GEN6833;
wire  _GEN8307 = io_x[42] ? _GEN8306 : _GEN8302;
wire  _GEN8308 = io_x[38] ? _GEN8307 : _GEN8299;
wire  _GEN8309 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8310 = io_x[6] ? _GEN6850 : _GEN8309;
wire  _GEN8311 = io_x[41] ? _GEN6836 : _GEN8310;
wire  _GEN8312 = io_x[14] ? _GEN6843 : _GEN8311;
wire  _GEN8313 = io_x[0] ? _GEN6845 : _GEN8312;
wire  _GEN8314 = io_x[76] ? _GEN8313 : _GEN6834;
wire  _GEN8315 = io_x[42] ? _GEN8314 : _GEN6874;
wire  _GEN8316 = io_x[38] ? _GEN6871 : _GEN8315;
wire  _GEN8317 = io_x[10] ? _GEN8316 : _GEN8308;
wire  _GEN8318 = io_x[71] ? _GEN8317 : _GEN8292;
wire  _GEN8319 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8320 = io_x[2] ? _GEN6837 : _GEN8319;
wire  _GEN8321 = io_x[6] ? _GEN6850 : _GEN8320;
wire  _GEN8322 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8323 = io_x[6] ? _GEN6850 : _GEN8322;
wire  _GEN8324 = io_x[41] ? _GEN8323 : _GEN8321;
wire  _GEN8325 = io_x[14] ? _GEN6843 : _GEN8324;
wire  _GEN8326 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8327 = io_x[0] ? _GEN8326 : _GEN8325;
wire  _GEN8328 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8329 = io_x[2] ? _GEN6837 : _GEN8328;
wire  _GEN8330 = io_x[6] ? _GEN6850 : _GEN8329;
wire  _GEN8331 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8332 = io_x[2] ? _GEN6837 : _GEN8331;
wire  _GEN8333 = io_x[6] ? _GEN6850 : _GEN8332;
wire  _GEN8334 = io_x[41] ? _GEN8333 : _GEN8330;
wire  _GEN8335 = io_x[14] ? _GEN6843 : _GEN8334;
wire  _GEN8336 = io_x[0] ? _GEN6858 : _GEN8335;
wire  _GEN8337 = io_x[76] ? _GEN8336 : _GEN8327;
wire  _GEN8338 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN8339 = io_x[42] ? _GEN8338 : _GEN8337;
wire  _GEN8340 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN8341 = io_x[0] ? _GEN6845 : _GEN8340;
wire  _GEN8342 = io_x[76] ? _GEN8341 : _GEN6834;
wire  _GEN8343 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8344 = io_x[6] ? _GEN6850 : _GEN8343;
wire  _GEN8345 = io_x[41] ? _GEN6836 : _GEN8344;
wire  _GEN8346 = io_x[14] ? _GEN6843 : _GEN8345;
wire  _GEN8347 = io_x[0] ? _GEN6845 : _GEN8346;
wire  _GEN8348 = io_x[76] ? _GEN8347 : _GEN6834;
wire  _GEN8349 = io_x[42] ? _GEN8348 : _GEN8342;
wire  _GEN8350 = io_x[38] ? _GEN8349 : _GEN8339;
wire  _GEN8351 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN8352 = io_x[42] ? _GEN8351 : _GEN6874;
wire  _GEN8353 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8354 = io_x[6] ? _GEN6850 : _GEN8353;
wire  _GEN8355 = io_x[41] ? _GEN6836 : _GEN8354;
wire  _GEN8356 = io_x[14] ? _GEN6856 : _GEN8355;
wire  _GEN8357 = io_x[0] ? _GEN6845 : _GEN8356;
wire  _GEN8358 = io_x[76] ? _GEN8357 : _GEN6834;
wire  _GEN8359 = io_x[42] ? _GEN8358 : _GEN6874;
wire  _GEN8360 = io_x[38] ? _GEN8359 : _GEN8352;
wire  _GEN8361 = io_x[10] ? _GEN8360 : _GEN8350;
wire  _GEN8362 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8363 = io_x[2] ? _GEN6837 : _GEN8362;
wire  _GEN8364 = io_x[6] ? _GEN6850 : _GEN8363;
wire  _GEN8365 = io_x[41] ? _GEN6836 : _GEN8364;
wire  _GEN8366 = io_x[14] ? _GEN6843 : _GEN8365;
wire  _GEN8367 = io_x[0] ? _GEN8366 : _GEN6845;
wire  _GEN8368 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN8369 = io_x[76] ? _GEN8368 : _GEN8367;
wire  _GEN8370 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8371 = io_x[6] ? _GEN6850 : _GEN8370;
wire  _GEN8372 = io_x[41] ? _GEN6836 : _GEN8371;
wire  _GEN8373 = io_x[14] ? _GEN6843 : _GEN8372;
wire  _GEN8374 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN8375 = io_x[0] ? _GEN8374 : _GEN8373;
wire  _GEN8376 = io_x[76] ? _GEN8375 : _GEN6834;
wire  _GEN8377 = io_x[42] ? _GEN8376 : _GEN8369;
wire  _GEN8378 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN8379 = io_x[76] ? _GEN8378 : _GEN6834;
wire  _GEN8380 = io_x[42] ? _GEN8379 : _GEN6863;
wire  _GEN8381 = io_x[38] ? _GEN8380 : _GEN8377;
wire  _GEN8382 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN8383 = io_x[10] ? _GEN8382 : _GEN8381;
wire  _GEN8384 = io_x[71] ? _GEN8383 : _GEN8361;
wire  _GEN8385 = io_x[70] ? _GEN8384 : _GEN8318;
wire  _GEN8386 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN8387 = io_x[0] ? _GEN6845 : _GEN8386;
wire  _GEN8388 = io_x[76] ? _GEN8387 : _GEN6833;
wire  _GEN8389 = io_x[42] ? _GEN8388 : _GEN6874;
wire  _GEN8390 = io_x[38] ? _GEN7036 : _GEN8389;
wire  _GEN8391 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8392 = io_x[6] ? _GEN6850 : _GEN8391;
wire  _GEN8393 = io_x[41] ? _GEN6836 : _GEN8392;
wire  _GEN8394 = io_x[14] ? _GEN6843 : _GEN8393;
wire  _GEN8395 = io_x[0] ? _GEN6845 : _GEN8394;
wire  _GEN8396 = io_x[76] ? _GEN8395 : _GEN6834;
wire  _GEN8397 = io_x[42] ? _GEN8396 : _GEN6874;
wire  _GEN8398 = io_x[38] ? _GEN6871 : _GEN8397;
wire  _GEN8399 = io_x[10] ? _GEN8398 : _GEN8390;
wire  _GEN8400 = io_x[71] ? _GEN8399 : _GEN7196;
wire  _GEN8401 = io_x[71] ? _GEN7196 : _GEN7203;
wire  _GEN8402 = io_x[70] ? _GEN8401 : _GEN8400;
wire  _GEN8403 = io_x[33] ? _GEN8402 : _GEN8385;
wire  _GEN8404 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN8405 = io_x[38] ? _GEN8404 : _GEN7036;
wire  _GEN8406 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8407 = io_x[0] ? _GEN8406 : _GEN6845;
wire  _GEN8408 = io_x[76] ? _GEN6834 : _GEN8407;
wire  _GEN8409 = io_x[42] ? _GEN8408 : _GEN6874;
wire  _GEN8410 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN8411 = io_x[0] ? _GEN8410 : _GEN6845;
wire  _GEN8412 = io_x[76] ? _GEN6834 : _GEN8411;
wire  _GEN8413 = io_x[42] ? _GEN8412 : _GEN6874;
wire  _GEN8414 = io_x[38] ? _GEN8413 : _GEN8409;
wire  _GEN8415 = io_x[10] ? _GEN8414 : _GEN8405;
wire  _GEN8416 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN8417 = io_x[76] ? _GEN8416 : _GEN6834;
wire  _GEN8418 = io_x[42] ? _GEN8417 : _GEN6863;
wire  _GEN8419 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN8420 = io_x[76] ? _GEN8419 : _GEN6833;
wire  _GEN8421 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN8422 = io_x[14] ? _GEN6843 : _GEN8421;
wire  _GEN8423 = io_x[0] ? _GEN6858 : _GEN8422;
wire  _GEN8424 = io_x[76] ? _GEN8423 : _GEN6834;
wire  _GEN8425 = io_x[42] ? _GEN8424 : _GEN8420;
wire  _GEN8426 = io_x[38] ? _GEN8425 : _GEN8418;
wire  _GEN8427 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN8428 = io_x[76] ? _GEN8427 : _GEN6834;
wire  _GEN8429 = io_x[42] ? _GEN8428 : _GEN6874;
wire  _GEN8430 = io_x[38] ? _GEN8429 : _GEN6871;
wire  _GEN8431 = io_x[10] ? _GEN8430 : _GEN8426;
wire  _GEN8432 = io_x[71] ? _GEN8431 : _GEN8415;
wire  _GEN8433 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8434 = io_x[0] ? _GEN6845 : _GEN8433;
wire  _GEN8435 = io_x[76] ? _GEN6833 : _GEN8434;
wire  _GEN8436 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8437 = io_x[41] ? _GEN6836 : _GEN8436;
wire  _GEN8438 = io_x[14] ? _GEN6843 : _GEN8437;
wire  _GEN8439 = io_x[0] ? _GEN6845 : _GEN8438;
wire  _GEN8440 = io_x[76] ? _GEN6834 : _GEN8439;
wire  _GEN8441 = io_x[42] ? _GEN8440 : _GEN8435;
wire  _GEN8442 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN8443 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN8444 = io_x[0] ? _GEN6845 : _GEN8443;
wire  _GEN8445 = io_x[76] ? _GEN8444 : _GEN6833;
wire  _GEN8446 = io_x[42] ? _GEN8445 : _GEN8442;
wire  _GEN8447 = io_x[38] ? _GEN8446 : _GEN8441;
wire  _GEN8448 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8449 = io_x[41] ? _GEN6836 : _GEN8448;
wire  _GEN8450 = io_x[14] ? _GEN8449 : _GEN6843;
wire  _GEN8451 = io_x[0] ? _GEN8450 : _GEN6858;
wire  _GEN8452 = io_x[76] ? _GEN6834 : _GEN8451;
wire  _GEN8453 = io_x[42] ? _GEN6863 : _GEN8452;
wire  _GEN8454 = io_x[38] ? _GEN7036 : _GEN8453;
wire  _GEN8455 = io_x[10] ? _GEN8454 : _GEN8447;
wire  _GEN8456 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN8457 = io_x[42] ? _GEN6874 : _GEN8456;
wire  _GEN8458 = io_x[38] ? _GEN7036 : _GEN8457;
wire  _GEN8459 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8460 = io_x[0] ? _GEN8459 : _GEN6845;
wire  _GEN8461 = io_x[76] ? _GEN8460 : _GEN6834;
wire  _GEN8462 = io_x[42] ? _GEN8461 : _GEN6874;
wire  _GEN8463 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN8464 = io_x[14] ? _GEN8463 : _GEN6843;
wire  _GEN8465 = io_x[0] ? _GEN8464 : _GEN6845;
wire  _GEN8466 = io_x[76] ? _GEN6833 : _GEN8465;
wire  _GEN8467 = io_x[42] ? _GEN6863 : _GEN8466;
wire  _GEN8468 = io_x[38] ? _GEN8467 : _GEN8462;
wire  _GEN8469 = io_x[10] ? _GEN8468 : _GEN8458;
wire  _GEN8470 = io_x[71] ? _GEN8469 : _GEN8455;
wire  _GEN8471 = io_x[70] ? _GEN8470 : _GEN8432;
wire  _GEN8472 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN8473 = io_x[71] ? _GEN8472 : _GEN7196;
wire  _GEN8474 = 1'b1;
wire  _GEN8475 = io_x[70] ? _GEN8474 : _GEN8473;
wire  _GEN8476 = io_x[33] ? _GEN8475 : _GEN8471;
wire  _GEN8477 = io_x[21] ? _GEN8476 : _GEN8403;
wire  _GEN8478 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8479 = io_x[6] ? _GEN6850 : _GEN8478;
wire  _GEN8480 = io_x[41] ? _GEN6836 : _GEN8479;
wire  _GEN8481 = io_x[14] ? _GEN6843 : _GEN8480;
wire  _GEN8482 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8483 = io_x[41] ? _GEN6924 : _GEN8482;
wire  _GEN8484 = io_x[14] ? _GEN6856 : _GEN8483;
wire  _GEN8485 = io_x[0] ? _GEN8484 : _GEN8481;
wire  _GEN8486 = io_x[76] ? _GEN6834 : _GEN8485;
wire  _GEN8487 = io_x[42] ? _GEN6874 : _GEN8486;
wire  _GEN8488 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN8489 = io_x[76] ? _GEN6834 : _GEN8488;
wire  _GEN8490 = io_x[42] ? _GEN8489 : _GEN6863;
wire  _GEN8491 = io_x[38] ? _GEN8490 : _GEN8487;
wire  _GEN8492 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN8493 = io_x[14] ? _GEN6856 : _GEN8492;
wire  _GEN8494 = io_x[0] ? _GEN6858 : _GEN8493;
wire  _GEN8495 = io_x[76] ? _GEN6834 : _GEN8494;
wire  _GEN8496 = io_x[42] ? _GEN6874 : _GEN8495;
wire  _GEN8497 = io_x[38] ? _GEN6871 : _GEN8496;
wire  _GEN8498 = io_x[10] ? _GEN8497 : _GEN8491;
wire  _GEN8499 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN8500 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN8501 = io_x[2] ? _GEN8500 : _GEN6838;
wire  _GEN8502 = io_x[6] ? _GEN6840 : _GEN8501;
wire  _GEN8503 = io_x[41] ? _GEN8502 : _GEN6836;
wire  _GEN8504 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8505 = io_x[6] ? _GEN6850 : _GEN8504;
wire  _GEN8506 = io_x[41] ? _GEN8505 : _GEN6836;
wire  _GEN8507 = io_x[14] ? _GEN8506 : _GEN8503;
wire  _GEN8508 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8509 = io_x[6] ? _GEN6850 : _GEN8508;
wire  _GEN8510 = io_x[41] ? _GEN8509 : _GEN6836;
wire  _GEN8511 = io_x[14] ? _GEN6843 : _GEN8510;
wire  _GEN8512 = io_x[0] ? _GEN8511 : _GEN8507;
wire  _GEN8513 = io_x[76] ? _GEN8512 : _GEN6834;
wire  _GEN8514 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8515 = io_x[6] ? _GEN6840 : _GEN8514;
wire  _GEN8516 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8517 = io_x[6] ? _GEN6850 : _GEN8516;
wire  _GEN8518 = io_x[41] ? _GEN8517 : _GEN8515;
wire  _GEN8519 = io_x[14] ? _GEN6843 : _GEN8518;
wire  _GEN8520 = io_x[0] ? _GEN6845 : _GEN8519;
wire  _GEN8521 = io_x[76] ? _GEN8520 : _GEN6834;
wire  _GEN8522 = io_x[42] ? _GEN8521 : _GEN8513;
wire  _GEN8523 = io_x[38] ? _GEN8522 : _GEN8499;
wire  _GEN8524 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8525 = io_x[41] ? _GEN8524 : _GEN6836;
wire  _GEN8526 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8527 = io_x[6] ? _GEN6840 : _GEN8526;
wire  _GEN8528 = io_x[41] ? _GEN8527 : _GEN6836;
wire  _GEN8529 = io_x[14] ? _GEN8528 : _GEN8525;
wire  _GEN8530 = io_x[0] ? _GEN6845 : _GEN8529;
wire  _GEN8531 = io_x[76] ? _GEN8530 : _GEN6834;
wire  _GEN8532 = io_x[42] ? _GEN6863 : _GEN8531;
wire  _GEN8533 = io_x[38] ? _GEN8532 : _GEN7036;
wire  _GEN8534 = io_x[10] ? _GEN8533 : _GEN8523;
wire  _GEN8535 = io_x[71] ? _GEN8534 : _GEN8498;
wire  _GEN8536 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8537 = io_x[2] ? _GEN6837 : _GEN8536;
wire  _GEN8538 = io_x[6] ? _GEN6840 : _GEN8537;
wire  _GEN8539 = io_x[41] ? _GEN6924 : _GEN8538;
wire  _GEN8540 = io_x[14] ? _GEN6843 : _GEN8539;
wire  _GEN8541 = io_x[0] ? _GEN8540 : _GEN6845;
wire  _GEN8542 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8543 = io_x[2] ? _GEN6837 : _GEN8542;
wire  _GEN8544 = io_x[6] ? _GEN6850 : _GEN8543;
wire  _GEN8545 = io_x[41] ? _GEN6924 : _GEN8544;
wire  _GEN8546 = io_x[14] ? _GEN6843 : _GEN8545;
wire  _GEN8547 = io_x[0] ? _GEN6845 : _GEN8546;
wire  _GEN8548 = io_x[76] ? _GEN8547 : _GEN8541;
wire  _GEN8549 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN8550 = io_x[14] ? _GEN6843 : _GEN8549;
wire  _GEN8551 = io_x[0] ? _GEN8550 : _GEN6845;
wire  _GEN8552 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8553 = io_x[2] ? _GEN6837 : _GEN8552;
wire  _GEN8554 = io_x[6] ? _GEN6850 : _GEN8553;
wire  _GEN8555 = io_x[41] ? _GEN8554 : _GEN6836;
wire  _GEN8556 = io_x[14] ? _GEN6843 : _GEN8555;
wire  _GEN8557 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN8558 = io_x[14] ? _GEN6843 : _GEN8557;
wire  _GEN8559 = io_x[0] ? _GEN8558 : _GEN8556;
wire  _GEN8560 = io_x[76] ? _GEN8559 : _GEN8551;
wire  _GEN8561 = io_x[42] ? _GEN8560 : _GEN8548;
wire  _GEN8562 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8563 = io_x[6] ? _GEN6850 : _GEN8562;
wire  _GEN8564 = io_x[41] ? _GEN8563 : _GEN6836;
wire  _GEN8565 = io_x[14] ? _GEN6856 : _GEN8564;
wire  _GEN8566 = io_x[0] ? _GEN6858 : _GEN8565;
wire  _GEN8567 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8568 = io_x[6] ? _GEN6850 : _GEN8567;
wire  _GEN8569 = io_x[41] ? _GEN8568 : _GEN6836;
wire  _GEN8570 = io_x[14] ? _GEN6843 : _GEN8569;
wire  _GEN8571 = io_x[0] ? _GEN8570 : _GEN6845;
wire  _GEN8572 = io_x[76] ? _GEN8571 : _GEN8566;
wire  _GEN8573 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8574 = io_x[41] ? _GEN6924 : _GEN8573;
wire  _GEN8575 = io_x[14] ? _GEN6843 : _GEN8574;
wire  _GEN8576 = io_x[0] ? _GEN6845 : _GEN8575;
wire  _GEN8577 = io_x[76] ? _GEN8576 : _GEN6834;
wire  _GEN8578 = io_x[42] ? _GEN8577 : _GEN8572;
wire  _GEN8579 = io_x[38] ? _GEN8578 : _GEN8561;
wire  _GEN8580 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8581 = io_x[41] ? _GEN8580 : _GEN6836;
wire  _GEN8582 = io_x[14] ? _GEN6843 : _GEN8581;
wire  _GEN8583 = io_x[0] ? _GEN8582 : _GEN6845;
wire  _GEN8584 = io_x[76] ? _GEN8583 : _GEN6834;
wire  _GEN8585 = io_x[42] ? _GEN6874 : _GEN8584;
wire  _GEN8586 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN8587 = io_x[38] ? _GEN8586 : _GEN8585;
wire  _GEN8588 = io_x[10] ? _GEN8587 : _GEN8579;
wire  _GEN8589 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN8590 = io_x[76] ? _GEN8589 : _GEN6834;
wire  _GEN8591 = io_x[42] ? _GEN6874 : _GEN8590;
wire  _GEN8592 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN8593 = io_x[0] ? _GEN6845 : _GEN8592;
wire  _GEN8594 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN8595 = io_x[76] ? _GEN8594 : _GEN8593;
wire  _GEN8596 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8597 = io_x[41] ? _GEN6836 : _GEN8596;
wire  _GEN8598 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8599 = io_x[41] ? _GEN6836 : _GEN8598;
wire  _GEN8600 = io_x[14] ? _GEN8599 : _GEN8597;
wire  _GEN8601 = io_x[0] ? _GEN6845 : _GEN8600;
wire  _GEN8602 = io_x[76] ? _GEN8601 : _GEN6834;
wire  _GEN8603 = io_x[42] ? _GEN8602 : _GEN8595;
wire  _GEN8604 = io_x[38] ? _GEN8603 : _GEN8591;
wire  _GEN8605 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8606 = io_x[41] ? _GEN8605 : _GEN6836;
wire  _GEN8607 = io_x[14] ? _GEN6843 : _GEN8606;
wire  _GEN8608 = io_x[0] ? _GEN6845 : _GEN8607;
wire  _GEN8609 = io_x[76] ? _GEN6834 : _GEN8608;
wire  _GEN8610 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8611 = io_x[41] ? _GEN6836 : _GEN8610;
wire  _GEN8612 = io_x[14] ? _GEN8611 : _GEN6843;
wire  _GEN8613 = io_x[0] ? _GEN6845 : _GEN8612;
wire  _GEN8614 = io_x[76] ? _GEN8613 : _GEN6834;
wire  _GEN8615 = io_x[42] ? _GEN8614 : _GEN8609;
wire  _GEN8616 = io_x[38] ? _GEN8615 : _GEN6871;
wire  _GEN8617 = io_x[10] ? _GEN8616 : _GEN8604;
wire  _GEN8618 = io_x[71] ? _GEN8617 : _GEN8588;
wire  _GEN8619 = io_x[70] ? _GEN8618 : _GEN8535;
wire  _GEN8620 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN8621 = io_x[38] ? _GEN7036 : _GEN8620;
wire  _GEN8622 = io_x[10] ? _GEN7044 : _GEN8621;
wire  _GEN8623 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8624 = io_x[41] ? _GEN6836 : _GEN8623;
wire  _GEN8625 = io_x[14] ? _GEN6843 : _GEN8624;
wire  _GEN8626 = io_x[0] ? _GEN6845 : _GEN8625;
wire  _GEN8627 = io_x[76] ? _GEN8626 : _GEN6834;
wire  _GEN8628 = io_x[42] ? _GEN8627 : _GEN6874;
wire  _GEN8629 = io_x[38] ? _GEN8628 : _GEN6871;
wire  _GEN8630 = io_x[10] ? _GEN7094 : _GEN8629;
wire  _GEN8631 = io_x[71] ? _GEN8630 : _GEN8622;
wire  _GEN8632 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN8633 = io_x[42] ? _GEN6863 : _GEN8632;
wire  _GEN8634 = io_x[38] ? _GEN7036 : _GEN8633;
wire  _GEN8635 = io_x[10] ? _GEN7044 : _GEN8634;
wire  _GEN8636 = io_x[71] ? _GEN8635 : _GEN7196;
wire  _GEN8637 = io_x[70] ? _GEN8636 : _GEN8631;
wire  _GEN8638 = io_x[33] ? _GEN8637 : _GEN8619;
wire  _GEN8639 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8640 = io_x[41] ? _GEN8639 : _GEN6836;
wire  _GEN8641 = io_x[14] ? _GEN6843 : _GEN8640;
wire  _GEN8642 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8643 = io_x[6] ? _GEN6850 : _GEN8642;
wire  _GEN8644 = io_x[41] ? _GEN6836 : _GEN8643;
wire  _GEN8645 = io_x[14] ? _GEN6843 : _GEN8644;
wire  _GEN8646 = io_x[0] ? _GEN8645 : _GEN8641;
wire  _GEN8647 = io_x[76] ? _GEN6833 : _GEN8646;
wire  _GEN8648 = io_x[42] ? _GEN6874 : _GEN8647;
wire  _GEN8649 = io_x[38] ? _GEN7036 : _GEN8648;
wire  _GEN8650 = io_x[10] ? _GEN7094 : _GEN8649;
wire  _GEN8651 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN8652 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8653 = io_x[41] ? _GEN6836 : _GEN8652;
wire  _GEN8654 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8655 = io_x[6] ? _GEN8654 : _GEN6840;
wire  _GEN8656 = io_x[41] ? _GEN6836 : _GEN8655;
wire  _GEN8657 = io_x[14] ? _GEN8656 : _GEN8653;
wire  _GEN8658 = io_x[0] ? _GEN6845 : _GEN8657;
wire  _GEN8659 = io_x[76] ? _GEN8658 : _GEN6834;
wire  _GEN8660 = io_x[42] ? _GEN8659 : _GEN6874;
wire  _GEN8661 = io_x[38] ? _GEN8660 : _GEN8651;
wire  _GEN8662 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8663 = io_x[6] ? _GEN8662 : _GEN6850;
wire  _GEN8664 = io_x[41] ? _GEN8663 : _GEN6836;
wire  _GEN8665 = io_x[14] ? _GEN8664 : _GEN6843;
wire  _GEN8666 = io_x[0] ? _GEN6845 : _GEN8665;
wire  _GEN8667 = io_x[76] ? _GEN8666 : _GEN6834;
wire  _GEN8668 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8669 = io_x[41] ? _GEN6836 : _GEN8668;
wire  _GEN8670 = io_x[14] ? _GEN8669 : _GEN6856;
wire  _GEN8671 = io_x[0] ? _GEN6845 : _GEN8670;
wire  _GEN8672 = io_x[76] ? _GEN8671 : _GEN6834;
wire  _GEN8673 = io_x[42] ? _GEN8672 : _GEN8667;
wire  _GEN8674 = io_x[38] ? _GEN8673 : _GEN6871;
wire  _GEN8675 = io_x[10] ? _GEN8674 : _GEN8661;
wire  _GEN8676 = io_x[71] ? _GEN8675 : _GEN8650;
wire  _GEN8677 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN8678 = io_x[76] ? _GEN8677 : _GEN6833;
wire  _GEN8679 = io_x[42] ? _GEN6863 : _GEN8678;
wire  _GEN8680 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8681 = io_x[41] ? _GEN6836 : _GEN8680;
wire  _GEN8682 = io_x[14] ? _GEN6843 : _GEN8681;
wire  _GEN8683 = io_x[0] ? _GEN6845 : _GEN8682;
wire  _GEN8684 = io_x[76] ? _GEN8683 : _GEN6834;
wire  _GEN8685 = io_x[42] ? _GEN8684 : _GEN6874;
wire  _GEN8686 = io_x[38] ? _GEN8685 : _GEN8679;
wire  _GEN8687 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN8688 = io_x[42] ? _GEN6863 : _GEN8687;
wire  _GEN8689 = io_x[38] ? _GEN8688 : _GEN6871;
wire  _GEN8690 = io_x[10] ? _GEN8689 : _GEN8686;
wire  _GEN8691 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8692 = io_x[41] ? _GEN8691 : _GEN6836;
wire  _GEN8693 = io_x[14] ? _GEN6843 : _GEN8692;
wire  _GEN8694 = io_x[0] ? _GEN6845 : _GEN8693;
wire  _GEN8695 = io_x[76] ? _GEN6833 : _GEN8694;
wire  _GEN8696 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8697 = io_x[41] ? _GEN6836 : _GEN8696;
wire  _GEN8698 = io_x[14] ? _GEN8697 : _GEN6856;
wire  _GEN8699 = io_x[0] ? _GEN6845 : _GEN8698;
wire  _GEN8700 = io_x[76] ? _GEN8699 : _GEN6834;
wire  _GEN8701 = io_x[42] ? _GEN8700 : _GEN8695;
wire  _GEN8702 = io_x[38] ? _GEN8701 : _GEN6871;
wire  _GEN8703 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8704 = io_x[41] ? _GEN6836 : _GEN8703;
wire  _GEN8705 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8706 = io_x[41] ? _GEN6836 : _GEN8705;
wire  _GEN8707 = io_x[14] ? _GEN8706 : _GEN8704;
wire  _GEN8708 = io_x[0] ? _GEN6845 : _GEN8707;
wire  _GEN8709 = io_x[76] ? _GEN8708 : _GEN6833;
wire  _GEN8710 = io_x[42] ? _GEN8709 : _GEN6863;
wire  _GEN8711 = io_x[38] ? _GEN8710 : _GEN6871;
wire  _GEN8712 = io_x[10] ? _GEN8711 : _GEN8702;
wire  _GEN8713 = io_x[71] ? _GEN8712 : _GEN8690;
wire  _GEN8714 = io_x[70] ? _GEN8713 : _GEN8676;
wire  _GEN8715 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8716 = io_x[41] ? _GEN6836 : _GEN8715;
wire  _GEN8717 = io_x[14] ? _GEN6843 : _GEN8716;
wire  _GEN8718 = io_x[0] ? _GEN6845 : _GEN8717;
wire  _GEN8719 = io_x[76] ? _GEN8718 : _GEN6834;
wire  _GEN8720 = io_x[42] ? _GEN8719 : _GEN6874;
wire  _GEN8721 = io_x[38] ? _GEN8720 : _GEN6871;
wire  _GEN8722 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN8723 = io_x[10] ? _GEN8722 : _GEN8721;
wire  _GEN8724 = io_x[71] ? _GEN8723 : _GEN7203;
wire  _GEN8725 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN8726 = io_x[10] ? _GEN7044 : _GEN8725;
wire  _GEN8727 = io_x[71] ? _GEN8726 : _GEN7196;
wire  _GEN8728 = io_x[70] ? _GEN8727 : _GEN8724;
wire  _GEN8729 = io_x[33] ? _GEN8728 : _GEN8714;
wire  _GEN8730 = io_x[21] ? _GEN8729 : _GEN8638;
wire  _GEN8731 = io_x[18] ? _GEN8730 : _GEN8477;
wire  _GEN8732 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8733 = io_x[6] ? _GEN6850 : _GEN8732;
wire  _GEN8734 = io_x[41] ? _GEN6836 : _GEN8733;
wire  _GEN8735 = io_x[14] ? _GEN6856 : _GEN8734;
wire  _GEN8736 = io_x[0] ? _GEN8735 : _GEN6858;
wire  _GEN8737 = io_x[76] ? _GEN6833 : _GEN8736;
wire  _GEN8738 = io_x[42] ? _GEN6874 : _GEN8737;
wire  _GEN8739 = io_x[38] ? _GEN6871 : _GEN8738;
wire  _GEN8740 = io_x[10] ? _GEN7044 : _GEN8739;
wire  _GEN8741 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN8742 = io_x[42] ? _GEN8741 : _GEN6874;
wire  _GEN8743 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN8744 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8745 = io_x[41] ? _GEN8744 : _GEN6836;
wire  _GEN8746 = io_x[14] ? _GEN8745 : _GEN6856;
wire  _GEN8747 = io_x[0] ? _GEN8746 : _GEN6858;
wire  _GEN8748 = io_x[76] ? _GEN8747 : _GEN8743;
wire  _GEN8749 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8750 = io_x[41] ? _GEN6836 : _GEN8749;
wire  _GEN8751 = io_x[14] ? _GEN6843 : _GEN8750;
wire  _GEN8752 = io_x[0] ? _GEN6858 : _GEN8751;
wire  _GEN8753 = io_x[76] ? _GEN8752 : _GEN6834;
wire  _GEN8754 = io_x[42] ? _GEN8753 : _GEN8748;
wire  _GEN8755 = io_x[38] ? _GEN8754 : _GEN8742;
wire  _GEN8756 = io_x[10] ? _GEN7044 : _GEN8755;
wire  _GEN8757 = io_x[71] ? _GEN8756 : _GEN8740;
wire  _GEN8758 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN8759 = io_x[42] ? _GEN8758 : _GEN6863;
wire  _GEN8760 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8761 = io_x[0] ? _GEN6845 : _GEN8760;
wire  _GEN8762 = io_x[76] ? _GEN8761 : _GEN6834;
wire  _GEN8763 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8764 = io_x[41] ? _GEN6836 : _GEN8763;
wire  _GEN8765 = io_x[14] ? _GEN6843 : _GEN8764;
wire  _GEN8766 = io_x[0] ? _GEN6845 : _GEN8765;
wire  _GEN8767 = io_x[76] ? _GEN8766 : _GEN6834;
wire  _GEN8768 = io_x[42] ? _GEN8767 : _GEN8762;
wire  _GEN8769 = io_x[38] ? _GEN8768 : _GEN8759;
wire  _GEN8770 = io_x[10] ? _GEN7044 : _GEN8769;
wire  _GEN8771 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8772 = io_x[2] ? _GEN6837 : _GEN8771;
wire  _GEN8773 = io_x[6] ? _GEN6850 : _GEN8772;
wire  _GEN8774 = io_x[41] ? _GEN6836 : _GEN8773;
wire  _GEN8775 = io_x[14] ? _GEN6843 : _GEN8774;
wire  _GEN8776 = io_x[0] ? _GEN6845 : _GEN8775;
wire  _GEN8777 = io_x[76] ? _GEN8776 : _GEN6834;
wire  _GEN8778 = io_x[42] ? _GEN6874 : _GEN8777;
wire  _GEN8779 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN8780 = io_x[14] ? _GEN6843 : _GEN8779;
wire  _GEN8781 = io_x[0] ? _GEN6845 : _GEN8780;
wire  _GEN8782 = io_x[76] ? _GEN8781 : _GEN6834;
wire  _GEN8783 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN8784 = io_x[0] ? _GEN6845 : _GEN8783;
wire  _GEN8785 = io_x[76] ? _GEN8784 : _GEN6834;
wire  _GEN8786 = io_x[42] ? _GEN8785 : _GEN8782;
wire  _GEN8787 = io_x[38] ? _GEN8786 : _GEN8778;
wire  _GEN8788 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8789 = io_x[41] ? _GEN6836 : _GEN8788;
wire  _GEN8790 = io_x[14] ? _GEN6843 : _GEN8789;
wire  _GEN8791 = io_x[0] ? _GEN6845 : _GEN8790;
wire  _GEN8792 = io_x[76] ? _GEN8791 : _GEN6834;
wire  _GEN8793 = io_x[42] ? _GEN8792 : _GEN6874;
wire  _GEN8794 = io_x[38] ? _GEN8793 : _GEN7036;
wire  _GEN8795 = io_x[10] ? _GEN8794 : _GEN8787;
wire  _GEN8796 = io_x[71] ? _GEN8795 : _GEN8770;
wire  _GEN8797 = io_x[70] ? _GEN8796 : _GEN8757;
wire  _GEN8798 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8799 = io_x[41] ? _GEN6836 : _GEN8798;
wire  _GEN8800 = io_x[14] ? _GEN6843 : _GEN8799;
wire  _GEN8801 = io_x[0] ? _GEN6845 : _GEN8800;
wire  _GEN8802 = io_x[76] ? _GEN8801 : _GEN6834;
wire  _GEN8803 = io_x[42] ? _GEN8802 : _GEN6874;
wire  _GEN8804 = io_x[38] ? _GEN8803 : _GEN6871;
wire  _GEN8805 = io_x[10] ? _GEN7044 : _GEN8804;
wire  _GEN8806 = io_x[71] ? _GEN8805 : _GEN7196;
wire  _GEN8807 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN8808 = io_x[38] ? _GEN6871 : _GEN8807;
wire  _GEN8809 = io_x[10] ? _GEN7044 : _GEN8808;
wire  _GEN8810 = io_x[71] ? _GEN8809 : _GEN7196;
wire  _GEN8811 = io_x[70] ? _GEN8810 : _GEN8806;
wire  _GEN8812 = io_x[33] ? _GEN8811 : _GEN8797;
wire  _GEN8813 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN8814 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN8815 = io_x[76] ? _GEN6834 : _GEN8814;
wire  _GEN8816 = io_x[42] ? _GEN6874 : _GEN8815;
wire  _GEN8817 = io_x[38] ? _GEN6871 : _GEN8816;
wire  _GEN8818 = io_x[10] ? _GEN8817 : _GEN8813;
wire  _GEN8819 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN8820 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN8821 = io_x[76] ? _GEN6833 : _GEN8820;
wire  _GEN8822 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8823 = io_x[6] ? _GEN6840 : _GEN8822;
wire  _GEN8824 = io_x[41] ? _GEN6836 : _GEN8823;
wire  _GEN8825 = io_x[14] ? _GEN6843 : _GEN8824;
wire  _GEN8826 = io_x[0] ? _GEN8825 : _GEN6845;
wire  _GEN8827 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN8828 = io_x[2] ? _GEN6837 : _GEN8827;
wire  _GEN8829 = io_x[6] ? _GEN8828 : _GEN6840;
wire  _GEN8830 = io_x[41] ? _GEN6836 : _GEN8829;
wire  _GEN8831 = io_x[14] ? _GEN6843 : _GEN8830;
wire  _GEN8832 = io_x[0] ? _GEN8831 : _GEN6845;
wire  _GEN8833 = io_x[76] ? _GEN8832 : _GEN8826;
wire  _GEN8834 = io_x[42] ? _GEN8833 : _GEN8821;
wire  _GEN8835 = io_x[38] ? _GEN8834 : _GEN8819;
wire  _GEN8836 = io_x[10] ? _GEN7044 : _GEN8835;
wire  _GEN8837 = io_x[71] ? _GEN8836 : _GEN8818;
wire  _GEN8838 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8839 = io_x[2] ? _GEN6837 : _GEN8838;
wire  _GEN8840 = io_x[6] ? _GEN6850 : _GEN8839;
wire  _GEN8841 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8842 = io_x[41] ? _GEN8841 : _GEN8840;
wire  _GEN8843 = io_x[14] ? _GEN6843 : _GEN8842;
wire  _GEN8844 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8845 = io_x[6] ? _GEN8844 : _GEN6840;
wire  _GEN8846 = io_x[41] ? _GEN8845 : _GEN6836;
wire  _GEN8847 = io_x[14] ? _GEN6843 : _GEN8846;
wire  _GEN8848 = io_x[0] ? _GEN8847 : _GEN8843;
wire  _GEN8849 = io_x[76] ? _GEN8848 : _GEN6833;
wire  _GEN8850 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8851 = io_x[41] ? _GEN6836 : _GEN8850;
wire  _GEN8852 = io_x[14] ? _GEN6843 : _GEN8851;
wire  _GEN8853 = io_x[0] ? _GEN6845 : _GEN8852;
wire  _GEN8854 = io_x[76] ? _GEN6834 : _GEN8853;
wire  _GEN8855 = io_x[42] ? _GEN8854 : _GEN8849;
wire  _GEN8856 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8857 = io_x[41] ? _GEN8856 : _GEN6924;
wire  _GEN8858 = io_x[14] ? _GEN6843 : _GEN8857;
wire  _GEN8859 = io_x[0] ? _GEN6845 : _GEN8858;
wire  _GEN8860 = io_x[76] ? _GEN8859 : _GEN6834;
wire  _GEN8861 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN8862 = io_x[14] ? _GEN6843 : _GEN8861;
wire  _GEN8863 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8864 = io_x[0] ? _GEN8863 : _GEN8862;
wire  _GEN8865 = io_x[76] ? _GEN8864 : _GEN6834;
wire  _GEN8866 = io_x[42] ? _GEN8865 : _GEN8860;
wire  _GEN8867 = io_x[38] ? _GEN8866 : _GEN8855;
wire  _GEN8868 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8869 = io_x[6] ? _GEN6850 : _GEN8868;
wire  _GEN8870 = io_x[41] ? _GEN6836 : _GEN8869;
wire  _GEN8871 = io_x[14] ? _GEN8870 : _GEN6843;
wire  _GEN8872 = io_x[0] ? _GEN6845 : _GEN8871;
wire  _GEN8873 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN8874 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN8875 = io_x[2] ? _GEN6837 : _GEN8874;
wire  _GEN8876 = io_x[6] ? _GEN8875 : _GEN6850;
wire  _GEN8877 = io_x[41] ? _GEN6924 : _GEN8876;
wire  _GEN8878 = io_x[14] ? _GEN8877 : _GEN8873;
wire  _GEN8879 = io_x[0] ? _GEN6858 : _GEN8878;
wire  _GEN8880 = io_x[76] ? _GEN8879 : _GEN8872;
wire  _GEN8881 = io_x[42] ? _GEN8880 : _GEN6874;
wire  _GEN8882 = io_x[38] ? _GEN6871 : _GEN8881;
wire  _GEN8883 = io_x[10] ? _GEN8882 : _GEN8867;
wire  _GEN8884 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN8885 = io_x[14] ? _GEN6843 : _GEN8884;
wire  _GEN8886 = io_x[0] ? _GEN8885 : _GEN6858;
wire  _GEN8887 = io_x[76] ? _GEN8886 : _GEN6834;
wire  _GEN8888 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8889 = io_x[41] ? _GEN6836 : _GEN8888;
wire  _GEN8890 = io_x[14] ? _GEN6843 : _GEN8889;
wire  _GEN8891 = io_x[0] ? _GEN6845 : _GEN8890;
wire  _GEN8892 = io_x[76] ? _GEN8891 : _GEN6834;
wire  _GEN8893 = io_x[42] ? _GEN8892 : _GEN8887;
wire  _GEN8894 = io_x[38] ? _GEN8893 : _GEN6871;
wire  _GEN8895 = io_x[10] ? _GEN7044 : _GEN8894;
wire  _GEN8896 = io_x[71] ? _GEN8895 : _GEN8883;
wire  _GEN8897 = io_x[70] ? _GEN8896 : _GEN8837;
wire  _GEN8898 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN8899 = io_x[76] ? _GEN8898 : _GEN6834;
wire  _GEN8900 = io_x[42] ? _GEN8899 : _GEN6874;
wire  _GEN8901 = io_x[38] ? _GEN8900 : _GEN6871;
wire  _GEN8902 = io_x[10] ? _GEN7044 : _GEN8901;
wire  _GEN8903 = io_x[71] ? _GEN8902 : _GEN7196;
wire  _GEN8904 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN8905 = io_x[42] ? _GEN6874 : _GEN8904;
wire  _GEN8906 = io_x[38] ? _GEN6871 : _GEN8905;
wire  _GEN8907 = io_x[10] ? _GEN7094 : _GEN8906;
wire  _GEN8908 = io_x[71] ? _GEN8907 : _GEN7196;
wire  _GEN8909 = io_x[70] ? _GEN8908 : _GEN8903;
wire  _GEN8910 = io_x[33] ? _GEN8909 : _GEN8897;
wire  _GEN8911 = io_x[21] ? _GEN8910 : _GEN8812;
wire  _GEN8912 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8913 = io_x[6] ? _GEN6850 : _GEN8912;
wire  _GEN8914 = io_x[41] ? _GEN6836 : _GEN8913;
wire  _GEN8915 = io_x[14] ? _GEN6856 : _GEN8914;
wire  _GEN8916 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8917 = io_x[41] ? _GEN6836 : _GEN8916;
wire  _GEN8918 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN8919 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8920 = io_x[6] ? _GEN8919 : _GEN8918;
wire  _GEN8921 = io_x[41] ? _GEN6836 : _GEN8920;
wire  _GEN8922 = io_x[14] ? _GEN8921 : _GEN8917;
wire  _GEN8923 = io_x[0] ? _GEN8922 : _GEN8915;
wire  _GEN8924 = io_x[76] ? _GEN6833 : _GEN8923;
wire  _GEN8925 = io_x[42] ? _GEN6874 : _GEN8924;
wire  _GEN8926 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8927 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8928 = io_x[6] ? _GEN6850 : _GEN8927;
wire  _GEN8929 = io_x[41] ? _GEN8928 : _GEN8926;
wire  _GEN8930 = io_x[14] ? _GEN6843 : _GEN8929;
wire  _GEN8931 = io_x[0] ? _GEN6845 : _GEN8930;
wire  _GEN8932 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN8933 = io_x[76] ? _GEN8932 : _GEN8931;
wire  _GEN8934 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN8935 = io_x[76] ? _GEN8934 : _GEN6834;
wire  _GEN8936 = io_x[42] ? _GEN8935 : _GEN8933;
wire  _GEN8937 = io_x[38] ? _GEN8936 : _GEN8925;
wire  _GEN8938 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8939 = io_x[0] ? _GEN8938 : _GEN6858;
wire  _GEN8940 = io_x[76] ? _GEN6834 : _GEN8939;
wire  _GEN8941 = io_x[42] ? _GEN6874 : _GEN8940;
wire  _GEN8942 = io_x[38] ? _GEN6871 : _GEN8941;
wire  _GEN8943 = io_x[10] ? _GEN8942 : _GEN8937;
wire  _GEN8944 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN8945 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN8946 = io_x[41] ? _GEN8945 : _GEN6836;
wire  _GEN8947 = io_x[14] ? _GEN6843 : _GEN8946;
wire  _GEN8948 = io_x[0] ? _GEN8947 : _GEN6858;
wire  _GEN8949 = io_x[76] ? _GEN8948 : _GEN6834;
wire  _GEN8950 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8951 = io_x[41] ? _GEN6836 : _GEN8950;
wire  _GEN8952 = io_x[14] ? _GEN6856 : _GEN8951;
wire  _GEN8953 = io_x[0] ? _GEN6845 : _GEN8952;
wire  _GEN8954 = io_x[76] ? _GEN8953 : _GEN6834;
wire  _GEN8955 = io_x[42] ? _GEN8954 : _GEN8949;
wire  _GEN8956 = io_x[38] ? _GEN8955 : _GEN8944;
wire  _GEN8957 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8958 = io_x[0] ? _GEN6858 : _GEN8957;
wire  _GEN8959 = io_x[76] ? _GEN8958 : _GEN6834;
wire  _GEN8960 = io_x[42] ? _GEN8959 : _GEN6874;
wire  _GEN8961 = io_x[38] ? _GEN8960 : _GEN6871;
wire  _GEN8962 = io_x[10] ? _GEN8961 : _GEN8956;
wire  _GEN8963 = io_x[71] ? _GEN8962 : _GEN8943;
wire  _GEN8964 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN8965 = io_x[6] ? _GEN6850 : _GEN8964;
wire  _GEN8966 = io_x[41] ? _GEN6836 : _GEN8965;
wire  _GEN8967 = io_x[14] ? _GEN6843 : _GEN8966;
wire  _GEN8968 = io_x[0] ? _GEN6845 : _GEN8967;
wire  _GEN8969 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN8970 = io_x[2] ? _GEN6837 : _GEN8969;
wire  _GEN8971 = io_x[6] ? _GEN6850 : _GEN8970;
wire  _GEN8972 = io_x[41] ? _GEN6924 : _GEN8971;
wire  _GEN8973 = io_x[14] ? _GEN6843 : _GEN8972;
wire  _GEN8974 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN8975 = io_x[0] ? _GEN8974 : _GEN8973;
wire  _GEN8976 = io_x[76] ? _GEN8975 : _GEN8968;
wire  _GEN8977 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN8978 = io_x[14] ? _GEN6843 : _GEN8977;
wire  _GEN8979 = io_x[0] ? _GEN6845 : _GEN8978;
wire  _GEN8980 = io_x[76] ? _GEN8979 : _GEN6834;
wire  _GEN8981 = io_x[42] ? _GEN8980 : _GEN8976;
wire  _GEN8982 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN8983 = io_x[41] ? _GEN6836 : _GEN8982;
wire  _GEN8984 = io_x[14] ? _GEN6856 : _GEN8983;
wire  _GEN8985 = io_x[0] ? _GEN6845 : _GEN8984;
wire  _GEN8986 = io_x[76] ? _GEN8985 : _GEN6834;
wire  _GEN8987 = io_x[42] ? _GEN8986 : _GEN6874;
wire  _GEN8988 = io_x[38] ? _GEN8987 : _GEN8981;
wire  _GEN8989 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN8990 = io_x[0] ? _GEN8989 : _GEN6845;
wire  _GEN8991 = io_x[76] ? _GEN8990 : _GEN6833;
wire  _GEN8992 = io_x[42] ? _GEN8991 : _GEN6874;
wire  _GEN8993 = io_x[38] ? _GEN6871 : _GEN8992;
wire  _GEN8994 = io_x[10] ? _GEN8993 : _GEN8988;
wire  _GEN8995 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN8996 = io_x[42] ? _GEN6863 : _GEN8995;
wire  _GEN8997 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN8998 = io_x[76] ? _GEN8997 : _GEN6834;
wire  _GEN8999 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9000 = io_x[41] ? _GEN6836 : _GEN8999;
wire  _GEN9001 = io_x[14] ? _GEN6843 : _GEN9000;
wire  _GEN9002 = io_x[0] ? _GEN6845 : _GEN9001;
wire  _GEN9003 = io_x[76] ? _GEN9002 : _GEN6834;
wire  _GEN9004 = io_x[42] ? _GEN9003 : _GEN8998;
wire  _GEN9005 = io_x[38] ? _GEN9004 : _GEN8996;
wire  _GEN9006 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9007 = io_x[6] ? _GEN9006 : _GEN6850;
wire  _GEN9008 = io_x[41] ? _GEN6836 : _GEN9007;
wire  _GEN9009 = io_x[14] ? _GEN9008 : _GEN6843;
wire  _GEN9010 = io_x[0] ? _GEN9009 : _GEN6845;
wire  _GEN9011 = io_x[76] ? _GEN9010 : _GEN6834;
wire  _GEN9012 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9013 = io_x[0] ? _GEN6845 : _GEN9012;
wire  _GEN9014 = io_x[76] ? _GEN9013 : _GEN6834;
wire  _GEN9015 = io_x[42] ? _GEN9014 : _GEN9011;
wire  _GEN9016 = io_x[38] ? _GEN9015 : _GEN6871;
wire  _GEN9017 = io_x[10] ? _GEN9016 : _GEN9005;
wire  _GEN9018 = io_x[71] ? _GEN9017 : _GEN8994;
wire  _GEN9019 = io_x[70] ? _GEN9018 : _GEN8963;
wire  _GEN9020 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9021 = io_x[41] ? _GEN6836 : _GEN9020;
wire  _GEN9022 = io_x[14] ? _GEN6856 : _GEN9021;
wire  _GEN9023 = io_x[0] ? _GEN6845 : _GEN9022;
wire  _GEN9024 = io_x[76] ? _GEN9023 : _GEN6834;
wire  _GEN9025 = io_x[42] ? _GEN9024 : _GEN6874;
wire  _GEN9026 = io_x[38] ? _GEN9025 : _GEN6871;
wire  _GEN9027 = io_x[10] ? _GEN7044 : _GEN9026;
wire  _GEN9028 = io_x[71] ? _GEN9027 : _GEN7203;
wire  _GEN9029 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN9030 = io_x[38] ? _GEN6871 : _GEN9029;
wire  _GEN9031 = io_x[10] ? _GEN7044 : _GEN9030;
wire  _GEN9032 = io_x[71] ? _GEN9031 : _GEN7196;
wire  _GEN9033 = io_x[70] ? _GEN9032 : _GEN9028;
wire  _GEN9034 = io_x[33] ? _GEN9033 : _GEN9019;
wire  _GEN9035 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9036 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9037 = io_x[41] ? _GEN9036 : _GEN9035;
wire  _GEN9038 = io_x[14] ? _GEN6843 : _GEN9037;
wire  _GEN9039 = io_x[0] ? _GEN9038 : _GEN6845;
wire  _GEN9040 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9041 = io_x[41] ? _GEN9040 : _GEN6924;
wire  _GEN9042 = io_x[14] ? _GEN6843 : _GEN9041;
wire  _GEN9043 = io_x[0] ? _GEN6858 : _GEN9042;
wire  _GEN9044 = io_x[76] ? _GEN9043 : _GEN9039;
wire  _GEN9045 = io_x[42] ? _GEN6863 : _GEN9044;
wire  _GEN9046 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN9047 = io_x[76] ? _GEN6834 : _GEN9046;
wire  _GEN9048 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9049 = io_x[2] ? _GEN6837 : _GEN9048;
wire  _GEN9050 = io_x[6] ? _GEN6850 : _GEN9049;
wire  _GEN9051 = io_x[41] ? _GEN9050 : _GEN6836;
wire  _GEN9052 = io_x[14] ? _GEN6843 : _GEN9051;
wire  _GEN9053 = io_x[0] ? _GEN6845 : _GEN9052;
wire  _GEN9054 = io_x[76] ? _GEN6834 : _GEN9053;
wire  _GEN9055 = io_x[42] ? _GEN9054 : _GEN9047;
wire  _GEN9056 = io_x[38] ? _GEN9055 : _GEN9045;
wire  _GEN9057 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9058 = io_x[41] ? _GEN6836 : _GEN9057;
wire  _GEN9059 = io_x[14] ? _GEN6843 : _GEN9058;
wire  _GEN9060 = io_x[0] ? _GEN9059 : _GEN6845;
wire  _GEN9061 = io_x[76] ? _GEN6834 : _GEN9060;
wire  _GEN9062 = io_x[42] ? _GEN6874 : _GEN9061;
wire  _GEN9063 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9064 = io_x[0] ? _GEN9063 : _GEN6845;
wire  _GEN9065 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9066 = io_x[2] ? _GEN9065 : _GEN6837;
wire  _GEN9067 = io_x[6] ? _GEN9066 : _GEN6850;
wire  _GEN9068 = io_x[41] ? _GEN6836 : _GEN9067;
wire  _GEN9069 = io_x[14] ? _GEN9068 : _GEN6843;
wire  _GEN9070 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN9071 = io_x[14] ? _GEN9070 : _GEN6843;
wire  _GEN9072 = io_x[0] ? _GEN9071 : _GEN9069;
wire  _GEN9073 = io_x[76] ? _GEN9072 : _GEN9064;
wire  _GEN9074 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9075 = io_x[6] ? _GEN9074 : _GEN6850;
wire  _GEN9076 = io_x[41] ? _GEN9075 : _GEN6836;
wire  _GEN9077 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9078 = io_x[6] ? _GEN9077 : _GEN6850;
wire  _GEN9079 = io_x[41] ? _GEN9078 : _GEN6836;
wire  _GEN9080 = io_x[14] ? _GEN9079 : _GEN9076;
wire  _GEN9081 = io_x[0] ? _GEN9080 : _GEN6845;
wire  _GEN9082 = io_x[76] ? _GEN6833 : _GEN9081;
wire  _GEN9083 = io_x[42] ? _GEN9082 : _GEN9073;
wire  _GEN9084 = io_x[38] ? _GEN9083 : _GEN9062;
wire  _GEN9085 = io_x[10] ? _GEN9084 : _GEN9056;
wire  _GEN9086 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9087 = io_x[0] ? _GEN9086 : _GEN6858;
wire  _GEN9088 = io_x[76] ? _GEN6834 : _GEN9087;
wire  _GEN9089 = io_x[42] ? _GEN6874 : _GEN9088;
wire  _GEN9090 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN9091 = io_x[76] ? _GEN6833 : _GEN9090;
wire  _GEN9092 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN9093 = io_x[14] ? _GEN6856 : _GEN9092;
wire  _GEN9094 = io_x[0] ? _GEN6858 : _GEN9093;
wire  _GEN9095 = io_x[76] ? _GEN9094 : _GEN6834;
wire  _GEN9096 = io_x[42] ? _GEN9095 : _GEN9091;
wire  _GEN9097 = io_x[38] ? _GEN9096 : _GEN9089;
wire  _GEN9098 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9099 = io_x[41] ? _GEN9098 : _GEN6836;
wire  _GEN9100 = io_x[14] ? _GEN6843 : _GEN9099;
wire  _GEN9101 = io_x[0] ? _GEN9100 : _GEN6845;
wire  _GEN9102 = io_x[76] ? _GEN9101 : _GEN6833;
wire  _GEN9103 = io_x[42] ? _GEN9102 : _GEN6863;
wire  _GEN9104 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN9105 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9106 = io_x[41] ? _GEN6836 : _GEN9105;
wire  _GEN9107 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9108 = io_x[41] ? _GEN6836 : _GEN9107;
wire  _GEN9109 = io_x[14] ? _GEN9108 : _GEN9106;
wire  _GEN9110 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9111 = io_x[0] ? _GEN9110 : _GEN9109;
wire  _GEN9112 = io_x[76] ? _GEN9111 : _GEN6834;
wire  _GEN9113 = io_x[42] ? _GEN9112 : _GEN9104;
wire  _GEN9114 = io_x[38] ? _GEN9113 : _GEN9103;
wire  _GEN9115 = io_x[10] ? _GEN9114 : _GEN9097;
wire  _GEN9116 = io_x[71] ? _GEN9115 : _GEN9085;
wire  _GEN9117 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9118 = io_x[0] ? _GEN9117 : _GEN6858;
wire  _GEN9119 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9120 = io_x[2] ? _GEN6837 : _GEN9119;
wire  _GEN9121 = io_x[6] ? _GEN6850 : _GEN9120;
wire  _GEN9122 = io_x[41] ? _GEN9121 : _GEN6924;
wire  _GEN9123 = io_x[14] ? _GEN6856 : _GEN9122;
wire  _GEN9124 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN9125 = io_x[2] ? _GEN9124 : _GEN6837;
wire  _GEN9126 = io_x[6] ? _GEN9125 : _GEN6850;
wire  _GEN9127 = io_x[41] ? _GEN9126 : _GEN6836;
wire  _GEN9128 = io_x[14] ? _GEN9127 : _GEN6843;
wire  _GEN9129 = io_x[0] ? _GEN9128 : _GEN9123;
wire  _GEN9130 = io_x[76] ? _GEN9129 : _GEN9118;
wire  _GEN9131 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9132 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9133 = io_x[41] ? _GEN9132 : _GEN9131;
wire  _GEN9134 = io_x[14] ? _GEN6843 : _GEN9133;
wire  _GEN9135 = io_x[0] ? _GEN9134 : _GEN6858;
wire  _GEN9136 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN9137 = io_x[14] ? _GEN6843 : _GEN9136;
wire  _GEN9138 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN9139 = io_x[14] ? _GEN6843 : _GEN9138;
wire  _GEN9140 = io_x[0] ? _GEN9139 : _GEN9137;
wire  _GEN9141 = io_x[76] ? _GEN9140 : _GEN9135;
wire  _GEN9142 = io_x[42] ? _GEN9141 : _GEN9130;
wire  _GEN9143 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN9144 = io_x[14] ? _GEN6843 : _GEN9143;
wire  _GEN9145 = io_x[0] ? _GEN6845 : _GEN9144;
wire  _GEN9146 = io_x[76] ? _GEN6833 : _GEN9145;
wire  _GEN9147 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9148 = io_x[6] ? _GEN6850 : _GEN9147;
wire  _GEN9149 = io_x[41] ? _GEN6836 : _GEN9148;
wire  _GEN9150 = io_x[14] ? _GEN6843 : _GEN9149;
wire  _GEN9151 = io_x[0] ? _GEN6858 : _GEN9150;
wire  _GEN9152 = io_x[76] ? _GEN9151 : _GEN6834;
wire  _GEN9153 = io_x[42] ? _GEN9152 : _GEN9146;
wire  _GEN9154 = io_x[38] ? _GEN9153 : _GEN9142;
wire  _GEN9155 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9156 = io_x[6] ? _GEN9155 : _GEN6850;
wire  _GEN9157 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9158 = io_x[41] ? _GEN9157 : _GEN9156;
wire  _GEN9159 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9160 = io_x[6] ? _GEN9159 : _GEN6850;
wire  _GEN9161 = io_x[41] ? _GEN6924 : _GEN9160;
wire  _GEN9162 = io_x[14] ? _GEN9161 : _GEN9158;
wire  _GEN9163 = io_x[0] ? _GEN9162 : _GEN6845;
wire  _GEN9164 = io_x[76] ? _GEN6834 : _GEN9163;
wire  _GEN9165 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9166 = io_x[41] ? _GEN9165 : _GEN6924;
wire  _GEN9167 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN9168 = io_x[2] ? _GEN9167 : _GEN6837;
wire  _GEN9169 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9170 = io_x[2] ? _GEN9169 : _GEN6837;
wire  _GEN9171 = io_x[6] ? _GEN9170 : _GEN9168;
wire  _GEN9172 = io_x[41] ? _GEN9171 : _GEN6836;
wire  _GEN9173 = io_x[14] ? _GEN9172 : _GEN9166;
wire  _GEN9174 = io_x[0] ? _GEN9173 : _GEN6858;
wire  _GEN9175 = io_x[76] ? _GEN9174 : _GEN6834;
wire  _GEN9176 = io_x[42] ? _GEN9175 : _GEN9164;
wire  _GEN9177 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN9178 = io_x[14] ? _GEN6843 : _GEN9177;
wire  _GEN9179 = io_x[0] ? _GEN9178 : _GEN6858;
wire  _GEN9180 = io_x[76] ? _GEN9179 : _GEN6833;
wire  _GEN9181 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN9182 = io_x[14] ? _GEN9181 : _GEN6843;
wire  _GEN9183 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9184 = io_x[2] ? _GEN9183 : _GEN6837;
wire  _GEN9185 = io_x[6] ? _GEN9184 : _GEN6850;
wire  _GEN9186 = io_x[41] ? _GEN6836 : _GEN9185;
wire  _GEN9187 = io_x[14] ? _GEN9186 : _GEN6843;
wire  _GEN9188 = io_x[0] ? _GEN9187 : _GEN9182;
wire  _GEN9189 = io_x[76] ? _GEN9188 : _GEN6834;
wire  _GEN9190 = io_x[42] ? _GEN9189 : _GEN9180;
wire  _GEN9191 = io_x[38] ? _GEN9190 : _GEN9176;
wire  _GEN9192 = io_x[10] ? _GEN9191 : _GEN9154;
wire  _GEN9193 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9194 = io_x[0] ? _GEN9193 : _GEN6845;
wire  _GEN9195 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9196 = io_x[2] ? _GEN6837 : _GEN9195;
wire  _GEN9197 = io_x[6] ? _GEN6850 : _GEN9196;
wire  _GEN9198 = io_x[41] ? _GEN6836 : _GEN9197;
wire  _GEN9199 = io_x[14] ? _GEN6843 : _GEN9198;
wire  _GEN9200 = io_x[0] ? _GEN6845 : _GEN9199;
wire  _GEN9201 = io_x[76] ? _GEN9200 : _GEN9194;
wire  _GEN9202 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9203 = io_x[2] ? _GEN6837 : _GEN9202;
wire  _GEN9204 = io_x[6] ? _GEN6850 : _GEN9203;
wire  _GEN9205 = io_x[41] ? _GEN6836 : _GEN9204;
wire  _GEN9206 = io_x[14] ? _GEN6843 : _GEN9205;
wire  _GEN9207 = io_x[0] ? _GEN6845 : _GEN9206;
wire  _GEN9208 = io_x[76] ? _GEN9207 : _GEN6834;
wire  _GEN9209 = io_x[42] ? _GEN9208 : _GEN9201;
wire  _GEN9210 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN9211 = io_x[76] ? _GEN6833 : _GEN9210;
wire  _GEN9212 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN9213 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9214 = io_x[41] ? _GEN6836 : _GEN9213;
wire  _GEN9215 = io_x[14] ? _GEN6856 : _GEN9214;
wire  _GEN9216 = io_x[0] ? _GEN6845 : _GEN9215;
wire  _GEN9217 = io_x[76] ? _GEN9216 : _GEN9212;
wire  _GEN9218 = io_x[42] ? _GEN9217 : _GEN9211;
wire  _GEN9219 = io_x[38] ? _GEN9218 : _GEN9209;
wire  _GEN9220 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN9221 = io_x[14] ? _GEN9220 : _GEN6843;
wire  _GEN9222 = io_x[0] ? _GEN9221 : _GEN6845;
wire  _GEN9223 = io_x[76] ? _GEN6833 : _GEN9222;
wire  _GEN9224 = io_x[42] ? _GEN6874 : _GEN9223;
wire  _GEN9225 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9226 = io_x[2] ? _GEN9225 : _GEN6837;
wire  _GEN9227 = io_x[6] ? _GEN9226 : _GEN6850;
wire  _GEN9228 = io_x[41] ? _GEN6836 : _GEN9227;
wire  _GEN9229 = io_x[14] ? _GEN9228 : _GEN6843;
wire  _GEN9230 = io_x[0] ? _GEN9229 : _GEN6845;
wire  _GEN9231 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9232 = io_x[0] ? _GEN9231 : _GEN6845;
wire  _GEN9233 = io_x[76] ? _GEN9232 : _GEN9230;
wire  _GEN9234 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9235 = io_x[41] ? _GEN6836 : _GEN9234;
wire  _GEN9236 = io_x[14] ? _GEN9235 : _GEN6843;
wire  _GEN9237 = io_x[0] ? _GEN9236 : _GEN6858;
wire  _GEN9238 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9239 = io_x[41] ? _GEN6836 : _GEN9238;
wire  _GEN9240 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9241 = io_x[41] ? _GEN6836 : _GEN9240;
wire  _GEN9242 = io_x[14] ? _GEN9241 : _GEN9239;
wire  _GEN9243 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9244 = io_x[41] ? _GEN9243 : _GEN6836;
wire  _GEN9245 = io_x[14] ? _GEN9244 : _GEN6856;
wire  _GEN9246 = io_x[0] ? _GEN9245 : _GEN9242;
wire  _GEN9247 = io_x[76] ? _GEN9246 : _GEN9237;
wire  _GEN9248 = io_x[42] ? _GEN9247 : _GEN9233;
wire  _GEN9249 = io_x[38] ? _GEN9248 : _GEN9224;
wire  _GEN9250 = io_x[10] ? _GEN9249 : _GEN9219;
wire  _GEN9251 = io_x[71] ? _GEN9250 : _GEN9192;
wire  _GEN9252 = io_x[70] ? _GEN9251 : _GEN9116;
wire  _GEN9253 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN9254 = io_x[10] ? _GEN9253 : _GEN7094;
wire  _GEN9255 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9256 = io_x[6] ? _GEN6850 : _GEN9255;
wire  _GEN9257 = io_x[41] ? _GEN6836 : _GEN9256;
wire  _GEN9258 = io_x[14] ? _GEN6843 : _GEN9257;
wire  _GEN9259 = io_x[0] ? _GEN6845 : _GEN9258;
wire  _GEN9260 = io_x[76] ? _GEN9259 : _GEN6834;
wire  _GEN9261 = io_x[42] ? _GEN9260 : _GEN6874;
wire  _GEN9262 = io_x[38] ? _GEN9261 : _GEN6871;
wire  _GEN9263 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9264 = io_x[0] ? _GEN6845 : _GEN9263;
wire  _GEN9265 = io_x[76] ? _GEN9264 : _GEN6834;
wire  _GEN9266 = io_x[42] ? _GEN9265 : _GEN6874;
wire  _GEN9267 = io_x[38] ? _GEN9266 : _GEN6871;
wire  _GEN9268 = io_x[10] ? _GEN9267 : _GEN9262;
wire  _GEN9269 = io_x[71] ? _GEN9268 : _GEN9254;
wire  _GEN9270 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9271 = io_x[6] ? _GEN9270 : _GEN6850;
wire  _GEN9272 = io_x[41] ? _GEN6836 : _GEN9271;
wire  _GEN9273 = io_x[14] ? _GEN9272 : _GEN6843;
wire  _GEN9274 = io_x[0] ? _GEN9273 : _GEN6858;
wire  _GEN9275 = io_x[76] ? _GEN9274 : _GEN6833;
wire  _GEN9276 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9277 = io_x[6] ? _GEN9276 : _GEN6850;
wire  _GEN9278 = io_x[41] ? _GEN9277 : _GEN6836;
wire  _GEN9279 = io_x[14] ? _GEN9278 : _GEN6843;
wire  _GEN9280 = io_x[0] ? _GEN9279 : _GEN6845;
wire  _GEN9281 = io_x[76] ? _GEN9280 : _GEN6834;
wire  _GEN9282 = io_x[42] ? _GEN9281 : _GEN9275;
wire  _GEN9283 = io_x[38] ? _GEN9282 : _GEN6871;
wire  _GEN9284 = io_x[10] ? _GEN9283 : _GEN7044;
wire  _GEN9285 = io_x[71] ? _GEN9284 : _GEN7196;
wire  _GEN9286 = io_x[70] ? _GEN9285 : _GEN9269;
wire  _GEN9287 = io_x[33] ? _GEN9286 : _GEN9252;
wire  _GEN9288 = io_x[21] ? _GEN9287 : _GEN9034;
wire  _GEN9289 = io_x[18] ? _GEN9288 : _GEN8911;
wire  _GEN9290 = io_x[20] ? _GEN9289 : _GEN8731;
wire  _GEN9291 = io_x[45] ? _GEN9290 : _GEN8263;
wire  _GEN9292 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9293 = io_x[6] ? _GEN6850 : _GEN9292;
wire  _GEN9294 = io_x[41] ? _GEN9293 : _GEN6836;
wire  _GEN9295 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9296 = io_x[41] ? _GEN9295 : _GEN6836;
wire  _GEN9297 = io_x[14] ? _GEN9296 : _GEN9294;
wire  _GEN9298 = io_x[0] ? _GEN6845 : _GEN9297;
wire  _GEN9299 = io_x[76] ? _GEN6833 : _GEN9298;
wire  _GEN9300 = io_x[42] ? _GEN9299 : _GEN6874;
wire  _GEN9301 = io_x[38] ? _GEN6871 : _GEN9300;
wire  _GEN9302 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9303 = io_x[2] ? _GEN9302 : _GEN6837;
wire  _GEN9304 = io_x[6] ? _GEN6840 : _GEN9303;
wire  _GEN9305 = io_x[41] ? _GEN9304 : _GEN6836;
wire  _GEN9306 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9307 = io_x[6] ? _GEN9306 : _GEN6850;
wire  _GEN9308 = io_x[41] ? _GEN9307 : _GEN6836;
wire  _GEN9309 = io_x[14] ? _GEN9308 : _GEN9305;
wire  _GEN9310 = io_x[0] ? _GEN6845 : _GEN9309;
wire  _GEN9311 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9312 = io_x[0] ? _GEN6845 : _GEN9311;
wire  _GEN9313 = io_x[76] ? _GEN9312 : _GEN9310;
wire  _GEN9314 = io_x[42] ? _GEN9313 : _GEN6874;
wire  _GEN9315 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9316 = io_x[0] ? _GEN6858 : _GEN9315;
wire  _GEN9317 = io_x[76] ? _GEN6834 : _GEN9316;
wire  _GEN9318 = io_x[42] ? _GEN9317 : _GEN6874;
wire  _GEN9319 = io_x[38] ? _GEN9318 : _GEN9314;
wire  _GEN9320 = io_x[10] ? _GEN9319 : _GEN9301;
wire  _GEN9321 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN9322 = io_x[42] ? _GEN9321 : _GEN6874;
wire  _GEN9323 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9324 = io_x[41] ? _GEN6836 : _GEN9323;
wire  _GEN9325 = io_x[14] ? _GEN9324 : _GEN6843;
wire  _GEN9326 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9327 = io_x[0] ? _GEN9326 : _GEN9325;
wire  _GEN9328 = io_x[76] ? _GEN9327 : _GEN6834;
wire  _GEN9329 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN9330 = io_x[76] ? _GEN6834 : _GEN9329;
wire  _GEN9331 = io_x[42] ? _GEN9330 : _GEN9328;
wire  _GEN9332 = io_x[38] ? _GEN9331 : _GEN9322;
wire  _GEN9333 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN9334 = io_x[76] ? _GEN6833 : _GEN9333;
wire  _GEN9335 = io_x[42] ? _GEN9334 : _GEN6863;
wire  _GEN9336 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9337 = io_x[41] ? _GEN6836 : _GEN9336;
wire  _GEN9338 = io_x[14] ? _GEN6843 : _GEN9337;
wire  _GEN9339 = io_x[0] ? _GEN6845 : _GEN9338;
wire  _GEN9340 = io_x[76] ? _GEN9339 : _GEN6833;
wire  _GEN9341 = io_x[42] ? _GEN6874 : _GEN9340;
wire  _GEN9342 = io_x[38] ? _GEN9341 : _GEN9335;
wire  _GEN9343 = io_x[10] ? _GEN9342 : _GEN9332;
wire  _GEN9344 = io_x[71] ? _GEN9343 : _GEN9320;
wire  _GEN9345 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN9346 = io_x[14] ? _GEN6843 : _GEN9345;
wire  _GEN9347 = io_x[0] ? _GEN6858 : _GEN9346;
wire  _GEN9348 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9349 = io_x[41] ? _GEN6924 : _GEN9348;
wire  _GEN9350 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9351 = io_x[41] ? _GEN6924 : _GEN9350;
wire  _GEN9352 = io_x[14] ? _GEN9351 : _GEN9349;
wire  _GEN9353 = io_x[0] ? _GEN6845 : _GEN9352;
wire  _GEN9354 = io_x[76] ? _GEN9353 : _GEN9347;
wire  _GEN9355 = io_x[42] ? _GEN9354 : _GEN6874;
wire  _GEN9356 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9357 = io_x[0] ? _GEN6845 : _GEN9356;
wire  _GEN9358 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN9359 = io_x[76] ? _GEN9358 : _GEN9357;
wire  _GEN9360 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9361 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9362 = io_x[2] ? _GEN6837 : _GEN9361;
wire  _GEN9363 = io_x[6] ? _GEN6850 : _GEN9362;
wire  _GEN9364 = io_x[41] ? _GEN9363 : _GEN9360;
wire  _GEN9365 = io_x[14] ? _GEN6843 : _GEN9364;
wire  _GEN9366 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9367 = io_x[41] ? _GEN6836 : _GEN9366;
wire  _GEN9368 = io_x[14] ? _GEN9367 : _GEN6843;
wire  _GEN9369 = io_x[0] ? _GEN9368 : _GEN9365;
wire  _GEN9370 = io_x[76] ? _GEN6833 : _GEN9369;
wire  _GEN9371 = io_x[42] ? _GEN9370 : _GEN9359;
wire  _GEN9372 = io_x[38] ? _GEN9371 : _GEN9355;
wire  _GEN9373 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9374 = io_x[6] ? _GEN9373 : _GEN6850;
wire  _GEN9375 = io_x[41] ? _GEN6836 : _GEN9374;
wire  _GEN9376 = io_x[14] ? _GEN6856 : _GEN9375;
wire  _GEN9377 = io_x[0] ? _GEN9376 : _GEN6845;
wire  _GEN9378 = io_x[76] ? _GEN9377 : _GEN6834;
wire  _GEN9379 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9380 = io_x[41] ? _GEN6836 : _GEN9379;
wire  _GEN9381 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9382 = io_x[41] ? _GEN6836 : _GEN9381;
wire  _GEN9383 = io_x[14] ? _GEN9382 : _GEN9380;
wire  _GEN9384 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN9385 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9386 = io_x[6] ? _GEN9385 : _GEN6850;
wire  _GEN9387 = io_x[41] ? _GEN6836 : _GEN9386;
wire  _GEN9388 = io_x[14] ? _GEN9387 : _GEN9384;
wire  _GEN9389 = io_x[0] ? _GEN9388 : _GEN9383;
wire  _GEN9390 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9391 = io_x[41] ? _GEN9390 : _GEN6924;
wire  _GEN9392 = io_x[14] ? _GEN9391 : _GEN6856;
wire  _GEN9393 = io_x[0] ? _GEN6845 : _GEN9392;
wire  _GEN9394 = io_x[76] ? _GEN9393 : _GEN9389;
wire  _GEN9395 = io_x[42] ? _GEN9394 : _GEN9378;
wire  _GEN9396 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9397 = io_x[6] ? _GEN9396 : _GEN6850;
wire  _GEN9398 = io_x[41] ? _GEN9397 : _GEN6924;
wire  _GEN9399 = io_x[14] ? _GEN9398 : _GEN6856;
wire  _GEN9400 = io_x[0] ? _GEN6845 : _GEN9399;
wire  _GEN9401 = io_x[76] ? _GEN6834 : _GEN9400;
wire  _GEN9402 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9403 = io_x[6] ? _GEN9402 : _GEN6850;
wire  _GEN9404 = io_x[41] ? _GEN6836 : _GEN9403;
wire  _GEN9405 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9406 = io_x[41] ? _GEN6836 : _GEN9405;
wire  _GEN9407 = io_x[14] ? _GEN9406 : _GEN9404;
wire  _GEN9408 = io_x[0] ? _GEN6845 : _GEN9407;
wire  _GEN9409 = io_x[76] ? _GEN6833 : _GEN9408;
wire  _GEN9410 = io_x[42] ? _GEN9409 : _GEN9401;
wire  _GEN9411 = io_x[38] ? _GEN9410 : _GEN9395;
wire  _GEN9412 = io_x[10] ? _GEN9411 : _GEN9372;
wire  _GEN9413 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN9414 = io_x[76] ? _GEN6834 : _GEN9413;
wire  _GEN9415 = io_x[42] ? _GEN6863 : _GEN9414;
wire  _GEN9416 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9417 = io_x[41] ? _GEN6836 : _GEN9416;
wire  _GEN9418 = io_x[14] ? _GEN9417 : _GEN6843;
wire  _GEN9419 = io_x[0] ? _GEN6858 : _GEN9418;
wire  _GEN9420 = io_x[76] ? _GEN6834 : _GEN9419;
wire  _GEN9421 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9422 = io_x[2] ? _GEN6837 : _GEN9421;
wire  _GEN9423 = io_x[6] ? _GEN6850 : _GEN9422;
wire  _GEN9424 = io_x[41] ? _GEN9423 : _GEN6836;
wire  _GEN9425 = io_x[14] ? _GEN6843 : _GEN9424;
wire  _GEN9426 = io_x[0] ? _GEN6845 : _GEN9425;
wire  _GEN9427 = io_x[76] ? _GEN6833 : _GEN9426;
wire  _GEN9428 = io_x[42] ? _GEN9427 : _GEN9420;
wire  _GEN9429 = io_x[38] ? _GEN9428 : _GEN9415;
wire  _GEN9430 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9431 = io_x[41] ? _GEN9430 : _GEN6924;
wire  _GEN9432 = io_x[14] ? _GEN6856 : _GEN9431;
wire  _GEN9433 = io_x[0] ? _GEN6845 : _GEN9432;
wire  _GEN9434 = io_x[76] ? _GEN6834 : _GEN9433;
wire  _GEN9435 = io_x[42] ? _GEN6874 : _GEN9434;
wire  _GEN9436 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9437 = io_x[6] ? _GEN9436 : _GEN6850;
wire  _GEN9438 = io_x[41] ? _GEN6924 : _GEN9437;
wire  _GEN9439 = io_x[14] ? _GEN9438 : _GEN6856;
wire  _GEN9440 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9441 = io_x[41] ? _GEN9440 : _GEN6836;
wire  _GEN9442 = io_x[14] ? _GEN9441 : _GEN6843;
wire  _GEN9443 = io_x[0] ? _GEN9442 : _GEN9439;
wire  _GEN9444 = io_x[76] ? _GEN6834 : _GEN9443;
wire  _GEN9445 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9446 = io_x[41] ? _GEN6836 : _GEN9445;
wire  _GEN9447 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9448 = io_x[41] ? _GEN6836 : _GEN9447;
wire  _GEN9449 = io_x[14] ? _GEN9448 : _GEN9446;
wire  _GEN9450 = io_x[0] ? _GEN6845 : _GEN9449;
wire  _GEN9451 = io_x[76] ? _GEN6833 : _GEN9450;
wire  _GEN9452 = io_x[42] ? _GEN9451 : _GEN9444;
wire  _GEN9453 = io_x[38] ? _GEN9452 : _GEN9435;
wire  _GEN9454 = io_x[10] ? _GEN9453 : _GEN9429;
wire  _GEN9455 = io_x[71] ? _GEN9454 : _GEN9412;
wire  _GEN9456 = io_x[70] ? _GEN9455 : _GEN9344;
wire  _GEN9457 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9458 = io_x[0] ? _GEN6845 : _GEN9457;
wire  _GEN9459 = io_x[76] ? _GEN6834 : _GEN9458;
wire  _GEN9460 = io_x[42] ? _GEN9459 : _GEN6874;
wire  _GEN9461 = io_x[38] ? _GEN9460 : _GEN6871;
wire  _GEN9462 = io_x[10] ? _GEN9461 : _GEN7044;
wire  _GEN9463 = io_x[71] ? _GEN9462 : _GEN7196;
wire  _GEN9464 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9465 = io_x[41] ? _GEN9464 : _GEN6836;
wire  _GEN9466 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9467 = io_x[41] ? _GEN9466 : _GEN6836;
wire  _GEN9468 = io_x[14] ? _GEN9467 : _GEN9465;
wire  _GEN9469 = io_x[0] ? _GEN9468 : _GEN6845;
wire  _GEN9470 = io_x[76] ? _GEN9469 : _GEN6834;
wire  _GEN9471 = io_x[42] ? _GEN6874 : _GEN9470;
wire  _GEN9472 = io_x[38] ? _GEN9471 : _GEN6871;
wire  _GEN9473 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9474 = io_x[41] ? _GEN9473 : _GEN6836;
wire  _GEN9475 = io_x[14] ? _GEN9474 : _GEN6843;
wire  _GEN9476 = io_x[0] ? _GEN9475 : _GEN6845;
wire  _GEN9477 = io_x[76] ? _GEN9476 : _GEN6834;
wire  _GEN9478 = io_x[42] ? _GEN6874 : _GEN9477;
wire  _GEN9479 = io_x[38] ? _GEN9478 : _GEN7036;
wire  _GEN9480 = io_x[10] ? _GEN9479 : _GEN9472;
wire  _GEN9481 = io_x[71] ? _GEN7203 : _GEN9480;
wire  _GEN9482 = io_x[70] ? _GEN9481 : _GEN9463;
wire  _GEN9483 = io_x[33] ? _GEN9482 : _GEN9456;
wire  _GEN9484 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN9485 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9486 = io_x[41] ? _GEN9485 : _GEN6836;
wire  _GEN9487 = io_x[14] ? _GEN9486 : _GEN6856;
wire  _GEN9488 = io_x[0] ? _GEN6845 : _GEN9487;
wire  _GEN9489 = io_x[76] ? _GEN6834 : _GEN9488;
wire  _GEN9490 = io_x[42] ? _GEN9489 : _GEN9484;
wire  _GEN9491 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9492 = io_x[0] ? _GEN9491 : _GEN6845;
wire  _GEN9493 = io_x[76] ? _GEN9492 : _GEN6834;
wire  _GEN9494 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN9495 = io_x[42] ? _GEN9494 : _GEN9493;
wire  _GEN9496 = io_x[38] ? _GEN9495 : _GEN9490;
wire  _GEN9497 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN9498 = io_x[2] ? _GEN9497 : _GEN6837;
wire  _GEN9499 = io_x[6] ? _GEN9498 : _GEN6850;
wire  _GEN9500 = io_x[41] ? _GEN9499 : _GEN6836;
wire  _GEN9501 = io_x[14] ? _GEN6856 : _GEN9500;
wire  _GEN9502 = io_x[0] ? _GEN6845 : _GEN9501;
wire  _GEN9503 = io_x[76] ? _GEN6833 : _GEN9502;
wire  _GEN9504 = io_x[42] ? _GEN9503 : _GEN6874;
wire  _GEN9505 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9506 = io_x[41] ? _GEN6836 : _GEN9505;
wire  _GEN9507 = io_x[14] ? _GEN6856 : _GEN9506;
wire  _GEN9508 = io_x[0] ? _GEN9507 : _GEN6845;
wire  _GEN9509 = io_x[76] ? _GEN9508 : _GEN6834;
wire  _GEN9510 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9511 = io_x[41] ? _GEN6836 : _GEN9510;
wire  _GEN9512 = io_x[14] ? _GEN9511 : _GEN6843;
wire  _GEN9513 = io_x[0] ? _GEN6845 : _GEN9512;
wire  _GEN9514 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN9515 = io_x[76] ? _GEN9514 : _GEN9513;
wire  _GEN9516 = io_x[42] ? _GEN9515 : _GEN9509;
wire  _GEN9517 = io_x[38] ? _GEN9516 : _GEN9504;
wire  _GEN9518 = io_x[10] ? _GEN9517 : _GEN9496;
wire  _GEN9519 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN9520 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN9521 = io_x[42] ? _GEN9520 : _GEN9519;
wire  _GEN9522 = io_x[38] ? _GEN9521 : _GEN7036;
wire  _GEN9523 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN9524 = io_x[76] ? _GEN6833 : _GEN9523;
wire  _GEN9525 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9526 = io_x[41] ? _GEN9525 : _GEN6836;
wire  _GEN9527 = io_x[14] ? _GEN9526 : _GEN6843;
wire  _GEN9528 = io_x[0] ? _GEN6845 : _GEN9527;
wire  _GEN9529 = io_x[76] ? _GEN6834 : _GEN9528;
wire  _GEN9530 = io_x[42] ? _GEN9529 : _GEN9524;
wire  _GEN9531 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN9532 = io_x[14] ? _GEN9531 : _GEN6843;
wire  _GEN9533 = io_x[0] ? _GEN6845 : _GEN9532;
wire  _GEN9534 = io_x[76] ? _GEN6834 : _GEN9533;
wire  _GEN9535 = io_x[42] ? _GEN6874 : _GEN9534;
wire  _GEN9536 = io_x[38] ? _GEN9535 : _GEN9530;
wire  _GEN9537 = io_x[10] ? _GEN9536 : _GEN9522;
wire  _GEN9538 = io_x[71] ? _GEN9537 : _GEN9518;
wire  _GEN9539 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9540 = io_x[0] ? _GEN9539 : _GEN6845;
wire  _GEN9541 = io_x[76] ? _GEN6833 : _GEN9540;
wire  _GEN9542 = io_x[42] ? _GEN9541 : _GEN6874;
wire  _GEN9543 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9544 = io_x[41] ? _GEN6836 : _GEN9543;
wire  _GEN9545 = io_x[14] ? _GEN6843 : _GEN9544;
wire  _GEN9546 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9547 = io_x[0] ? _GEN9546 : _GEN9545;
wire  _GEN9548 = io_x[76] ? _GEN9547 : _GEN6833;
wire  _GEN9549 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN9550 = io_x[42] ? _GEN9549 : _GEN9548;
wire  _GEN9551 = io_x[38] ? _GEN9550 : _GEN9542;
wire  _GEN9552 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN9553 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9554 = io_x[41] ? _GEN6836 : _GEN9553;
wire  _GEN9555 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9556 = io_x[41] ? _GEN6836 : _GEN9555;
wire  _GEN9557 = io_x[14] ? _GEN9556 : _GEN9554;
wire  _GEN9558 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9559 = io_x[6] ? _GEN6840 : _GEN9558;
wire  _GEN9560 = io_x[41] ? _GEN6836 : _GEN9559;
wire  _GEN9561 = io_x[14] ? _GEN9560 : _GEN6843;
wire  _GEN9562 = io_x[0] ? _GEN9561 : _GEN9557;
wire  _GEN9563 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN9564 = io_x[2] ? _GEN6837 : _GEN9563;
wire  _GEN9565 = io_x[6] ? _GEN6840 : _GEN9564;
wire  _GEN9566 = io_x[41] ? _GEN9565 : _GEN6836;
wire  _GEN9567 = io_x[14] ? _GEN6843 : _GEN9566;
wire  _GEN9568 = io_x[0] ? _GEN6845 : _GEN9567;
wire  _GEN9569 = io_x[76] ? _GEN9568 : _GEN9562;
wire  _GEN9570 = io_x[42] ? _GEN9569 : _GEN9552;
wire  _GEN9571 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9572 = io_x[41] ? _GEN6836 : _GEN9571;
wire  _GEN9573 = io_x[14] ? _GEN9572 : _GEN6856;
wire  _GEN9574 = io_x[0] ? _GEN6845 : _GEN9573;
wire  _GEN9575 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9576 = io_x[41] ? _GEN6836 : _GEN9575;
wire  _GEN9577 = io_x[14] ? _GEN6856 : _GEN9576;
wire  _GEN9578 = io_x[0] ? _GEN9577 : _GEN6845;
wire  _GEN9579 = io_x[76] ? _GEN9578 : _GEN9574;
wire  _GEN9580 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9581 = io_x[41] ? _GEN6836 : _GEN9580;
wire  _GEN9582 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9583 = io_x[41] ? _GEN6836 : _GEN9582;
wire  _GEN9584 = io_x[14] ? _GEN9583 : _GEN9581;
wire  _GEN9585 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9586 = io_x[41] ? _GEN6836 : _GEN9585;
wire  _GEN9587 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9588 = io_x[41] ? _GEN6836 : _GEN9587;
wire  _GEN9589 = io_x[14] ? _GEN9588 : _GEN9586;
wire  _GEN9590 = io_x[0] ? _GEN9589 : _GEN9584;
wire  _GEN9591 = io_x[76] ? _GEN6833 : _GEN9590;
wire  _GEN9592 = io_x[42] ? _GEN9591 : _GEN9579;
wire  _GEN9593 = io_x[38] ? _GEN9592 : _GEN9570;
wire  _GEN9594 = io_x[10] ? _GEN9593 : _GEN9551;
wire  _GEN9595 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9596 = io_x[0] ? _GEN6845 : _GEN9595;
wire  _GEN9597 = io_x[76] ? _GEN6834 : _GEN9596;
wire  _GEN9598 = io_x[42] ? _GEN6863 : _GEN9597;
wire  _GEN9599 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9600 = io_x[41] ? _GEN6836 : _GEN9599;
wire  _GEN9601 = io_x[14] ? _GEN6843 : _GEN9600;
wire  _GEN9602 = io_x[0] ? _GEN6858 : _GEN9601;
wire  _GEN9603 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9604 = io_x[6] ? _GEN6850 : _GEN9603;
wire  _GEN9605 = io_x[41] ? _GEN9604 : _GEN6836;
wire  _GEN9606 = io_x[14] ? _GEN9605 : _GEN6843;
wire  _GEN9607 = io_x[0] ? _GEN9606 : _GEN6845;
wire  _GEN9608 = io_x[76] ? _GEN9607 : _GEN9602;
wire  _GEN9609 = io_x[42] ? _GEN9608 : _GEN6863;
wire  _GEN9610 = io_x[38] ? _GEN9609 : _GEN9598;
wire  _GEN9611 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9612 = io_x[0] ? _GEN6845 : _GEN9611;
wire  _GEN9613 = io_x[76] ? _GEN6833 : _GEN9612;
wire  _GEN9614 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN9615 = io_x[76] ? _GEN9614 : _GEN6833;
wire  _GEN9616 = io_x[42] ? _GEN9615 : _GEN9613;
wire  _GEN9617 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9618 = io_x[41] ? _GEN6836 : _GEN9617;
wire  _GEN9619 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9620 = io_x[41] ? _GEN6836 : _GEN9619;
wire  _GEN9621 = io_x[14] ? _GEN9620 : _GEN9618;
wire  _GEN9622 = io_x[0] ? _GEN6845 : _GEN9621;
wire  _GEN9623 = io_x[76] ? _GEN6834 : _GEN9622;
wire  _GEN9624 = io_x[42] ? _GEN9623 : _GEN6863;
wire  _GEN9625 = io_x[38] ? _GEN9624 : _GEN9616;
wire  _GEN9626 = io_x[10] ? _GEN9625 : _GEN9610;
wire  _GEN9627 = io_x[71] ? _GEN9626 : _GEN9594;
wire  _GEN9628 = io_x[70] ? _GEN9627 : _GEN9538;
wire  _GEN9629 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9630 = io_x[0] ? _GEN6845 : _GEN9629;
wire  _GEN9631 = io_x[76] ? _GEN6834 : _GEN9630;
wire  _GEN9632 = io_x[42] ? _GEN9631 : _GEN6863;
wire  _GEN9633 = io_x[38] ? _GEN9632 : _GEN6871;
wire  _GEN9634 = io_x[10] ? _GEN9633 : _GEN7044;
wire  _GEN9635 = io_x[71] ? _GEN7196 : _GEN9634;
wire  _GEN9636 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9637 = io_x[41] ? _GEN6836 : _GEN9636;
wire  _GEN9638 = io_x[14] ? _GEN9637 : _GEN6843;
wire  _GEN9639 = io_x[0] ? _GEN6845 : _GEN9638;
wire  _GEN9640 = io_x[76] ? _GEN6834 : _GEN9639;
wire  _GEN9641 = io_x[42] ? _GEN9640 : _GEN6874;
wire  _GEN9642 = io_x[38] ? _GEN9641 : _GEN6871;
wire  _GEN9643 = io_x[10] ? _GEN9642 : _GEN7044;
wire  _GEN9644 = io_x[71] ? _GEN9643 : _GEN7203;
wire  _GEN9645 = io_x[70] ? _GEN9644 : _GEN9635;
wire  _GEN9646 = io_x[33] ? _GEN9645 : _GEN9628;
wire  _GEN9647 = io_x[21] ? _GEN9646 : _GEN9483;
wire  _GEN9648 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN9649 = io_x[76] ? _GEN9648 : _GEN6834;
wire  _GEN9650 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9651 = io_x[41] ? _GEN6836 : _GEN9650;
wire  _GEN9652 = io_x[14] ? _GEN9651 : _GEN6856;
wire  _GEN9653 = io_x[0] ? _GEN9652 : _GEN6858;
wire  _GEN9654 = io_x[76] ? _GEN6834 : _GEN9653;
wire  _GEN9655 = io_x[42] ? _GEN9654 : _GEN9649;
wire  _GEN9656 = io_x[38] ? _GEN9655 : _GEN7036;
wire  _GEN9657 = io_x[10] ? _GEN9656 : _GEN7044;
wire  _GEN9658 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9659 = io_x[6] ? _GEN9658 : _GEN6850;
wire  _GEN9660 = io_x[41] ? _GEN9659 : _GEN6836;
wire  _GEN9661 = io_x[14] ? _GEN9660 : _GEN6843;
wire  _GEN9662 = io_x[0] ? _GEN9661 : _GEN6858;
wire  _GEN9663 = io_x[76] ? _GEN6834 : _GEN9662;
wire  _GEN9664 = io_x[42] ? _GEN9663 : _GEN6874;
wire  _GEN9665 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN9666 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9667 = io_x[0] ? _GEN6845 : _GEN9666;
wire  _GEN9668 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9669 = io_x[6] ? _GEN6850 : _GEN9668;
wire  _GEN9670 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9671 = io_x[2] ? _GEN6837 : _GEN9670;
wire  _GEN9672 = io_x[6] ? _GEN6850 : _GEN9671;
wire  _GEN9673 = io_x[41] ? _GEN9672 : _GEN9669;
wire  _GEN9674 = io_x[14] ? _GEN6843 : _GEN9673;
wire  _GEN9675 = io_x[0] ? _GEN6845 : _GEN9674;
wire  _GEN9676 = io_x[76] ? _GEN9675 : _GEN9667;
wire  _GEN9677 = io_x[42] ? _GEN9676 : _GEN9665;
wire  _GEN9678 = io_x[38] ? _GEN9677 : _GEN9664;
wire  _GEN9679 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9680 = io_x[41] ? _GEN9679 : _GEN6836;
wire  _GEN9681 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9682 = io_x[6] ? _GEN6850 : _GEN9681;
wire  _GEN9683 = io_x[41] ? _GEN9682 : _GEN6836;
wire  _GEN9684 = io_x[14] ? _GEN9683 : _GEN9680;
wire  _GEN9685 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9686 = io_x[6] ? _GEN9685 : _GEN6850;
wire  _GEN9687 = io_x[41] ? _GEN9686 : _GEN6836;
wire  _GEN9688 = io_x[14] ? _GEN6856 : _GEN9687;
wire  _GEN9689 = io_x[0] ? _GEN9688 : _GEN9684;
wire  _GEN9690 = io_x[76] ? _GEN6834 : _GEN9689;
wire  _GEN9691 = io_x[42] ? _GEN9690 : _GEN6874;
wire  _GEN9692 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9693 = io_x[41] ? _GEN6836 : _GEN9692;
wire  _GEN9694 = io_x[14] ? _GEN9693 : _GEN6856;
wire  _GEN9695 = io_x[0] ? _GEN6858 : _GEN9694;
wire  _GEN9696 = io_x[76] ? _GEN6834 : _GEN9695;
wire  _GEN9697 = io_x[42] ? _GEN9696 : _GEN6863;
wire  _GEN9698 = io_x[38] ? _GEN9697 : _GEN9691;
wire  _GEN9699 = io_x[10] ? _GEN9698 : _GEN9678;
wire  _GEN9700 = io_x[71] ? _GEN9699 : _GEN9657;
wire  _GEN9701 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9702 = io_x[0] ? _GEN9701 : _GEN6858;
wire  _GEN9703 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9704 = io_x[6] ? _GEN6850 : _GEN9703;
wire  _GEN9705 = io_x[41] ? _GEN9704 : _GEN6836;
wire  _GEN9706 = io_x[14] ? _GEN6856 : _GEN9705;
wire  _GEN9707 = io_x[0] ? _GEN6845 : _GEN9706;
wire  _GEN9708 = io_x[76] ? _GEN9707 : _GEN9702;
wire  _GEN9709 = io_x[42] ? _GEN9708 : _GEN6874;
wire  _GEN9710 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN9711 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9712 = io_x[6] ? _GEN6840 : _GEN9711;
wire  _GEN9713 = io_x[41] ? _GEN6836 : _GEN9712;
wire  _GEN9714 = io_x[14] ? _GEN6843 : _GEN9713;
wire  _GEN9715 = io_x[0] ? _GEN6845 : _GEN9714;
wire  _GEN9716 = io_x[76] ? _GEN6834 : _GEN9715;
wire  _GEN9717 = io_x[42] ? _GEN9716 : _GEN9710;
wire  _GEN9718 = io_x[38] ? _GEN9717 : _GEN9709;
wire  _GEN9719 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9720 = io_x[41] ? _GEN9719 : _GEN6836;
wire  _GEN9721 = io_x[14] ? _GEN9720 : _GEN6843;
wire  _GEN9722 = io_x[0] ? _GEN6845 : _GEN9721;
wire  _GEN9723 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9724 = io_x[6] ? _GEN6850 : _GEN9723;
wire  _GEN9725 = io_x[41] ? _GEN6836 : _GEN9724;
wire  _GEN9726 = io_x[14] ? _GEN9725 : _GEN6843;
wire  _GEN9727 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9728 = io_x[0] ? _GEN9727 : _GEN9726;
wire  _GEN9729 = io_x[76] ? _GEN9728 : _GEN9722;
wire  _GEN9730 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9731 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN9732 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9733 = io_x[6] ? _GEN6850 : _GEN9732;
wire  _GEN9734 = io_x[41] ? _GEN6836 : _GEN9733;
wire  _GEN9735 = io_x[14] ? _GEN9734 : _GEN9731;
wire  _GEN9736 = io_x[0] ? _GEN9735 : _GEN9730;
wire  _GEN9737 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9738 = io_x[0] ? _GEN6845 : _GEN9737;
wire  _GEN9739 = io_x[76] ? _GEN9738 : _GEN9736;
wire  _GEN9740 = io_x[42] ? _GEN9739 : _GEN9729;
wire  _GEN9741 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9742 = io_x[0] ? _GEN9741 : _GEN6845;
wire  _GEN9743 = io_x[76] ? _GEN9742 : _GEN6834;
wire  _GEN9744 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9745 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9746 = io_x[6] ? _GEN9745 : _GEN9744;
wire  _GEN9747 = io_x[41] ? _GEN6836 : _GEN9746;
wire  _GEN9748 = io_x[14] ? _GEN9747 : _GEN6856;
wire  _GEN9749 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9750 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9751 = io_x[6] ? _GEN9750 : _GEN9749;
wire  _GEN9752 = io_x[41] ? _GEN6836 : _GEN9751;
wire  _GEN9753 = io_x[14] ? _GEN9752 : _GEN6856;
wire  _GEN9754 = io_x[0] ? _GEN9753 : _GEN9748;
wire  _GEN9755 = io_x[76] ? _GEN6834 : _GEN9754;
wire  _GEN9756 = io_x[42] ? _GEN9755 : _GEN9743;
wire  _GEN9757 = io_x[38] ? _GEN9756 : _GEN9740;
wire  _GEN9758 = io_x[10] ? _GEN9757 : _GEN9718;
wire  _GEN9759 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9760 = io_x[0] ? _GEN6845 : _GEN9759;
wire  _GEN9761 = io_x[76] ? _GEN6834 : _GEN9760;
wire  _GEN9762 = io_x[42] ? _GEN9761 : _GEN6874;
wire  _GEN9763 = io_x[38] ? _GEN9762 : _GEN6871;
wire  _GEN9764 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN9765 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN9766 = io_x[14] ? _GEN9765 : _GEN9764;
wire  _GEN9767 = io_x[0] ? _GEN6845 : _GEN9766;
wire  _GEN9768 = io_x[76] ? _GEN6834 : _GEN9767;
wire  _GEN9769 = io_x[42] ? _GEN6874 : _GEN9768;
wire  _GEN9770 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9771 = io_x[41] ? _GEN6836 : _GEN9770;
wire  _GEN9772 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9773 = io_x[41] ? _GEN6836 : _GEN9772;
wire  _GEN9774 = io_x[14] ? _GEN9773 : _GEN9771;
wire  _GEN9775 = io_x[0] ? _GEN9774 : _GEN6845;
wire  _GEN9776 = io_x[76] ? _GEN6834 : _GEN9775;
wire  _GEN9777 = io_x[42] ? _GEN9776 : _GEN6863;
wire  _GEN9778 = io_x[38] ? _GEN9777 : _GEN9769;
wire  _GEN9779 = io_x[10] ? _GEN9778 : _GEN9763;
wire  _GEN9780 = io_x[71] ? _GEN9779 : _GEN9758;
wire  _GEN9781 = io_x[70] ? _GEN9780 : _GEN9700;
wire  _GEN9782 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9783 = io_x[0] ? _GEN9782 : _GEN6845;
wire  _GEN9784 = io_x[76] ? _GEN6834 : _GEN9783;
wire  _GEN9785 = io_x[42] ? _GEN9784 : _GEN6874;
wire  _GEN9786 = io_x[38] ? _GEN9785 : _GEN6871;
wire  _GEN9787 = io_x[10] ? _GEN9786 : _GEN7044;
wire  _GEN9788 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9789 = io_x[6] ? _GEN6840 : _GEN9788;
wire  _GEN9790 = io_x[41] ? _GEN6836 : _GEN9789;
wire  _GEN9791 = io_x[14] ? _GEN6856 : _GEN9790;
wire  _GEN9792 = io_x[0] ? _GEN9791 : _GEN6845;
wire  _GEN9793 = io_x[76] ? _GEN6834 : _GEN9792;
wire  _GEN9794 = io_x[42] ? _GEN9793 : _GEN6874;
wire  _GEN9795 = io_x[38] ? _GEN9794 : _GEN6871;
wire  _GEN9796 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9797 = io_x[0] ? _GEN9796 : _GEN6845;
wire  _GEN9798 = io_x[76] ? _GEN6834 : _GEN9797;
wire  _GEN9799 = io_x[42] ? _GEN9798 : _GEN6874;
wire  _GEN9800 = io_x[38] ? _GEN9799 : _GEN6871;
wire  _GEN9801 = io_x[10] ? _GEN9800 : _GEN9795;
wire  _GEN9802 = io_x[71] ? _GEN9801 : _GEN9787;
wire  _GEN9803 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9804 = io_x[0] ? _GEN9803 : _GEN6845;
wire  _GEN9805 = io_x[76] ? _GEN9804 : _GEN6834;
wire  _GEN9806 = io_x[42] ? _GEN6874 : _GEN9805;
wire  _GEN9807 = io_x[38] ? _GEN9806 : _GEN7036;
wire  _GEN9808 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9809 = io_x[41] ? _GEN6836 : _GEN9808;
wire  _GEN9810 = io_x[14] ? _GEN9809 : _GEN6856;
wire  _GEN9811 = io_x[0] ? _GEN6845 : _GEN9810;
wire  _GEN9812 = io_x[76] ? _GEN6834 : _GEN9811;
wire  _GEN9813 = io_x[42] ? _GEN9812 : _GEN6874;
wire  _GEN9814 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9815 = io_x[41] ? _GEN9814 : _GEN6924;
wire  _GEN9816 = io_x[14] ? _GEN9815 : _GEN6843;
wire  _GEN9817 = io_x[0] ? _GEN9816 : _GEN6845;
wire  _GEN9818 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9819 = io_x[0] ? _GEN9818 : _GEN6845;
wire  _GEN9820 = io_x[76] ? _GEN9819 : _GEN9817;
wire  _GEN9821 = io_x[42] ? _GEN6874 : _GEN9820;
wire  _GEN9822 = io_x[38] ? _GEN9821 : _GEN9813;
wire  _GEN9823 = io_x[10] ? _GEN9822 : _GEN9807;
wire  _GEN9824 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9825 = io_x[41] ? _GEN6836 : _GEN9824;
wire  _GEN9826 = io_x[14] ? _GEN9825 : _GEN6856;
wire  _GEN9827 = io_x[0] ? _GEN9826 : _GEN6845;
wire  _GEN9828 = io_x[76] ? _GEN6834 : _GEN9827;
wire  _GEN9829 = io_x[42] ? _GEN9828 : _GEN6874;
wire  _GEN9830 = io_x[38] ? _GEN9829 : _GEN6871;
wire  _GEN9831 = io_x[10] ? _GEN9830 : _GEN7044;
wire  _GEN9832 = io_x[71] ? _GEN9831 : _GEN9823;
wire  _GEN9833 = io_x[70] ? _GEN9832 : _GEN9802;
wire  _GEN9834 = io_x[33] ? _GEN9833 : _GEN9781;
wire  _GEN9835 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9836 = io_x[0] ? _GEN9835 : _GEN6858;
wire  _GEN9837 = io_x[76] ? _GEN6834 : _GEN9836;
wire  _GEN9838 = io_x[42] ? _GEN9837 : _GEN6863;
wire  _GEN9839 = io_x[38] ? _GEN9838 : _GEN6871;
wire  _GEN9840 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9841 = io_x[41] ? _GEN9840 : _GEN6836;
wire  _GEN9842 = io_x[14] ? _GEN9841 : _GEN6843;
wire  _GEN9843 = io_x[0] ? _GEN9842 : _GEN6858;
wire  _GEN9844 = io_x[76] ? _GEN6834 : _GEN9843;
wire  _GEN9845 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN9846 = io_x[42] ? _GEN9845 : _GEN9844;
wire  _GEN9847 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN9848 = io_x[76] ? _GEN6833 : _GEN9847;
wire  _GEN9849 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9850 = io_x[6] ? _GEN9849 : _GEN6850;
wire  _GEN9851 = io_x[41] ? _GEN6924 : _GEN9850;
wire  _GEN9852 = io_x[14] ? _GEN9851 : _GEN6856;
wire  _GEN9853 = io_x[0] ? _GEN9852 : _GEN6845;
wire  _GEN9854 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9855 = io_x[41] ? _GEN9854 : _GEN6836;
wire  _GEN9856 = io_x[14] ? _GEN9855 : _GEN6843;
wire  _GEN9857 = io_x[0] ? _GEN6845 : _GEN9856;
wire  _GEN9858 = io_x[76] ? _GEN9857 : _GEN9853;
wire  _GEN9859 = io_x[42] ? _GEN9858 : _GEN9848;
wire  _GEN9860 = io_x[38] ? _GEN9859 : _GEN9846;
wire  _GEN9861 = io_x[10] ? _GEN9860 : _GEN9839;
wire  _GEN9862 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9863 = io_x[0] ? _GEN9862 : _GEN6845;
wire  _GEN9864 = io_x[76] ? _GEN6834 : _GEN9863;
wire  _GEN9865 = io_x[42] ? _GEN9864 : _GEN6874;
wire  _GEN9866 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN9867 = io_x[14] ? _GEN6843 : _GEN9866;
wire  _GEN9868 = io_x[0] ? _GEN6845 : _GEN9867;
wire  _GEN9869 = io_x[76] ? _GEN9868 : _GEN6833;
wire  _GEN9870 = io_x[42] ? _GEN9869 : _GEN6874;
wire  _GEN9871 = io_x[38] ? _GEN9870 : _GEN9865;
wire  _GEN9872 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9873 = io_x[6] ? _GEN9872 : _GEN6850;
wire  _GEN9874 = io_x[41] ? _GEN9873 : _GEN6836;
wire  _GEN9875 = io_x[14] ? _GEN9874 : _GEN6856;
wire  _GEN9876 = io_x[0] ? _GEN9875 : _GEN6858;
wire  _GEN9877 = io_x[76] ? _GEN6834 : _GEN9876;
wire  _GEN9878 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9879 = io_x[6] ? _GEN6850 : _GEN9878;
wire  _GEN9880 = io_x[41] ? _GEN9879 : _GEN6924;
wire  _GEN9881 = io_x[14] ? _GEN9880 : _GEN6843;
wire  _GEN9882 = io_x[0] ? _GEN9881 : _GEN6858;
wire  _GEN9883 = io_x[76] ? _GEN6834 : _GEN9882;
wire  _GEN9884 = io_x[42] ? _GEN9883 : _GEN9877;
wire  _GEN9885 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9886 = io_x[41] ? _GEN6836 : _GEN9885;
wire  _GEN9887 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9888 = io_x[41] ? _GEN6836 : _GEN9887;
wire  _GEN9889 = io_x[14] ? _GEN9888 : _GEN9886;
wire  _GEN9890 = io_x[0] ? _GEN9889 : _GEN6845;
wire  _GEN9891 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9892 = io_x[0] ? _GEN9891 : _GEN6845;
wire  _GEN9893 = io_x[76] ? _GEN9892 : _GEN9890;
wire  _GEN9894 = io_x[42] ? _GEN9893 : _GEN6863;
wire  _GEN9895 = io_x[38] ? _GEN9894 : _GEN9884;
wire  _GEN9896 = io_x[10] ? _GEN9895 : _GEN9871;
wire  _GEN9897 = io_x[71] ? _GEN9896 : _GEN9861;
wire  _GEN9898 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN9899 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9900 = io_x[41] ? _GEN6836 : _GEN9899;
wire  _GEN9901 = io_x[14] ? _GEN9900 : _GEN6843;
wire  _GEN9902 = io_x[0] ? _GEN6845 : _GEN9901;
wire  _GEN9903 = io_x[76] ? _GEN9902 : _GEN9898;
wire  _GEN9904 = io_x[42] ? _GEN9903 : _GEN6863;
wire  _GEN9905 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN9906 = io_x[76] ? _GEN6833 : _GEN9905;
wire  _GEN9907 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN9908 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9909 = io_x[2] ? _GEN6837 : _GEN9908;
wire  _GEN9910 = io_x[6] ? _GEN6850 : _GEN9909;
wire  _GEN9911 = io_x[41] ? _GEN9910 : _GEN6836;
wire  _GEN9912 = io_x[14] ? _GEN6843 : _GEN9911;
wire  _GEN9913 = io_x[0] ? _GEN6845 : _GEN9912;
wire  _GEN9914 = io_x[76] ? _GEN9913 : _GEN9907;
wire  _GEN9915 = io_x[42] ? _GEN9914 : _GEN9906;
wire  _GEN9916 = io_x[38] ? _GEN9915 : _GEN9904;
wire  _GEN9917 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9918 = io_x[41] ? _GEN9917 : _GEN6836;
wire  _GEN9919 = io_x[14] ? _GEN6856 : _GEN9918;
wire  _GEN9920 = io_x[0] ? _GEN9919 : _GEN6845;
wire  _GEN9921 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9922 = io_x[6] ? _GEN9921 : _GEN6850;
wire  _GEN9923 = io_x[41] ? _GEN6836 : _GEN9922;
wire  _GEN9924 = io_x[14] ? _GEN9923 : _GEN6856;
wire  _GEN9925 = io_x[0] ? _GEN6845 : _GEN9924;
wire  _GEN9926 = io_x[76] ? _GEN9925 : _GEN9920;
wire  _GEN9927 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9928 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9929 = io_x[6] ? _GEN9928 : _GEN6850;
wire  _GEN9930 = io_x[41] ? _GEN6836 : _GEN9929;
wire  _GEN9931 = io_x[14] ? _GEN9930 : _GEN6843;
wire  _GEN9932 = io_x[0] ? _GEN9931 : _GEN9927;
wire  _GEN9933 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9934 = io_x[41] ? _GEN9933 : _GEN6924;
wire  _GEN9935 = io_x[14] ? _GEN9934 : _GEN6856;
wire  _GEN9936 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9937 = io_x[2] ? _GEN6837 : _GEN9936;
wire  _GEN9938 = io_x[6] ? _GEN9937 : _GEN6850;
wire  _GEN9939 = io_x[41] ? _GEN9938 : _GEN6836;
wire  _GEN9940 = io_x[14] ? _GEN6856 : _GEN9939;
wire  _GEN9941 = io_x[0] ? _GEN9940 : _GEN9935;
wire  _GEN9942 = io_x[76] ? _GEN9941 : _GEN9932;
wire  _GEN9943 = io_x[42] ? _GEN9942 : _GEN9926;
wire  _GEN9944 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9945 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9946 = io_x[6] ? _GEN9945 : _GEN6850;
wire  _GEN9947 = io_x[41] ? _GEN6836 : _GEN9946;
wire  _GEN9948 = io_x[14] ? _GEN6856 : _GEN9947;
wire  _GEN9949 = io_x[0] ? _GEN9948 : _GEN9944;
wire  _GEN9950 = io_x[76] ? _GEN6833 : _GEN9949;
wire  _GEN9951 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN9952 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN9953 = io_x[6] ? _GEN9952 : _GEN6840;
wire  _GEN9954 = io_x[41] ? _GEN6836 : _GEN9953;
wire  _GEN9955 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9956 = io_x[6] ? _GEN9955 : _GEN6850;
wire  _GEN9957 = io_x[41] ? _GEN6836 : _GEN9956;
wire  _GEN9958 = io_x[14] ? _GEN9957 : _GEN9954;
wire  _GEN9959 = io_x[0] ? _GEN9958 : _GEN9951;
wire  _GEN9960 = io_x[76] ? _GEN6834 : _GEN9959;
wire  _GEN9961 = io_x[42] ? _GEN9960 : _GEN9950;
wire  _GEN9962 = io_x[38] ? _GEN9961 : _GEN9943;
wire  _GEN9963 = io_x[10] ? _GEN9962 : _GEN9916;
wire  _GEN9964 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN9965 = io_x[14] ? _GEN9964 : _GEN6843;
wire  _GEN9966 = io_x[0] ? _GEN6845 : _GEN9965;
wire  _GEN9967 = io_x[76] ? _GEN6834 : _GEN9966;
wire  _GEN9968 = io_x[42] ? _GEN6874 : _GEN9967;
wire  _GEN9969 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN9970 = io_x[2] ? _GEN6837 : _GEN9969;
wire  _GEN9971 = io_x[6] ? _GEN6850 : _GEN9970;
wire  _GEN9972 = io_x[41] ? _GEN9971 : _GEN6836;
wire  _GEN9973 = io_x[14] ? _GEN6843 : _GEN9972;
wire  _GEN9974 = io_x[0] ? _GEN6845 : _GEN9973;
wire  _GEN9975 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN9976 = io_x[14] ? _GEN6843 : _GEN9975;
wire  _GEN9977 = io_x[0] ? _GEN6845 : _GEN9976;
wire  _GEN9978 = io_x[76] ? _GEN9977 : _GEN9974;
wire  _GEN9979 = io_x[42] ? _GEN9978 : _GEN6863;
wire  _GEN9980 = io_x[38] ? _GEN9979 : _GEN9968;
wire  _GEN9981 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN9982 = io_x[6] ? _GEN9981 : _GEN6850;
wire  _GEN9983 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN9984 = io_x[41] ? _GEN9983 : _GEN9982;
wire  _GEN9985 = io_x[14] ? _GEN9984 : _GEN6843;
wire  _GEN9986 = io_x[0] ? _GEN9985 : _GEN6858;
wire  _GEN9987 = io_x[76] ? _GEN6834 : _GEN9986;
wire  _GEN9988 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9989 = io_x[41] ? _GEN9988 : _GEN6836;
wire  _GEN9990 = io_x[14] ? _GEN9989 : _GEN6843;
wire  _GEN9991 = io_x[0] ? _GEN6845 : _GEN9990;
wire  _GEN9992 = io_x[76] ? _GEN6834 : _GEN9991;
wire  _GEN9993 = io_x[42] ? _GEN9992 : _GEN9987;
wire  _GEN9994 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN9995 = io_x[76] ? _GEN6834 : _GEN9994;
wire  _GEN9996 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN9997 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN9998 = io_x[41] ? _GEN6836 : _GEN9997;
wire  _GEN9999 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10000 = io_x[41] ? _GEN6836 : _GEN9999;
wire  _GEN10001 = io_x[14] ? _GEN10000 : _GEN9998;
wire  _GEN10002 = io_x[0] ? _GEN10001 : _GEN9996;
wire  _GEN10003 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10004 = io_x[0] ? _GEN6845 : _GEN10003;
wire  _GEN10005 = io_x[76] ? _GEN10004 : _GEN10002;
wire  _GEN10006 = io_x[42] ? _GEN10005 : _GEN9995;
wire  _GEN10007 = io_x[38] ? _GEN10006 : _GEN9993;
wire  _GEN10008 = io_x[10] ? _GEN10007 : _GEN9980;
wire  _GEN10009 = io_x[71] ? _GEN10008 : _GEN9963;
wire  _GEN10010 = io_x[70] ? _GEN10009 : _GEN9897;
wire  _GEN10011 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10012 = io_x[41] ? _GEN10011 : _GEN6836;
wire  _GEN10013 = io_x[14] ? _GEN10012 : _GEN6843;
wire  _GEN10014 = io_x[0] ? _GEN10013 : _GEN6845;
wire  _GEN10015 = io_x[76] ? _GEN6834 : _GEN10014;
wire  _GEN10016 = io_x[42] ? _GEN6874 : _GEN10015;
wire  _GEN10017 = io_x[38] ? _GEN6871 : _GEN10016;
wire  _GEN10018 = io_x[10] ? _GEN10017 : _GEN7044;
wire  _GEN10019 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10020 = io_x[0] ? _GEN10019 : _GEN6845;
wire  _GEN10021 = io_x[76] ? _GEN6834 : _GEN10020;
wire  _GEN10022 = io_x[42] ? _GEN10021 : _GEN6863;
wire  _GEN10023 = io_x[38] ? _GEN10022 : _GEN6871;
wire  _GEN10024 = io_x[10] ? _GEN10023 : _GEN7044;
wire  _GEN10025 = io_x[71] ? _GEN10024 : _GEN10018;
wire  _GEN10026 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10027 = io_x[0] ? _GEN10026 : _GEN6845;
wire  _GEN10028 = io_x[76] ? _GEN6834 : _GEN10027;
wire  _GEN10029 = io_x[42] ? _GEN10028 : _GEN6863;
wire  _GEN10030 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10031 = io_x[41] ? _GEN10030 : _GEN6836;
wire  _GEN10032 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10033 = io_x[41] ? _GEN10032 : _GEN6924;
wire  _GEN10034 = io_x[14] ? _GEN10033 : _GEN10031;
wire  _GEN10035 = io_x[0] ? _GEN10034 : _GEN6845;
wire  _GEN10036 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10037 = io_x[0] ? _GEN10036 : _GEN6845;
wire  _GEN10038 = io_x[76] ? _GEN10037 : _GEN10035;
wire  _GEN10039 = io_x[42] ? _GEN6874 : _GEN10038;
wire  _GEN10040 = io_x[38] ? _GEN10039 : _GEN10029;
wire  _GEN10041 = io_x[10] ? _GEN10040 : _GEN7044;
wire  _GEN10042 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10043 = io_x[41] ? _GEN6836 : _GEN10042;
wire  _GEN10044 = io_x[14] ? _GEN6843 : _GEN10043;
wire  _GEN10045 = io_x[0] ? _GEN10044 : _GEN6845;
wire  _GEN10046 = io_x[76] ? _GEN6834 : _GEN10045;
wire  _GEN10047 = io_x[42] ? _GEN10046 : _GEN6863;
wire  _GEN10048 = io_x[38] ? _GEN10047 : _GEN6871;
wire  _GEN10049 = io_x[10] ? _GEN10048 : _GEN7044;
wire  _GEN10050 = io_x[71] ? _GEN10049 : _GEN10041;
wire  _GEN10051 = io_x[70] ? _GEN10050 : _GEN10025;
wire  _GEN10052 = io_x[33] ? _GEN10051 : _GEN10010;
wire  _GEN10053 = io_x[21] ? _GEN10052 : _GEN9834;
wire  _GEN10054 = io_x[18] ? _GEN10053 : _GEN9647;
wire  _GEN10055 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10056 = io_x[0] ? _GEN6845 : _GEN10055;
wire  _GEN10057 = io_x[76] ? _GEN6834 : _GEN10056;
wire  _GEN10058 = io_x[42] ? _GEN10057 : _GEN6874;
wire  _GEN10059 = io_x[38] ? _GEN10058 : _GEN7036;
wire  _GEN10060 = io_x[10] ? _GEN10059 : _GEN7044;
wire  _GEN10061 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10062 = io_x[0] ? _GEN6845 : _GEN10061;
wire  _GEN10063 = io_x[76] ? _GEN10062 : _GEN6833;
wire  _GEN10064 = io_x[42] ? _GEN10063 : _GEN6874;
wire  _GEN10065 = io_x[38] ? _GEN10064 : _GEN7036;
wire  _GEN10066 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10067 = io_x[0] ? _GEN6845 : _GEN10066;
wire  _GEN10068 = io_x[76] ? _GEN6834 : _GEN10067;
wire  _GEN10069 = io_x[42] ? _GEN10068 : _GEN6874;
wire  _GEN10070 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10071 = io_x[0] ? _GEN10070 : _GEN6845;
wire  _GEN10072 = io_x[76] ? _GEN10071 : _GEN6834;
wire  _GEN10073 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10074 = io_x[0] ? _GEN6845 : _GEN10073;
wire  _GEN10075 = io_x[76] ? _GEN10074 : _GEN6834;
wire  _GEN10076 = io_x[42] ? _GEN10075 : _GEN10072;
wire  _GEN10077 = io_x[38] ? _GEN10076 : _GEN10069;
wire  _GEN10078 = io_x[10] ? _GEN10077 : _GEN10065;
wire  _GEN10079 = io_x[71] ? _GEN10078 : _GEN10060;
wire  _GEN10080 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN10081 = io_x[42] ? _GEN10080 : _GEN6874;
wire  _GEN10082 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN10083 = io_x[42] ? _GEN6874 : _GEN10082;
wire  _GEN10084 = io_x[38] ? _GEN10083 : _GEN10081;
wire  _GEN10085 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN10086 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10087 = io_x[6] ? _GEN6840 : _GEN10086;
wire  _GEN10088 = io_x[41] ? _GEN6836 : _GEN10087;
wire  _GEN10089 = io_x[14] ? _GEN10088 : _GEN6843;
wire  _GEN10090 = io_x[0] ? _GEN10089 : _GEN6845;
wire  _GEN10091 = io_x[76] ? _GEN6833 : _GEN10090;
wire  _GEN10092 = io_x[42] ? _GEN10091 : _GEN10085;
wire  _GEN10093 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10094 = io_x[0] ? _GEN6845 : _GEN10093;
wire  _GEN10095 = io_x[76] ? _GEN6834 : _GEN10094;
wire  _GEN10096 = io_x[42] ? _GEN10095 : _GEN6874;
wire  _GEN10097 = io_x[38] ? _GEN10096 : _GEN10092;
wire  _GEN10098 = io_x[10] ? _GEN10097 : _GEN10084;
wire  _GEN10099 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10100 = io_x[6] ? _GEN6850 : _GEN10099;
wire  _GEN10101 = io_x[41] ? _GEN10100 : _GEN6836;
wire  _GEN10102 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10103 = io_x[41] ? _GEN10102 : _GEN6836;
wire  _GEN10104 = io_x[14] ? _GEN10103 : _GEN10101;
wire  _GEN10105 = io_x[0] ? _GEN6845 : _GEN10104;
wire  _GEN10106 = io_x[76] ? _GEN6833 : _GEN10105;
wire  _GEN10107 = io_x[42] ? _GEN6863 : _GEN10106;
wire  _GEN10108 = io_x[38] ? _GEN6871 : _GEN10107;
wire  _GEN10109 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10110 = io_x[6] ? _GEN10109 : _GEN6850;
wire  _GEN10111 = io_x[41] ? _GEN10110 : _GEN6836;
wire  _GEN10112 = io_x[14] ? _GEN10111 : _GEN6843;
wire  _GEN10113 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10114 = io_x[0] ? _GEN10113 : _GEN10112;
wire  _GEN10115 = io_x[76] ? _GEN6834 : _GEN10114;
wire  _GEN10116 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10117 = io_x[0] ? _GEN10116 : _GEN6845;
wire  _GEN10118 = io_x[76] ? _GEN6834 : _GEN10117;
wire  _GEN10119 = io_x[42] ? _GEN10118 : _GEN10115;
wire  _GEN10120 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10121 = io_x[41] ? _GEN10120 : _GEN6836;
wire  _GEN10122 = io_x[14] ? _GEN10121 : _GEN6843;
wire  _GEN10123 = io_x[0] ? _GEN6845 : _GEN10122;
wire  _GEN10124 = io_x[76] ? _GEN6834 : _GEN10123;
wire  _GEN10125 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10126 = io_x[41] ? _GEN6836 : _GEN10125;
wire  _GEN10127 = io_x[14] ? _GEN10126 : _GEN6843;
wire  _GEN10128 = io_x[0] ? _GEN6858 : _GEN10127;
wire  _GEN10129 = io_x[76] ? _GEN6834 : _GEN10128;
wire  _GEN10130 = io_x[42] ? _GEN10129 : _GEN10124;
wire  _GEN10131 = io_x[38] ? _GEN10130 : _GEN10119;
wire  _GEN10132 = io_x[10] ? _GEN10131 : _GEN10108;
wire  _GEN10133 = io_x[71] ? _GEN10132 : _GEN10098;
wire  _GEN10134 = io_x[70] ? _GEN10133 : _GEN10079;
wire  _GEN10135 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10136 = io_x[0] ? _GEN10135 : _GEN6845;
wire  _GEN10137 = io_x[76] ? _GEN10136 : _GEN6834;
wire  _GEN10138 = io_x[42] ? _GEN6874 : _GEN10137;
wire  _GEN10139 = io_x[38] ? _GEN10138 : _GEN6871;
wire  _GEN10140 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10141 = io_x[0] ? _GEN10140 : _GEN6845;
wire  _GEN10142 = io_x[76] ? _GEN10141 : _GEN6834;
wire  _GEN10143 = io_x[42] ? _GEN6874 : _GEN10142;
wire  _GEN10144 = io_x[38] ? _GEN10143 : _GEN6871;
wire  _GEN10145 = io_x[10] ? _GEN10144 : _GEN10139;
wire  _GEN10146 = io_x[71] ? _GEN10145 : _GEN7196;
wire  _GEN10147 = io_x[70] ? _GEN8474 : _GEN10146;
wire  _GEN10148 = io_x[33] ? _GEN10147 : _GEN10134;
wire  _GEN10149 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN10150 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10151 = io_x[6] ? _GEN6850 : _GEN10150;
wire  _GEN10152 = io_x[41] ? _GEN10151 : _GEN6836;
wire  _GEN10153 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10154 = io_x[41] ? _GEN10153 : _GEN6836;
wire  _GEN10155 = io_x[14] ? _GEN10154 : _GEN10152;
wire  _GEN10156 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10157 = io_x[6] ? _GEN6840 : _GEN10156;
wire  _GEN10158 = io_x[41] ? _GEN10157 : _GEN6924;
wire  _GEN10159 = io_x[14] ? _GEN10158 : _GEN6843;
wire  _GEN10160 = io_x[0] ? _GEN10159 : _GEN10155;
wire  _GEN10161 = io_x[76] ? _GEN6834 : _GEN10160;
wire  _GEN10162 = io_x[42] ? _GEN10161 : _GEN10149;
wire  _GEN10163 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN10164 = io_x[42] ? _GEN6863 : _GEN10163;
wire  _GEN10165 = io_x[38] ? _GEN10164 : _GEN10162;
wire  _GEN10166 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10167 = io_x[6] ? _GEN10166 : _GEN6850;
wire  _GEN10168 = io_x[41] ? _GEN10167 : _GEN6836;
wire  _GEN10169 = io_x[14] ? _GEN10168 : _GEN6843;
wire  _GEN10170 = io_x[0] ? _GEN10169 : _GEN6858;
wire  _GEN10171 = io_x[76] ? _GEN6833 : _GEN10170;
wire  _GEN10172 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10173 = io_x[41] ? _GEN10172 : _GEN6836;
wire  _GEN10174 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10175 = io_x[6] ? _GEN6850 : _GEN10174;
wire  _GEN10176 = io_x[41] ? _GEN10175 : _GEN6924;
wire  _GEN10177 = io_x[14] ? _GEN10176 : _GEN10173;
wire  _GEN10178 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10179 = io_x[0] ? _GEN10178 : _GEN10177;
wire  _GEN10180 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10181 = io_x[0] ? _GEN6845 : _GEN10180;
wire  _GEN10182 = io_x[76] ? _GEN10181 : _GEN10179;
wire  _GEN10183 = io_x[42] ? _GEN10182 : _GEN10171;
wire  _GEN10184 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10185 = io_x[41] ? _GEN10184 : _GEN6836;
wire  _GEN10186 = io_x[14] ? _GEN10185 : _GEN6843;
wire  _GEN10187 = io_x[0] ? _GEN6845 : _GEN10186;
wire  _GEN10188 = io_x[76] ? _GEN6833 : _GEN10187;
wire  _GEN10189 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10190 = io_x[6] ? _GEN10189 : _GEN6850;
wire  _GEN10191 = io_x[41] ? _GEN6836 : _GEN10190;
wire  _GEN10192 = io_x[14] ? _GEN10191 : _GEN6843;
wire  _GEN10193 = io_x[0] ? _GEN10192 : _GEN6845;
wire  _GEN10194 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10195 = io_x[2] ? _GEN10194 : _GEN6837;
wire  _GEN10196 = io_x[6] ? _GEN10195 : _GEN6850;
wire  _GEN10197 = io_x[41] ? _GEN6836 : _GEN10196;
wire  _GEN10198 = io_x[14] ? _GEN10197 : _GEN6856;
wire  _GEN10199 = io_x[0] ? _GEN10198 : _GEN6845;
wire  _GEN10200 = io_x[76] ? _GEN10199 : _GEN10193;
wire  _GEN10201 = io_x[42] ? _GEN10200 : _GEN10188;
wire  _GEN10202 = io_x[38] ? _GEN10201 : _GEN10183;
wire  _GEN10203 = io_x[10] ? _GEN10202 : _GEN10165;
wire  _GEN10204 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN10205 = io_x[76] ? _GEN6834 : _GEN10204;
wire  _GEN10206 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10207 = io_x[0] ? _GEN10206 : _GEN6845;
wire  _GEN10208 = io_x[76] ? _GEN6833 : _GEN10207;
wire  _GEN10209 = io_x[42] ? _GEN10208 : _GEN10205;
wire  _GEN10210 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10211 = io_x[6] ? _GEN10210 : _GEN6850;
wire  _GEN10212 = io_x[41] ? _GEN6836 : _GEN10211;
wire  _GEN10213 = io_x[14] ? _GEN10212 : _GEN6843;
wire  _GEN10214 = io_x[0] ? _GEN6845 : _GEN10213;
wire  _GEN10215 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10216 = io_x[6] ? _GEN6850 : _GEN10215;
wire  _GEN10217 = io_x[41] ? _GEN6836 : _GEN10216;
wire  _GEN10218 = io_x[14] ? _GEN6843 : _GEN10217;
wire  _GEN10219 = io_x[0] ? _GEN10218 : _GEN6845;
wire  _GEN10220 = io_x[76] ? _GEN10219 : _GEN10214;
wire  _GEN10221 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10222 = io_x[2] ? _GEN6837 : _GEN10221;
wire  _GEN10223 = io_x[6] ? _GEN6850 : _GEN10222;
wire  _GEN10224 = io_x[41] ? _GEN10223 : _GEN6836;
wire  _GEN10225 = io_x[14] ? _GEN6843 : _GEN10224;
wire  _GEN10226 = io_x[0] ? _GEN6845 : _GEN10225;
wire  _GEN10227 = io_x[76] ? _GEN10226 : _GEN6833;
wire  _GEN10228 = io_x[42] ? _GEN10227 : _GEN10220;
wire  _GEN10229 = io_x[38] ? _GEN10228 : _GEN10209;
wire  _GEN10230 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10231 = io_x[6] ? _GEN10230 : _GEN6850;
wire  _GEN10232 = io_x[41] ? _GEN10231 : _GEN6836;
wire  _GEN10233 = io_x[14] ? _GEN10232 : _GEN6843;
wire  _GEN10234 = io_x[0] ? _GEN10233 : _GEN6858;
wire  _GEN10235 = io_x[76] ? _GEN6834 : _GEN10234;
wire  _GEN10236 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10237 = io_x[6] ? _GEN10236 : _GEN6840;
wire  _GEN10238 = io_x[41] ? _GEN10237 : _GEN6836;
wire  _GEN10239 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10240 = io_x[6] ? _GEN10239 : _GEN6850;
wire  _GEN10241 = io_x[41] ? _GEN10240 : _GEN6836;
wire  _GEN10242 = io_x[14] ? _GEN10241 : _GEN10238;
wire  _GEN10243 = io_x[0] ? _GEN10242 : _GEN6845;
wire  _GEN10244 = io_x[76] ? _GEN6834 : _GEN10243;
wire  _GEN10245 = io_x[42] ? _GEN10244 : _GEN10235;
wire  _GEN10246 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10247 = io_x[0] ? _GEN10246 : _GEN6858;
wire  _GEN10248 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10249 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10250 = io_x[6] ? _GEN10249 : _GEN10248;
wire  _GEN10251 = io_x[41] ? _GEN6836 : _GEN10250;
wire  _GEN10252 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10253 = io_x[6] ? _GEN10252 : _GEN6850;
wire  _GEN10254 = io_x[41] ? _GEN6836 : _GEN10253;
wire  _GEN10255 = io_x[14] ? _GEN10254 : _GEN10251;
wire  _GEN10256 = io_x[0] ? _GEN10255 : _GEN6845;
wire  _GEN10257 = io_x[76] ? _GEN10256 : _GEN10247;
wire  _GEN10258 = io_x[42] ? _GEN6874 : _GEN10257;
wire  _GEN10259 = io_x[38] ? _GEN10258 : _GEN10245;
wire  _GEN10260 = io_x[10] ? _GEN10259 : _GEN10229;
wire  _GEN10261 = io_x[71] ? _GEN10260 : _GEN10203;
wire  _GEN10262 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10263 = io_x[2] ? _GEN6837 : _GEN10262;
wire  _GEN10264 = io_x[6] ? _GEN6840 : _GEN10263;
wire  _GEN10265 = io_x[41] ? _GEN10264 : _GEN6836;
wire  _GEN10266 = io_x[14] ? _GEN6843 : _GEN10265;
wire  _GEN10267 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10268 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10269 = io_x[6] ? _GEN10268 : _GEN10267;
wire  _GEN10270 = io_x[41] ? _GEN6836 : _GEN10269;
wire  _GEN10271 = io_x[14] ? _GEN10270 : _GEN6843;
wire  _GEN10272 = io_x[0] ? _GEN10271 : _GEN10266;
wire  _GEN10273 = io_x[76] ? _GEN6834 : _GEN10272;
wire  _GEN10274 = io_x[42] ? _GEN10273 : _GEN6874;
wire  _GEN10275 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10276 = io_x[0] ? _GEN6845 : _GEN10275;
wire  _GEN10277 = io_x[76] ? _GEN6834 : _GEN10276;
wire  _GEN10278 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10279 = io_x[41] ? _GEN6836 : _GEN10278;
wire  _GEN10280 = io_x[14] ? _GEN10279 : _GEN6843;
wire  _GEN10281 = io_x[0] ? _GEN10280 : _GEN6858;
wire  _GEN10282 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10283 = io_x[2] ? _GEN6837 : _GEN10282;
wire  _GEN10284 = io_x[6] ? _GEN6850 : _GEN10283;
wire  _GEN10285 = io_x[41] ? _GEN10284 : _GEN6836;
wire  _GEN10286 = io_x[14] ? _GEN6843 : _GEN10285;
wire  _GEN10287 = io_x[0] ? _GEN6845 : _GEN10286;
wire  _GEN10288 = io_x[76] ? _GEN10287 : _GEN10281;
wire  _GEN10289 = io_x[42] ? _GEN10288 : _GEN10277;
wire  _GEN10290 = io_x[38] ? _GEN10289 : _GEN10274;
wire  _GEN10291 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10292 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10293 = io_x[6] ? _GEN10292 : _GEN10291;
wire  _GEN10294 = io_x[41] ? _GEN10293 : _GEN6836;
wire  _GEN10295 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10296 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10297 = io_x[6] ? _GEN10296 : _GEN10295;
wire  _GEN10298 = io_x[41] ? _GEN10297 : _GEN6836;
wire  _GEN10299 = io_x[14] ? _GEN10298 : _GEN10294;
wire  _GEN10300 = io_x[0] ? _GEN6845 : _GEN10299;
wire  _GEN10301 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10302 = io_x[6] ? _GEN10301 : _GEN6840;
wire  _GEN10303 = io_x[41] ? _GEN6836 : _GEN10302;
wire  _GEN10304 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10305 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10306 = io_x[6] ? _GEN10305 : _GEN10304;
wire  _GEN10307 = io_x[41] ? _GEN6836 : _GEN10306;
wire  _GEN10308 = io_x[14] ? _GEN10307 : _GEN10303;
wire  _GEN10309 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10310 = io_x[41] ? _GEN6836 : _GEN10309;
wire  _GEN10311 = io_x[14] ? _GEN10310 : _GEN6856;
wire  _GEN10312 = io_x[0] ? _GEN10311 : _GEN10308;
wire  _GEN10313 = io_x[76] ? _GEN10312 : _GEN10300;
wire  _GEN10314 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10315 = io_x[41] ? _GEN6836 : _GEN10314;
wire  _GEN10316 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10317 = io_x[6] ? _GEN10316 : _GEN6850;
wire  _GEN10318 = io_x[41] ? _GEN6836 : _GEN10317;
wire  _GEN10319 = io_x[14] ? _GEN10318 : _GEN10315;
wire  _GEN10320 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10321 = io_x[6] ? _GEN10320 : _GEN6840;
wire  _GEN10322 = io_x[41] ? _GEN10321 : _GEN6836;
wire  _GEN10323 = io_x[14] ? _GEN6856 : _GEN10322;
wire  _GEN10324 = io_x[0] ? _GEN10323 : _GEN10319;
wire  _GEN10325 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10326 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN10327 = io_x[14] ? _GEN10326 : _GEN6843;
wire  _GEN10328 = io_x[0] ? _GEN10327 : _GEN10325;
wire  _GEN10329 = io_x[76] ? _GEN10328 : _GEN10324;
wire  _GEN10330 = io_x[42] ? _GEN10329 : _GEN10313;
wire  _GEN10331 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10332 = io_x[6] ? _GEN10331 : _GEN6840;
wire  _GEN10333 = io_x[41] ? _GEN10332 : _GEN6924;
wire  _GEN10334 = io_x[14] ? _GEN10333 : _GEN6843;
wire  _GEN10335 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10336 = io_x[0] ? _GEN10335 : _GEN10334;
wire  _GEN10337 = io_x[76] ? _GEN6833 : _GEN10336;
wire  _GEN10338 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10339 = io_x[41] ? _GEN6836 : _GEN10338;
wire  _GEN10340 = io_x[14] ? _GEN10339 : _GEN6843;
wire  _GEN10341 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10342 = io_x[41] ? _GEN6836 : _GEN10341;
wire  _GEN10343 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10344 = io_x[41] ? _GEN6836 : _GEN10343;
wire  _GEN10345 = io_x[14] ? _GEN10344 : _GEN10342;
wire  _GEN10346 = io_x[0] ? _GEN10345 : _GEN10340;
wire  _GEN10347 = io_x[76] ? _GEN6834 : _GEN10346;
wire  _GEN10348 = io_x[42] ? _GEN10347 : _GEN10337;
wire  _GEN10349 = io_x[38] ? _GEN10348 : _GEN10330;
wire  _GEN10350 = io_x[10] ? _GEN10349 : _GEN10290;
wire  _GEN10351 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN10352 = io_x[76] ? _GEN6834 : _GEN10351;
wire  _GEN10353 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN10354 = io_x[42] ? _GEN10353 : _GEN10352;
wire  _GEN10355 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10356 = io_x[2] ? _GEN6837 : _GEN10355;
wire  _GEN10357 = io_x[6] ? _GEN6850 : _GEN10356;
wire  _GEN10358 = io_x[41] ? _GEN10357 : _GEN6836;
wire  _GEN10359 = io_x[14] ? _GEN6843 : _GEN10358;
wire  _GEN10360 = io_x[0] ? _GEN6845 : _GEN10359;
wire  _GEN10361 = io_x[76] ? _GEN6834 : _GEN10360;
wire  _GEN10362 = io_x[42] ? _GEN10361 : _GEN6863;
wire  _GEN10363 = io_x[38] ? _GEN10362 : _GEN10354;
wire  _GEN10364 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10365 = io_x[41] ? _GEN10364 : _GEN6836;
wire  _GEN10366 = io_x[14] ? _GEN6856 : _GEN10365;
wire  _GEN10367 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10368 = io_x[6] ? _GEN10367 : _GEN6850;
wire  _GEN10369 = io_x[41] ? _GEN10368 : _GEN6924;
wire  _GEN10370 = io_x[14] ? _GEN10369 : _GEN6856;
wire  _GEN10371 = io_x[0] ? _GEN10370 : _GEN10366;
wire  _GEN10372 = io_x[76] ? _GEN6834 : _GEN10371;
wire  _GEN10373 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN10374 = io_x[76] ? _GEN10373 : _GEN6833;
wire  _GEN10375 = io_x[42] ? _GEN10374 : _GEN10372;
wire  _GEN10376 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN10377 = io_x[76] ? _GEN6833 : _GEN10376;
wire  _GEN10378 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10379 = io_x[41] ? _GEN6836 : _GEN10378;
wire  _GEN10380 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10381 = io_x[41] ? _GEN6836 : _GEN10380;
wire  _GEN10382 = io_x[14] ? _GEN10381 : _GEN10379;
wire  _GEN10383 = io_x[0] ? _GEN6858 : _GEN10382;
wire  _GEN10384 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10385 = io_x[0] ? _GEN6845 : _GEN10384;
wire  _GEN10386 = io_x[76] ? _GEN10385 : _GEN10383;
wire  _GEN10387 = io_x[42] ? _GEN10386 : _GEN10377;
wire  _GEN10388 = io_x[38] ? _GEN10387 : _GEN10375;
wire  _GEN10389 = io_x[10] ? _GEN10388 : _GEN10363;
wire  _GEN10390 = io_x[71] ? _GEN10389 : _GEN10350;
wire  _GEN10391 = io_x[70] ? _GEN10390 : _GEN10261;
wire  _GEN10392 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10393 = io_x[0] ? _GEN10392 : _GEN6845;
wire  _GEN10394 = io_x[76] ? _GEN10393 : _GEN6834;
wire  _GEN10395 = io_x[42] ? _GEN6874 : _GEN10394;
wire  _GEN10396 = io_x[38] ? _GEN10395 : _GEN6871;
wire  _GEN10397 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10398 = io_x[6] ? _GEN10397 : _GEN6850;
wire  _GEN10399 = io_x[41] ? _GEN6836 : _GEN10398;
wire  _GEN10400 = io_x[14] ? _GEN10399 : _GEN6843;
wire  _GEN10401 = io_x[0] ? _GEN10400 : _GEN6845;
wire  _GEN10402 = io_x[76] ? _GEN10401 : _GEN6834;
wire  _GEN10403 = io_x[42] ? _GEN6874 : _GEN10402;
wire  _GEN10404 = io_x[38] ? _GEN10403 : _GEN7036;
wire  _GEN10405 = io_x[10] ? _GEN10404 : _GEN10396;
wire  _GEN10406 = io_x[71] ? _GEN10405 : _GEN7196;
wire  _GEN10407 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10408 = io_x[0] ? _GEN10407 : _GEN6845;
wire  _GEN10409 = io_x[76] ? _GEN6833 : _GEN10408;
wire  _GEN10410 = io_x[42] ? _GEN6874 : _GEN10409;
wire  _GEN10411 = io_x[38] ? _GEN10410 : _GEN6871;
wire  _GEN10412 = io_x[10] ? _GEN10411 : _GEN7044;
wire  _GEN10413 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN10414 = io_x[38] ? _GEN6871 : _GEN10413;
wire  _GEN10415 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10416 = io_x[41] ? _GEN6836 : _GEN10415;
wire  _GEN10417 = io_x[14] ? _GEN10416 : _GEN6856;
wire  _GEN10418 = io_x[0] ? _GEN6845 : _GEN10417;
wire  _GEN10419 = io_x[76] ? _GEN6834 : _GEN10418;
wire  _GEN10420 = io_x[42] ? _GEN10419 : _GEN6874;
wire  _GEN10421 = io_x[38] ? _GEN10420 : _GEN6871;
wire  _GEN10422 = io_x[10] ? _GEN10421 : _GEN10414;
wire  _GEN10423 = io_x[71] ? _GEN10422 : _GEN10412;
wire  _GEN10424 = io_x[70] ? _GEN10423 : _GEN10406;
wire  _GEN10425 = io_x[33] ? _GEN10424 : _GEN10391;
wire  _GEN10426 = io_x[21] ? _GEN10425 : _GEN10148;
wire  _GEN10427 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN10428 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10429 = io_x[0] ? _GEN6845 : _GEN10428;
wire  _GEN10430 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10431 = io_x[0] ? _GEN6845 : _GEN10430;
wire  _GEN10432 = io_x[76] ? _GEN10431 : _GEN10429;
wire  _GEN10433 = io_x[42] ? _GEN10432 : _GEN10427;
wire  _GEN10434 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN10435 = io_x[14] ? _GEN10434 : _GEN6843;
wire  _GEN10436 = io_x[0] ? _GEN10435 : _GEN6845;
wire  _GEN10437 = io_x[76] ? _GEN10436 : _GEN6834;
wire  _GEN10438 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10439 = io_x[6] ? _GEN6850 : _GEN10438;
wire  _GEN10440 = io_x[41] ? _GEN6836 : _GEN10439;
wire  _GEN10441 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10442 = io_x[6] ? _GEN10441 : _GEN6850;
wire  _GEN10443 = io_x[41] ? _GEN6836 : _GEN10442;
wire  _GEN10444 = io_x[14] ? _GEN10443 : _GEN10440;
wire  _GEN10445 = io_x[0] ? _GEN10444 : _GEN6858;
wire  _GEN10446 = io_x[76] ? _GEN6834 : _GEN10445;
wire  _GEN10447 = io_x[42] ? _GEN10446 : _GEN10437;
wire  _GEN10448 = io_x[38] ? _GEN10447 : _GEN10433;
wire  _GEN10449 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN10450 = io_x[76] ? _GEN6834 : _GEN10449;
wire  _GEN10451 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10452 = io_x[6] ? _GEN10451 : _GEN6840;
wire  _GEN10453 = io_x[41] ? _GEN10452 : _GEN6836;
wire  _GEN10454 = io_x[14] ? _GEN10453 : _GEN6856;
wire  _GEN10455 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10456 = io_x[6] ? _GEN10455 : _GEN6850;
wire  _GEN10457 = io_x[41] ? _GEN6836 : _GEN10456;
wire  _GEN10458 = io_x[14] ? _GEN10457 : _GEN6843;
wire  _GEN10459 = io_x[0] ? _GEN10458 : _GEN10454;
wire  _GEN10460 = io_x[76] ? _GEN6834 : _GEN10459;
wire  _GEN10461 = io_x[42] ? _GEN10460 : _GEN10450;
wire  _GEN10462 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10463 = io_x[0] ? _GEN10462 : _GEN6845;
wire  _GEN10464 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10465 = io_x[41] ? _GEN6836 : _GEN10464;
wire  _GEN10466 = io_x[14] ? _GEN10465 : _GEN6856;
wire  _GEN10467 = io_x[0] ? _GEN10466 : _GEN6845;
wire  _GEN10468 = io_x[76] ? _GEN10467 : _GEN10463;
wire  _GEN10469 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10470 = io_x[41] ? _GEN6836 : _GEN10469;
wire  _GEN10471 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10472 = io_x[41] ? _GEN6924 : _GEN10471;
wire  _GEN10473 = io_x[14] ? _GEN10472 : _GEN10470;
wire  _GEN10474 = io_x[0] ? _GEN10473 : _GEN6858;
wire  _GEN10475 = io_x[76] ? _GEN6834 : _GEN10474;
wire  _GEN10476 = io_x[42] ? _GEN10475 : _GEN10468;
wire  _GEN10477 = io_x[38] ? _GEN10476 : _GEN10461;
wire  _GEN10478 = io_x[10] ? _GEN10477 : _GEN10448;
wire  _GEN10479 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN10480 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10481 = io_x[2] ? _GEN6837 : _GEN10480;
wire  _GEN10482 = io_x[6] ? _GEN6840 : _GEN10481;
wire  _GEN10483 = io_x[41] ? _GEN10482 : _GEN6836;
wire  _GEN10484 = io_x[14] ? _GEN6843 : _GEN10483;
wire  _GEN10485 = io_x[0] ? _GEN6845 : _GEN10484;
wire  _GEN10486 = io_x[76] ? _GEN10485 : _GEN6833;
wire  _GEN10487 = io_x[42] ? _GEN10486 : _GEN6863;
wire  _GEN10488 = io_x[38] ? _GEN10487 : _GEN10479;
wire  _GEN10489 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10490 = io_x[0] ? _GEN10489 : _GEN6858;
wire  _GEN10491 = io_x[76] ? _GEN6834 : _GEN10490;
wire  _GEN10492 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10493 = io_x[0] ? _GEN10492 : _GEN6845;
wire  _GEN10494 = io_x[76] ? _GEN10493 : _GEN6833;
wire  _GEN10495 = io_x[42] ? _GEN10494 : _GEN10491;
wire  _GEN10496 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN10497 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10498 = io_x[2] ? _GEN10497 : _GEN6838;
wire  _GEN10499 = io_x[6] ? _GEN10498 : _GEN6840;
wire  _GEN10500 = io_x[41] ? _GEN6836 : _GEN10499;
wire  _GEN10501 = io_x[14] ? _GEN10500 : _GEN10496;
wire  _GEN10502 = io_x[0] ? _GEN10501 : _GEN6858;
wire  _GEN10503 = io_x[76] ? _GEN6834 : _GEN10502;
wire  _GEN10504 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10505 = io_x[0] ? _GEN10504 : _GEN6845;
wire  _GEN10506 = io_x[76] ? _GEN6834 : _GEN10505;
wire  _GEN10507 = io_x[42] ? _GEN10506 : _GEN10503;
wire  _GEN10508 = io_x[38] ? _GEN10507 : _GEN10495;
wire  _GEN10509 = io_x[10] ? _GEN10508 : _GEN10488;
wire  _GEN10510 = io_x[71] ? _GEN10509 : _GEN10478;
wire  _GEN10511 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN10512 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10513 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10514 = io_x[41] ? _GEN6836 : _GEN10513;
wire  _GEN10515 = io_x[14] ? _GEN10514 : _GEN6843;
wire  _GEN10516 = io_x[0] ? _GEN10515 : _GEN10512;
wire  _GEN10517 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10518 = io_x[0] ? _GEN6845 : _GEN10517;
wire  _GEN10519 = io_x[76] ? _GEN10518 : _GEN10516;
wire  _GEN10520 = io_x[42] ? _GEN10519 : _GEN10511;
wire  _GEN10521 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10522 = io_x[0] ? _GEN6845 : _GEN10521;
wire  _GEN10523 = io_x[76] ? _GEN6834 : _GEN10522;
wire  _GEN10524 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10525 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10526 = io_x[6] ? _GEN10525 : _GEN10524;
wire  _GEN10527 = io_x[41] ? _GEN6836 : _GEN10526;
wire  _GEN10528 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10529 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10530 = io_x[6] ? _GEN10529 : _GEN10528;
wire  _GEN10531 = io_x[41] ? _GEN6836 : _GEN10530;
wire  _GEN10532 = io_x[14] ? _GEN10531 : _GEN10527;
wire  _GEN10533 = io_x[0] ? _GEN6845 : _GEN10532;
wire  _GEN10534 = io_x[76] ? _GEN6834 : _GEN10533;
wire  _GEN10535 = io_x[42] ? _GEN10534 : _GEN10523;
wire  _GEN10536 = io_x[38] ? _GEN10535 : _GEN10520;
wire  _GEN10537 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10538 = io_x[0] ? _GEN10537 : _GEN6845;
wire  _GEN10539 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10540 = io_x[41] ? _GEN6836 : _GEN10539;
wire  _GEN10541 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10542 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10543 = io_x[6] ? _GEN10542 : _GEN10541;
wire  _GEN10544 = io_x[41] ? _GEN6836 : _GEN10543;
wire  _GEN10545 = io_x[14] ? _GEN10544 : _GEN10540;
wire  _GEN10546 = io_x[0] ? _GEN10545 : _GEN6845;
wire  _GEN10547 = io_x[76] ? _GEN10546 : _GEN10538;
wire  _GEN10548 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10549 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10550 = io_x[6] ? _GEN10549 : _GEN6850;
wire  _GEN10551 = io_x[41] ? _GEN6836 : _GEN10550;
wire  _GEN10552 = io_x[14] ? _GEN10551 : _GEN6843;
wire  _GEN10553 = io_x[0] ? _GEN10552 : _GEN10548;
wire  _GEN10554 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10555 = io_x[41] ? _GEN6836 : _GEN10554;
wire  _GEN10556 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10557 = io_x[41] ? _GEN6924 : _GEN10556;
wire  _GEN10558 = io_x[14] ? _GEN10557 : _GEN10555;
wire  _GEN10559 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10560 = io_x[0] ? _GEN10559 : _GEN10558;
wire  _GEN10561 = io_x[76] ? _GEN10560 : _GEN10553;
wire  _GEN10562 = io_x[42] ? _GEN10561 : _GEN10547;
wire  _GEN10563 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10564 = io_x[41] ? _GEN6924 : _GEN10563;
wire  _GEN10565 = io_x[14] ? _GEN10564 : _GEN6856;
wire  _GEN10566 = io_x[0] ? _GEN10565 : _GEN6845;
wire  _GEN10567 = io_x[76] ? _GEN10566 : _GEN6833;
wire  _GEN10568 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10569 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10570 = io_x[6] ? _GEN10569 : _GEN10568;
wire  _GEN10571 = io_x[41] ? _GEN6836 : _GEN10570;
wire  _GEN10572 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10573 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10574 = io_x[6] ? _GEN10573 : _GEN10572;
wire  _GEN10575 = io_x[41] ? _GEN6836 : _GEN10574;
wire  _GEN10576 = io_x[14] ? _GEN10575 : _GEN10571;
wire  _GEN10577 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10578 = io_x[41] ? _GEN6836 : _GEN10577;
wire  _GEN10579 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10580 = io_x[41] ? _GEN6836 : _GEN10579;
wire  _GEN10581 = io_x[14] ? _GEN10580 : _GEN10578;
wire  _GEN10582 = io_x[0] ? _GEN10581 : _GEN10576;
wire  _GEN10583 = io_x[76] ? _GEN6834 : _GEN10582;
wire  _GEN10584 = io_x[42] ? _GEN10583 : _GEN10567;
wire  _GEN10585 = io_x[38] ? _GEN10584 : _GEN10562;
wire  _GEN10586 = io_x[10] ? _GEN10585 : _GEN10536;
wire  _GEN10587 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10588 = io_x[41] ? _GEN6836 : _GEN10587;
wire  _GEN10589 = io_x[14] ? _GEN10588 : _GEN6843;
wire  _GEN10590 = io_x[0] ? _GEN6845 : _GEN10589;
wire  _GEN10591 = io_x[76] ? _GEN6834 : _GEN10590;
wire  _GEN10592 = io_x[42] ? _GEN6863 : _GEN10591;
wire  _GEN10593 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN10594 = io_x[14] ? _GEN10593 : _GEN6843;
wire  _GEN10595 = io_x[0] ? _GEN6845 : _GEN10594;
wire  _GEN10596 = io_x[76] ? _GEN6834 : _GEN10595;
wire  _GEN10597 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10598 = io_x[2] ? _GEN6838 : _GEN10597;
wire  _GEN10599 = io_x[6] ? _GEN6850 : _GEN10598;
wire  _GEN10600 = io_x[41] ? _GEN6836 : _GEN10599;
wire  _GEN10601 = io_x[14] ? _GEN6843 : _GEN10600;
wire  _GEN10602 = io_x[0] ? _GEN6858 : _GEN10601;
wire  _GEN10603 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN10604 = io_x[14] ? _GEN6843 : _GEN10603;
wire  _GEN10605 = io_x[0] ? _GEN6845 : _GEN10604;
wire  _GEN10606 = io_x[76] ? _GEN10605 : _GEN10602;
wire  _GEN10607 = io_x[42] ? _GEN10606 : _GEN10596;
wire  _GEN10608 = io_x[38] ? _GEN10607 : _GEN10592;
wire  _GEN10609 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10610 = io_x[41] ? _GEN6836 : _GEN10609;
wire  _GEN10611 = io_x[14] ? _GEN10610 : _GEN6843;
wire  _GEN10612 = io_x[0] ? _GEN6858 : _GEN10611;
wire  _GEN10613 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN10614 = io_x[14] ? _GEN6843 : _GEN10613;
wire  _GEN10615 = io_x[0] ? _GEN10614 : _GEN6845;
wire  _GEN10616 = io_x[76] ? _GEN10615 : _GEN10612;
wire  _GEN10617 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10618 = io_x[0] ? _GEN10617 : _GEN6858;
wire  _GEN10619 = io_x[76] ? _GEN6834 : _GEN10618;
wire  _GEN10620 = io_x[42] ? _GEN10619 : _GEN10616;
wire  _GEN10621 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN10622 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10623 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10624 = io_x[41] ? _GEN6836 : _GEN10623;
wire  _GEN10625 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10626 = io_x[41] ? _GEN6836 : _GEN10625;
wire  _GEN10627 = io_x[14] ? _GEN10626 : _GEN10624;
wire  _GEN10628 = io_x[0] ? _GEN10627 : _GEN10622;
wire  _GEN10629 = io_x[76] ? _GEN6834 : _GEN10628;
wire  _GEN10630 = io_x[42] ? _GEN10629 : _GEN10621;
wire  _GEN10631 = io_x[38] ? _GEN10630 : _GEN10620;
wire  _GEN10632 = io_x[10] ? _GEN10631 : _GEN10608;
wire  _GEN10633 = io_x[71] ? _GEN10632 : _GEN10586;
wire  _GEN10634 = io_x[70] ? _GEN10633 : _GEN10510;
wire  _GEN10635 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN10636 = io_x[14] ? _GEN6843 : _GEN10635;
wire  _GEN10637 = io_x[0] ? _GEN6858 : _GEN10636;
wire  _GEN10638 = io_x[76] ? _GEN10637 : _GEN6833;
wire  _GEN10639 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10640 = io_x[41] ? _GEN6836 : _GEN10639;
wire  _GEN10641 = io_x[14] ? _GEN10640 : _GEN6856;
wire  _GEN10642 = io_x[0] ? _GEN10641 : _GEN6845;
wire  _GEN10643 = io_x[76] ? _GEN6834 : _GEN10642;
wire  _GEN10644 = io_x[42] ? _GEN10643 : _GEN10638;
wire  _GEN10645 = io_x[38] ? _GEN10644 : _GEN7036;
wire  _GEN10646 = io_x[10] ? _GEN10645 : _GEN7044;
wire  _GEN10647 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN10648 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10649 = io_x[6] ? _GEN6850 : _GEN10648;
wire  _GEN10650 = io_x[41] ? _GEN6836 : _GEN10649;
wire  _GEN10651 = io_x[14] ? _GEN6856 : _GEN10650;
wire  _GEN10652 = io_x[0] ? _GEN10651 : _GEN6845;
wire  _GEN10653 = io_x[76] ? _GEN6834 : _GEN10652;
wire  _GEN10654 = io_x[42] ? _GEN10653 : _GEN6874;
wire  _GEN10655 = io_x[38] ? _GEN10654 : _GEN10647;
wire  _GEN10656 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10657 = io_x[41] ? _GEN10656 : _GEN6836;
wire  _GEN10658 = io_x[14] ? _GEN6856 : _GEN10657;
wire  _GEN10659 = io_x[0] ? _GEN10658 : _GEN6845;
wire  _GEN10660 = io_x[76] ? _GEN6834 : _GEN10659;
wire  _GEN10661 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10662 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10663 = io_x[6] ? _GEN10662 : _GEN10661;
wire  _GEN10664 = io_x[41] ? _GEN6836 : _GEN10663;
wire  _GEN10665 = io_x[14] ? _GEN10664 : _GEN6843;
wire  _GEN10666 = io_x[0] ? _GEN10665 : _GEN6845;
wire  _GEN10667 = io_x[76] ? _GEN6834 : _GEN10666;
wire  _GEN10668 = io_x[42] ? _GEN10667 : _GEN10660;
wire  _GEN10669 = io_x[38] ? _GEN10668 : _GEN6871;
wire  _GEN10670 = io_x[10] ? _GEN10669 : _GEN10655;
wire  _GEN10671 = io_x[71] ? _GEN10670 : _GEN10646;
wire  _GEN10672 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10673 = io_x[6] ? _GEN6840 : _GEN10672;
wire  _GEN10674 = io_x[41] ? _GEN10673 : _GEN6836;
wire  _GEN10675 = io_x[14] ? _GEN10674 : _GEN6843;
wire  _GEN10676 = io_x[0] ? _GEN10675 : _GEN6845;
wire  _GEN10677 = io_x[76] ? _GEN10676 : _GEN6834;
wire  _GEN10678 = io_x[42] ? _GEN6874 : _GEN10677;
wire  _GEN10679 = io_x[38] ? _GEN10678 : _GEN7036;
wire  _GEN10680 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10681 = io_x[0] ? _GEN10680 : _GEN6845;
wire  _GEN10682 = io_x[76] ? _GEN6833 : _GEN10681;
wire  _GEN10683 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN10684 = io_x[42] ? _GEN10683 : _GEN10682;
wire  _GEN10685 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10686 = io_x[41] ? _GEN10685 : _GEN6924;
wire  _GEN10687 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10688 = io_x[41] ? _GEN10687 : _GEN6836;
wire  _GEN10689 = io_x[14] ? _GEN10688 : _GEN10686;
wire  _GEN10690 = io_x[0] ? _GEN10689 : _GEN6845;
wire  _GEN10691 = io_x[76] ? _GEN10690 : _GEN6833;
wire  _GEN10692 = io_x[42] ? _GEN6874 : _GEN10691;
wire  _GEN10693 = io_x[38] ? _GEN10692 : _GEN10684;
wire  _GEN10694 = io_x[10] ? _GEN10693 : _GEN10679;
wire  _GEN10695 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN10696 = io_x[71] ? _GEN10695 : _GEN10694;
wire  _GEN10697 = io_x[70] ? _GEN10696 : _GEN10671;
wire  _GEN10698 = io_x[33] ? _GEN10697 : _GEN10634;
wire  _GEN10699 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN10700 = io_x[76] ? _GEN6834 : _GEN10699;
wire  _GEN10701 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10702 = io_x[2] ? _GEN6837 : _GEN10701;
wire  _GEN10703 = io_x[6] ? _GEN6850 : _GEN10702;
wire  _GEN10704 = io_x[41] ? _GEN10703 : _GEN6836;
wire  _GEN10705 = io_x[14] ? _GEN6843 : _GEN10704;
wire  _GEN10706 = io_x[0] ? _GEN6845 : _GEN10705;
wire  _GEN10707 = io_x[76] ? _GEN6834 : _GEN10706;
wire  _GEN10708 = io_x[42] ? _GEN10707 : _GEN10700;
wire  _GEN10709 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10710 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10711 = io_x[6] ? _GEN10710 : _GEN6850;
wire  _GEN10712 = io_x[41] ? _GEN6836 : _GEN10711;
wire  _GEN10713 = io_x[14] ? _GEN6843 : _GEN10712;
wire  _GEN10714 = io_x[0] ? _GEN10713 : _GEN10709;
wire  _GEN10715 = io_x[76] ? _GEN6833 : _GEN10714;
wire  _GEN10716 = io_x[42] ? _GEN10715 : _GEN6863;
wire  _GEN10717 = io_x[38] ? _GEN10716 : _GEN10708;
wire  _GEN10718 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN10719 = io_x[14] ? _GEN6856 : _GEN10718;
wire  _GEN10720 = io_x[0] ? _GEN10719 : _GEN6858;
wire  _GEN10721 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN10722 = io_x[76] ? _GEN10721 : _GEN10720;
wire  _GEN10723 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10724 = io_x[41] ? _GEN6924 : _GEN10723;
wire  _GEN10725 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10726 = io_x[41] ? _GEN6836 : _GEN10725;
wire  _GEN10727 = io_x[14] ? _GEN10726 : _GEN10724;
wire  _GEN10728 = io_x[0] ? _GEN10727 : _GEN6858;
wire  _GEN10729 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10730 = io_x[2] ? _GEN10729 : _GEN6837;
wire  _GEN10731 = io_x[6] ? _GEN10730 : _GEN6850;
wire  _GEN10732 = io_x[41] ? _GEN10731 : _GEN6836;
wire  _GEN10733 = io_x[14] ? _GEN10732 : _GEN6843;
wire  _GEN10734 = io_x[0] ? _GEN6858 : _GEN10733;
wire  _GEN10735 = io_x[76] ? _GEN10734 : _GEN10728;
wire  _GEN10736 = io_x[42] ? _GEN10735 : _GEN10722;
wire  _GEN10737 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10738 = io_x[41] ? _GEN6836 : _GEN10737;
wire  _GEN10739 = io_x[14] ? _GEN10738 : _GEN6843;
wire  _GEN10740 = io_x[0] ? _GEN10739 : _GEN6858;
wire  _GEN10741 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10742 = io_x[41] ? _GEN6924 : _GEN10741;
wire  _GEN10743 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10744 = io_x[41] ? _GEN6836 : _GEN10743;
wire  _GEN10745 = io_x[14] ? _GEN10744 : _GEN10742;
wire  _GEN10746 = io_x[0] ? _GEN10745 : _GEN6845;
wire  _GEN10747 = io_x[76] ? _GEN10746 : _GEN10740;
wire  _GEN10748 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10749 = io_x[6] ? _GEN10748 : _GEN6850;
wire  _GEN10750 = io_x[41] ? _GEN6924 : _GEN10749;
wire  _GEN10751 = io_x[14] ? _GEN10750 : _GEN6843;
wire  _GEN10752 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10753 = io_x[6] ? _GEN10752 : _GEN6840;
wire  _GEN10754 = io_x[41] ? _GEN6836 : _GEN10753;
wire  _GEN10755 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10756 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10757 = io_x[6] ? _GEN10756 : _GEN10755;
wire  _GEN10758 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10759 = io_x[41] ? _GEN10758 : _GEN10757;
wire  _GEN10760 = io_x[14] ? _GEN10759 : _GEN10754;
wire  _GEN10761 = io_x[0] ? _GEN10760 : _GEN10751;
wire  _GEN10762 = io_x[76] ? _GEN6834 : _GEN10761;
wire  _GEN10763 = io_x[42] ? _GEN10762 : _GEN10747;
wire  _GEN10764 = io_x[38] ? _GEN10763 : _GEN10736;
wire  _GEN10765 = io_x[10] ? _GEN10764 : _GEN10717;
wire  _GEN10766 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10767 = io_x[41] ? _GEN10766 : _GEN6836;
wire  _GEN10768 = io_x[14] ? _GEN10767 : _GEN6843;
wire  _GEN10769 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10770 = io_x[0] ? _GEN10769 : _GEN10768;
wire  _GEN10771 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10772 = io_x[0] ? _GEN6845 : _GEN10771;
wire  _GEN10773 = io_x[76] ? _GEN10772 : _GEN10770;
wire  _GEN10774 = io_x[42] ? _GEN10773 : _GEN6874;
wire  _GEN10775 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10776 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10777 = io_x[6] ? _GEN10776 : _GEN6850;
wire  _GEN10778 = io_x[41] ? _GEN6836 : _GEN10777;
wire  _GEN10779 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10780 = io_x[6] ? _GEN10779 : _GEN6840;
wire  _GEN10781 = io_x[41] ? _GEN6836 : _GEN10780;
wire  _GEN10782 = io_x[14] ? _GEN10781 : _GEN10778;
wire  _GEN10783 = io_x[0] ? _GEN10782 : _GEN10775;
wire  _GEN10784 = io_x[76] ? _GEN6834 : _GEN10783;
wire  _GEN10785 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10786 = io_x[2] ? _GEN6837 : _GEN10785;
wire  _GEN10787 = io_x[6] ? _GEN6850 : _GEN10786;
wire  _GEN10788 = io_x[41] ? _GEN10787 : _GEN6924;
wire  _GEN10789 = io_x[14] ? _GEN6843 : _GEN10788;
wire  _GEN10790 = io_x[0] ? _GEN6845 : _GEN10789;
wire  _GEN10791 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10792 = io_x[2] ? _GEN6837 : _GEN10791;
wire  _GEN10793 = io_x[6] ? _GEN6850 : _GEN10792;
wire  _GEN10794 = io_x[41] ? _GEN10793 : _GEN6836;
wire  _GEN10795 = io_x[14] ? _GEN6843 : _GEN10794;
wire  _GEN10796 = io_x[0] ? _GEN6845 : _GEN10795;
wire  _GEN10797 = io_x[76] ? _GEN10796 : _GEN10790;
wire  _GEN10798 = io_x[42] ? _GEN10797 : _GEN10784;
wire  _GEN10799 = io_x[38] ? _GEN10798 : _GEN10774;
wire  _GEN10800 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN10801 = io_x[14] ? _GEN10800 : _GEN6856;
wire  _GEN10802 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10803 = io_x[41] ? _GEN6836 : _GEN10802;
wire  _GEN10804 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10805 = io_x[41] ? _GEN6836 : _GEN10804;
wire  _GEN10806 = io_x[14] ? _GEN10805 : _GEN10803;
wire  _GEN10807 = io_x[0] ? _GEN10806 : _GEN10801;
wire  _GEN10808 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10809 = io_x[41] ? _GEN6836 : _GEN10808;
wire  _GEN10810 = io_x[14] ? _GEN10809 : _GEN6856;
wire  _GEN10811 = io_x[0] ? _GEN6845 : _GEN10810;
wire  _GEN10812 = io_x[76] ? _GEN10811 : _GEN10807;
wire  _GEN10813 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10814 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN10815 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10816 = io_x[6] ? _GEN10815 : _GEN6850;
wire  _GEN10817 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10818 = io_x[2] ? _GEN10817 : _GEN6837;
wire  _GEN10819 = io_x[6] ? _GEN10818 : _GEN6850;
wire  _GEN10820 = io_x[41] ? _GEN10819 : _GEN10816;
wire  _GEN10821 = io_x[14] ? _GEN10820 : _GEN10814;
wire  _GEN10822 = io_x[0] ? _GEN10821 : _GEN10813;
wire  _GEN10823 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10824 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10825 = io_x[0] ? _GEN10824 : _GEN10823;
wire  _GEN10826 = io_x[76] ? _GEN10825 : _GEN10822;
wire  _GEN10827 = io_x[42] ? _GEN10826 : _GEN10812;
wire  _GEN10828 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10829 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10830 = io_x[6] ? _GEN6850 : _GEN10829;
wire  _GEN10831 = io_x[41] ? _GEN6836 : _GEN10830;
wire  _GEN10832 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10833 = io_x[2] ? _GEN10832 : _GEN6837;
wire  _GEN10834 = io_x[6] ? _GEN10833 : _GEN6840;
wire  _GEN10835 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10836 = io_x[6] ? _GEN10835 : _GEN6850;
wire  _GEN10837 = io_x[41] ? _GEN10836 : _GEN10834;
wire  _GEN10838 = io_x[14] ? _GEN10837 : _GEN10831;
wire  _GEN10839 = io_x[0] ? _GEN10838 : _GEN10828;
wire  _GEN10840 = io_x[76] ? _GEN6834 : _GEN10839;
wire  _GEN10841 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10842 = io_x[6] ? _GEN10841 : _GEN6840;
wire  _GEN10843 = io_x[41] ? _GEN6836 : _GEN10842;
wire  _GEN10844 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10845 = io_x[41] ? _GEN6836 : _GEN10844;
wire  _GEN10846 = io_x[14] ? _GEN10845 : _GEN10843;
wire  _GEN10847 = io_x[0] ? _GEN10846 : _GEN6858;
wire  _GEN10848 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN10849 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10850 = io_x[0] ? _GEN10849 : _GEN10848;
wire  _GEN10851 = io_x[76] ? _GEN10850 : _GEN10847;
wire  _GEN10852 = io_x[42] ? _GEN10851 : _GEN10840;
wire  _GEN10853 = io_x[38] ? _GEN10852 : _GEN10827;
wire  _GEN10854 = io_x[10] ? _GEN10853 : _GEN10799;
wire  _GEN10855 = io_x[71] ? _GEN10854 : _GEN10765;
wire  _GEN10856 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN10857 = io_x[0] ? _GEN6845 : _GEN10856;
wire  _GEN10858 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10859 = io_x[6] ? _GEN10858 : _GEN6840;
wire  _GEN10860 = io_x[41] ? _GEN6836 : _GEN10859;
wire  _GEN10861 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10862 = io_x[6] ? _GEN10861 : _GEN6850;
wire  _GEN10863 = io_x[41] ? _GEN6836 : _GEN10862;
wire  _GEN10864 = io_x[14] ? _GEN10863 : _GEN10860;
wire  _GEN10865 = io_x[0] ? _GEN10864 : _GEN6845;
wire  _GEN10866 = io_x[76] ? _GEN10865 : _GEN10857;
wire  _GEN10867 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN10868 = io_x[14] ? _GEN6843 : _GEN10867;
wire  _GEN10869 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10870 = io_x[41] ? _GEN6836 : _GEN10869;
wire  _GEN10871 = io_x[14] ? _GEN10870 : _GEN6856;
wire  _GEN10872 = io_x[0] ? _GEN10871 : _GEN10868;
wire  _GEN10873 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10874 = io_x[2] ? _GEN6837 : _GEN10873;
wire  _GEN10875 = io_x[6] ? _GEN6840 : _GEN10874;
wire  _GEN10876 = io_x[41] ? _GEN10875 : _GEN6836;
wire  _GEN10877 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN10878 = io_x[14] ? _GEN10877 : _GEN10876;
wire  _GEN10879 = io_x[0] ? _GEN6845 : _GEN10878;
wire  _GEN10880 = io_x[76] ? _GEN10879 : _GEN10872;
wire  _GEN10881 = io_x[42] ? _GEN10880 : _GEN10866;
wire  _GEN10882 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10883 = io_x[41] ? _GEN10882 : _GEN6836;
wire  _GEN10884 = io_x[14] ? _GEN6843 : _GEN10883;
wire  _GEN10885 = io_x[0] ? _GEN6858 : _GEN10884;
wire  _GEN10886 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN10887 = io_x[76] ? _GEN10886 : _GEN10885;
wire  _GEN10888 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10889 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10890 = io_x[6] ? _GEN10889 : _GEN10888;
wire  _GEN10891 = io_x[41] ? _GEN6924 : _GEN10890;
wire  _GEN10892 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10893 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10894 = io_x[6] ? _GEN10893 : _GEN10892;
wire  _GEN10895 = io_x[41] ? _GEN6836 : _GEN10894;
wire  _GEN10896 = io_x[14] ? _GEN10895 : _GEN10891;
wire  _GEN10897 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10898 = io_x[41] ? _GEN6836 : _GEN10897;
wire  _GEN10899 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10900 = io_x[41] ? _GEN6836 : _GEN10899;
wire  _GEN10901 = io_x[14] ? _GEN10900 : _GEN10898;
wire  _GEN10902 = io_x[0] ? _GEN10901 : _GEN10896;
wire  _GEN10903 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10904 = io_x[2] ? _GEN6837 : _GEN10903;
wire  _GEN10905 = io_x[6] ? _GEN6850 : _GEN10904;
wire  _GEN10906 = io_x[41] ? _GEN10905 : _GEN6836;
wire  _GEN10907 = io_x[14] ? _GEN6843 : _GEN10906;
wire  _GEN10908 = io_x[0] ? _GEN6845 : _GEN10907;
wire  _GEN10909 = io_x[76] ? _GEN10908 : _GEN10902;
wire  _GEN10910 = io_x[42] ? _GEN10909 : _GEN10887;
wire  _GEN10911 = io_x[38] ? _GEN10910 : _GEN10881;
wire  _GEN10912 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10913 = io_x[41] ? _GEN6924 : _GEN10912;
wire  _GEN10914 = io_x[14] ? _GEN10913 : _GEN6843;
wire  _GEN10915 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10916 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10917 = io_x[6] ? _GEN10916 : _GEN6840;
wire  _GEN10918 = io_x[41] ? _GEN10917 : _GEN10915;
wire  _GEN10919 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10920 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10921 = io_x[6] ? _GEN10920 : _GEN6850;
wire  _GEN10922 = io_x[41] ? _GEN10921 : _GEN10919;
wire  _GEN10923 = io_x[14] ? _GEN10922 : _GEN10918;
wire  _GEN10924 = io_x[0] ? _GEN10923 : _GEN10914;
wire  _GEN10925 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10926 = io_x[6] ? _GEN10925 : _GEN6840;
wire  _GEN10927 = io_x[41] ? _GEN6836 : _GEN10926;
wire  _GEN10928 = io_x[14] ? _GEN10927 : _GEN6856;
wire  _GEN10929 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10930 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10931 = io_x[6] ? _GEN10930 : _GEN10929;
wire  _GEN10932 = io_x[41] ? _GEN6836 : _GEN10931;
wire  _GEN10933 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10934 = io_x[6] ? _GEN10933 : _GEN6840;
wire  _GEN10935 = io_x[41] ? _GEN6836 : _GEN10934;
wire  _GEN10936 = io_x[14] ? _GEN10935 : _GEN10932;
wire  _GEN10937 = io_x[0] ? _GEN10936 : _GEN10928;
wire  _GEN10938 = io_x[76] ? _GEN10937 : _GEN10924;
wire  _GEN10939 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10940 = io_x[41] ? _GEN6836 : _GEN10939;
wire  _GEN10941 = io_x[14] ? _GEN10940 : _GEN6843;
wire  _GEN10942 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10943 = io_x[6] ? _GEN10942 : _GEN6840;
wire  _GEN10944 = io_x[41] ? _GEN6836 : _GEN10943;
wire  _GEN10945 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10946 = io_x[6] ? _GEN6840 : _GEN10945;
wire  _GEN10947 = io_x[41] ? _GEN6924 : _GEN10946;
wire  _GEN10948 = io_x[14] ? _GEN10947 : _GEN10944;
wire  _GEN10949 = io_x[0] ? _GEN10948 : _GEN10941;
wire  _GEN10950 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10951 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10952 = io_x[2] ? _GEN10951 : _GEN6837;
wire  _GEN10953 = io_x[6] ? _GEN10952 : _GEN6850;
wire  _GEN10954 = io_x[41] ? _GEN10953 : _GEN10950;
wire  _GEN10955 = io_x[14] ? _GEN10954 : _GEN6843;
wire  _GEN10956 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10957 = io_x[41] ? _GEN6836 : _GEN10956;
wire  _GEN10958 = io_x[14] ? _GEN6843 : _GEN10957;
wire  _GEN10959 = io_x[0] ? _GEN10958 : _GEN10955;
wire  _GEN10960 = io_x[76] ? _GEN10959 : _GEN10949;
wire  _GEN10961 = io_x[42] ? _GEN10960 : _GEN10938;
wire  _GEN10962 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10963 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10964 = io_x[6] ? _GEN10963 : _GEN10962;
wire  _GEN10965 = io_x[41] ? _GEN10964 : _GEN6924;
wire  _GEN10966 = io_x[14] ? _GEN10965 : _GEN6843;
wire  _GEN10967 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN10968 = io_x[14] ? _GEN10967 : _GEN6843;
wire  _GEN10969 = io_x[0] ? _GEN10968 : _GEN10966;
wire  _GEN10970 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10971 = io_x[41] ? _GEN6924 : _GEN10970;
wire  _GEN10972 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10973 = io_x[41] ? _GEN6924 : _GEN10972;
wire  _GEN10974 = io_x[14] ? _GEN10973 : _GEN10971;
wire  _GEN10975 = io_x[0] ? _GEN10974 : _GEN6845;
wire  _GEN10976 = io_x[76] ? _GEN10975 : _GEN10969;
wire  _GEN10977 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10978 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10979 = io_x[6] ? _GEN10978 : _GEN10977;
wire  _GEN10980 = io_x[41] ? _GEN6836 : _GEN10979;
wire  _GEN10981 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN10982 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN10983 = io_x[6] ? _GEN10982 : _GEN10981;
wire  _GEN10984 = io_x[41] ? _GEN6924 : _GEN10983;
wire  _GEN10985 = io_x[14] ? _GEN10984 : _GEN10980;
wire  _GEN10986 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN10987 = io_x[41] ? _GEN6836 : _GEN10986;
wire  _GEN10988 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN10989 = io_x[41] ? _GEN6836 : _GEN10988;
wire  _GEN10990 = io_x[14] ? _GEN10989 : _GEN10987;
wire  _GEN10991 = io_x[0] ? _GEN10990 : _GEN10985;
wire  _GEN10992 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN10993 = io_x[2] ? _GEN10992 : _GEN6837;
wire  _GEN10994 = io_x[6] ? _GEN10993 : _GEN6850;
wire  _GEN10995 = io_x[41] ? _GEN10994 : _GEN6836;
wire  _GEN10996 = io_x[14] ? _GEN10995 : _GEN6843;
wire  _GEN10997 = io_x[0] ? _GEN6845 : _GEN10996;
wire  _GEN10998 = io_x[76] ? _GEN10997 : _GEN10991;
wire  _GEN10999 = io_x[42] ? _GEN10998 : _GEN10976;
wire  _GEN11000 = io_x[38] ? _GEN10999 : _GEN10961;
wire  _GEN11001 = io_x[10] ? _GEN11000 : _GEN10911;
wire  _GEN11002 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11003 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11004 = io_x[6] ? _GEN11003 : _GEN6850;
wire  _GEN11005 = io_x[41] ? _GEN6836 : _GEN11004;
wire  _GEN11006 = io_x[14] ? _GEN11005 : _GEN6843;
wire  _GEN11007 = io_x[0] ? _GEN11006 : _GEN11002;
wire  _GEN11008 = io_x[76] ? _GEN6834 : _GEN11007;
wire  _GEN11009 = io_x[42] ? _GEN6863 : _GEN11008;
wire  _GEN11010 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11011 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN11012 = io_x[14] ? _GEN11011 : _GEN11010;
wire  _GEN11013 = io_x[0] ? _GEN11012 : _GEN6858;
wire  _GEN11014 = io_x[76] ? _GEN6834 : _GEN11013;
wire  _GEN11015 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11016 = io_x[2] ? _GEN6838 : _GEN11015;
wire  _GEN11017 = io_x[6] ? _GEN6850 : _GEN11016;
wire  _GEN11018 = io_x[41] ? _GEN6836 : _GEN11017;
wire  _GEN11019 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11020 = io_x[41] ? _GEN6836 : _GEN11019;
wire  _GEN11021 = io_x[14] ? _GEN11020 : _GEN11018;
wire  _GEN11022 = io_x[0] ? _GEN6845 : _GEN11021;
wire  _GEN11023 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN11024 = io_x[14] ? _GEN6843 : _GEN11023;
wire  _GEN11025 = io_x[0] ? _GEN6845 : _GEN11024;
wire  _GEN11026 = io_x[76] ? _GEN11025 : _GEN11022;
wire  _GEN11027 = io_x[42] ? _GEN11026 : _GEN11014;
wire  _GEN11028 = io_x[38] ? _GEN11027 : _GEN11009;
wire  _GEN11029 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11030 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11031 = io_x[6] ? _GEN6840 : _GEN11030;
wire  _GEN11032 = io_x[41] ? _GEN11031 : _GEN11029;
wire  _GEN11033 = io_x[14] ? _GEN11032 : _GEN6843;
wire  _GEN11034 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11035 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11036 = io_x[41] ? _GEN11035 : _GEN11034;
wire  _GEN11037 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11038 = io_x[6] ? _GEN11037 : _GEN6850;
wire  _GEN11039 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11040 = io_x[6] ? _GEN6840 : _GEN11039;
wire  _GEN11041 = io_x[41] ? _GEN11040 : _GEN11038;
wire  _GEN11042 = io_x[14] ? _GEN11041 : _GEN11036;
wire  _GEN11043 = io_x[0] ? _GEN11042 : _GEN11033;
wire  _GEN11044 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11045 = io_x[41] ? _GEN11044 : _GEN6836;
wire  _GEN11046 = io_x[14] ? _GEN11045 : _GEN6843;
wire  _GEN11047 = io_x[0] ? _GEN6845 : _GEN11046;
wire  _GEN11048 = io_x[76] ? _GEN11047 : _GEN11043;
wire  _GEN11049 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11050 = io_x[41] ? _GEN6924 : _GEN11049;
wire  _GEN11051 = io_x[14] ? _GEN11050 : _GEN6843;
wire  _GEN11052 = io_x[0] ? _GEN11051 : _GEN6845;
wire  _GEN11053 = io_x[76] ? _GEN6834 : _GEN11052;
wire  _GEN11054 = io_x[42] ? _GEN11053 : _GEN11048;
wire  _GEN11055 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11056 = io_x[2] ? _GEN11055 : _GEN6837;
wire  _GEN11057 = io_x[6] ? _GEN11056 : _GEN6850;
wire  _GEN11058 = io_x[41] ? _GEN11057 : _GEN6924;
wire  _GEN11059 = io_x[14] ? _GEN11058 : _GEN6843;
wire  _GEN11060 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11061 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11062 = io_x[41] ? _GEN6836 : _GEN11061;
wire  _GEN11063 = io_x[14] ? _GEN11062 : _GEN11060;
wire  _GEN11064 = io_x[0] ? _GEN11063 : _GEN11059;
wire  _GEN11065 = io_x[76] ? _GEN6834 : _GEN11064;
wire  _GEN11066 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11067 = io_x[41] ? _GEN6836 : _GEN11066;
wire  _GEN11068 = io_x[14] ? _GEN6843 : _GEN11067;
wire  _GEN11069 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11070 = io_x[41] ? _GEN6836 : _GEN11069;
wire  _GEN11071 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11072 = io_x[41] ? _GEN6924 : _GEN11071;
wire  _GEN11073 = io_x[14] ? _GEN11072 : _GEN11070;
wire  _GEN11074 = io_x[0] ? _GEN11073 : _GEN11068;
wire  _GEN11075 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN11076 = io_x[76] ? _GEN11075 : _GEN11074;
wire  _GEN11077 = io_x[42] ? _GEN11076 : _GEN11065;
wire  _GEN11078 = io_x[38] ? _GEN11077 : _GEN11054;
wire  _GEN11079 = io_x[10] ? _GEN11078 : _GEN11028;
wire  _GEN11080 = io_x[71] ? _GEN11079 : _GEN11001;
wire  _GEN11081 = io_x[70] ? _GEN11080 : _GEN10855;
wire  _GEN11082 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11083 = io_x[41] ? _GEN11082 : _GEN6836;
wire  _GEN11084 = io_x[14] ? _GEN11083 : _GEN6843;
wire  _GEN11085 = io_x[0] ? _GEN11084 : _GEN6845;
wire  _GEN11086 = io_x[76] ? _GEN6834 : _GEN11085;
wire  _GEN11087 = io_x[42] ? _GEN6874 : _GEN11086;
wire  _GEN11088 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11089 = io_x[41] ? _GEN6836 : _GEN11088;
wire  _GEN11090 = io_x[14] ? _GEN6843 : _GEN11089;
wire  _GEN11091 = io_x[0] ? _GEN11090 : _GEN6845;
wire  _GEN11092 = io_x[76] ? _GEN6834 : _GEN11091;
wire  _GEN11093 = io_x[42] ? _GEN11092 : _GEN6863;
wire  _GEN11094 = io_x[38] ? _GEN11093 : _GEN11087;
wire  _GEN11095 = io_x[10] ? _GEN11094 : _GEN7044;
wire  _GEN11096 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN11097 = io_x[42] ? _GEN6874 : _GEN11096;
wire  _GEN11098 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN11099 = io_x[76] ? _GEN6834 : _GEN11098;
wire  _GEN11100 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11101 = io_x[6] ? _GEN6850 : _GEN11100;
wire  _GEN11102 = io_x[41] ? _GEN6836 : _GEN11101;
wire  _GEN11103 = io_x[14] ? _GEN6843 : _GEN11102;
wire  _GEN11104 = io_x[0] ? _GEN11103 : _GEN6845;
wire  _GEN11105 = io_x[76] ? _GEN6834 : _GEN11104;
wire  _GEN11106 = io_x[42] ? _GEN11105 : _GEN11099;
wire  _GEN11107 = io_x[38] ? _GEN11106 : _GEN11097;
wire  _GEN11108 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11109 = io_x[0] ? _GEN6845 : _GEN11108;
wire  _GEN11110 = io_x[76] ? _GEN6834 : _GEN11109;
wire  _GEN11111 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11112 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11113 = io_x[0] ? _GEN11112 : _GEN11111;
wire  _GEN11114 = io_x[76] ? _GEN6834 : _GEN11113;
wire  _GEN11115 = io_x[42] ? _GEN11114 : _GEN11110;
wire  _GEN11116 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11117 = io_x[41] ? _GEN11116 : _GEN6836;
wire  _GEN11118 = io_x[14] ? _GEN11117 : _GEN6843;
wire  _GEN11119 = io_x[0] ? _GEN11118 : _GEN6845;
wire  _GEN11120 = io_x[76] ? _GEN6834 : _GEN11119;
wire  _GEN11121 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11122 = io_x[6] ? _GEN6850 : _GEN11121;
wire  _GEN11123 = io_x[41] ? _GEN6836 : _GEN11122;
wire  _GEN11124 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11125 = io_x[41] ? _GEN6836 : _GEN11124;
wire  _GEN11126 = io_x[14] ? _GEN11125 : _GEN11123;
wire  _GEN11127 = io_x[0] ? _GEN11126 : _GEN6845;
wire  _GEN11128 = io_x[76] ? _GEN6834 : _GEN11127;
wire  _GEN11129 = io_x[42] ? _GEN11128 : _GEN11120;
wire  _GEN11130 = io_x[38] ? _GEN11129 : _GEN11115;
wire  _GEN11131 = io_x[10] ? _GEN11130 : _GEN11107;
wire  _GEN11132 = io_x[71] ? _GEN11131 : _GEN11095;
wire  _GEN11133 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11134 = io_x[41] ? _GEN6836 : _GEN11133;
wire  _GEN11135 = io_x[14] ? _GEN11134 : _GEN6843;
wire  _GEN11136 = io_x[0] ? _GEN11135 : _GEN6845;
wire  _GEN11137 = io_x[76] ? _GEN6834 : _GEN11136;
wire  _GEN11138 = io_x[42] ? _GEN11137 : _GEN6874;
wire  _GEN11139 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN11140 = io_x[76] ? _GEN11139 : _GEN6834;
wire  _GEN11141 = io_x[42] ? _GEN6874 : _GEN11140;
wire  _GEN11142 = io_x[38] ? _GEN11141 : _GEN11138;
wire  _GEN11143 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11144 = io_x[41] ? _GEN6836 : _GEN11143;
wire  _GEN11145 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11146 = io_x[41] ? _GEN6836 : _GEN11145;
wire  _GEN11147 = io_x[14] ? _GEN11146 : _GEN11144;
wire  _GEN11148 = io_x[0] ? _GEN11147 : _GEN6845;
wire  _GEN11149 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11150 = io_x[41] ? _GEN6836 : _GEN11149;
wire  _GEN11151 = io_x[14] ? _GEN11150 : _GEN6856;
wire  _GEN11152 = io_x[0] ? _GEN11151 : _GEN6845;
wire  _GEN11153 = io_x[76] ? _GEN11152 : _GEN11148;
wire  _GEN11154 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11155 = io_x[41] ? _GEN6836 : _GEN11154;
wire  _GEN11156 = io_x[14] ? _GEN11155 : _GEN6843;
wire  _GEN11157 = io_x[0] ? _GEN11156 : _GEN6845;
wire  _GEN11158 = io_x[76] ? _GEN6834 : _GEN11157;
wire  _GEN11159 = io_x[42] ? _GEN11158 : _GEN11153;
wire  _GEN11160 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11161 = io_x[41] ? _GEN11160 : _GEN6836;
wire  _GEN11162 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN11163 = io_x[14] ? _GEN11162 : _GEN11161;
wire  _GEN11164 = io_x[0] ? _GEN11163 : _GEN6845;
wire  _GEN11165 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11166 = io_x[6] ? _GEN11165 : _GEN6850;
wire  _GEN11167 = io_x[41] ? _GEN11166 : _GEN6836;
wire  _GEN11168 = io_x[14] ? _GEN11167 : _GEN6843;
wire  _GEN11169 = io_x[0] ? _GEN11168 : _GEN6845;
wire  _GEN11170 = io_x[76] ? _GEN11169 : _GEN11164;
wire  _GEN11171 = io_x[42] ? _GEN6863 : _GEN11170;
wire  _GEN11172 = io_x[38] ? _GEN11171 : _GEN11159;
wire  _GEN11173 = io_x[10] ? _GEN11172 : _GEN11142;
wire  _GEN11174 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11175 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11176 = io_x[6] ? _GEN11175 : _GEN11174;
wire  _GEN11177 = io_x[41] ? _GEN6836 : _GEN11176;
wire  _GEN11178 = io_x[14] ? _GEN11177 : _GEN6843;
wire  _GEN11179 = io_x[0] ? _GEN11178 : _GEN6845;
wire  _GEN11180 = io_x[76] ? _GEN6834 : _GEN11179;
wire  _GEN11181 = io_x[42] ? _GEN6874 : _GEN11180;
wire  _GEN11182 = io_x[38] ? _GEN11181 : _GEN6871;
wire  _GEN11183 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11184 = io_x[6] ? _GEN11183 : _GEN6840;
wire  _GEN11185 = io_x[41] ? _GEN6836 : _GEN11184;
wire  _GEN11186 = io_x[14] ? _GEN11185 : _GEN6856;
wire  _GEN11187 = io_x[0] ? _GEN11186 : _GEN6845;
wire  _GEN11188 = io_x[76] ? _GEN6834 : _GEN11187;
wire  _GEN11189 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11190 = io_x[41] ? _GEN6836 : _GEN11189;
wire  _GEN11191 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11192 = io_x[41] ? _GEN6924 : _GEN11191;
wire  _GEN11193 = io_x[14] ? _GEN11192 : _GEN11190;
wire  _GEN11194 = io_x[0] ? _GEN11193 : _GEN6845;
wire  _GEN11195 = io_x[76] ? _GEN6834 : _GEN11194;
wire  _GEN11196 = io_x[42] ? _GEN11195 : _GEN11188;
wire  _GEN11197 = io_x[38] ? _GEN11196 : _GEN6871;
wire  _GEN11198 = io_x[10] ? _GEN11197 : _GEN11182;
wire  _GEN11199 = io_x[71] ? _GEN11198 : _GEN11173;
wire  _GEN11200 = io_x[70] ? _GEN11199 : _GEN11132;
wire  _GEN11201 = io_x[33] ? _GEN11200 : _GEN11081;
wire  _GEN11202 = io_x[21] ? _GEN11201 : _GEN10698;
wire  _GEN11203 = io_x[18] ? _GEN11202 : _GEN10426;
wire  _GEN11204 = io_x[20] ? _GEN11203 : _GEN10054;
wire  _GEN11205 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11206 = io_x[0] ? _GEN6845 : _GEN11205;
wire  _GEN11207 = io_x[76] ? _GEN6834 : _GEN11206;
wire  _GEN11208 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN11209 = io_x[76] ? _GEN6834 : _GEN11208;
wire  _GEN11210 = io_x[42] ? _GEN11209 : _GEN11207;
wire  _GEN11211 = io_x[38] ? _GEN11210 : _GEN7036;
wire  _GEN11212 = io_x[10] ? _GEN7044 : _GEN11211;
wire  _GEN11213 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11214 = io_x[0] ? _GEN11213 : _GEN6845;
wire  _GEN11215 = io_x[76] ? _GEN11214 : _GEN6833;
wire  _GEN11216 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN11217 = io_x[76] ? _GEN11216 : _GEN6834;
wire  _GEN11218 = io_x[42] ? _GEN11217 : _GEN11215;
wire  _GEN11219 = io_x[38] ? _GEN11218 : _GEN6871;
wire  _GEN11220 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN11221 = io_x[42] ? _GEN11220 : _GEN6863;
wire  _GEN11222 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11223 = io_x[0] ? _GEN11222 : _GEN6845;
wire  _GEN11224 = io_x[76] ? _GEN6834 : _GEN11223;
wire  _GEN11225 = io_x[42] ? _GEN6874 : _GEN11224;
wire  _GEN11226 = io_x[38] ? _GEN11225 : _GEN11221;
wire  _GEN11227 = io_x[10] ? _GEN11226 : _GEN11219;
wire  _GEN11228 = io_x[71] ? _GEN11227 : _GEN11212;
wire  _GEN11229 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11230 = io_x[2] ? _GEN6837 : _GEN11229;
wire  _GEN11231 = io_x[6] ? _GEN6850 : _GEN11230;
wire  _GEN11232 = io_x[41] ? _GEN6836 : _GEN11231;
wire  _GEN11233 = io_x[14] ? _GEN6843 : _GEN11232;
wire  _GEN11234 = io_x[0] ? _GEN6845 : _GEN11233;
wire  _GEN11235 = io_x[76] ? _GEN11234 : _GEN6834;
wire  _GEN11236 = io_x[42] ? _GEN11235 : _GEN6863;
wire  _GEN11237 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN11238 = io_x[42] ? _GEN6874 : _GEN11237;
wire  _GEN11239 = io_x[38] ? _GEN11238 : _GEN11236;
wire  _GEN11240 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11241 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN11242 = io_x[14] ? _GEN11241 : _GEN6843;
wire  _GEN11243 = io_x[0] ? _GEN11242 : _GEN11240;
wire  _GEN11244 = io_x[76] ? _GEN6834 : _GEN11243;
wire  _GEN11245 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11246 = io_x[0] ? _GEN6845 : _GEN11245;
wire  _GEN11247 = io_x[76] ? _GEN6834 : _GEN11246;
wire  _GEN11248 = io_x[42] ? _GEN11247 : _GEN11244;
wire  _GEN11249 = io_x[38] ? _GEN6871 : _GEN11248;
wire  _GEN11250 = io_x[10] ? _GEN11249 : _GEN11239;
wire  _GEN11251 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN11252 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN11253 = io_x[38] ? _GEN11252 : _GEN11251;
wire  _GEN11254 = io_x[10] ? _GEN7094 : _GEN11253;
wire  _GEN11255 = io_x[71] ? _GEN11254 : _GEN11250;
wire  _GEN11256 = io_x[70] ? _GEN11255 : _GEN11228;
wire  _GEN11257 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11258 = io_x[41] ? _GEN6836 : _GEN11257;
wire  _GEN11259 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11260 = io_x[41] ? _GEN6836 : _GEN11259;
wire  _GEN11261 = io_x[14] ? _GEN11260 : _GEN11258;
wire  _GEN11262 = io_x[0] ? _GEN6845 : _GEN11261;
wire  _GEN11263 = io_x[76] ? _GEN11262 : _GEN6834;
wire  _GEN11264 = io_x[42] ? _GEN11263 : _GEN6874;
wire  _GEN11265 = io_x[38] ? _GEN6871 : _GEN11264;
wire  _GEN11266 = io_x[10] ? _GEN11265 : _GEN7094;
wire  _GEN11267 = io_x[71] ? _GEN11266 : _GEN7196;
wire  _GEN11268 = io_x[70] ? _GEN8474 : _GEN11267;
wire  _GEN11269 = io_x[33] ? _GEN11268 : _GEN11256;
wire  _GEN11270 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11271 = io_x[6] ? _GEN11270 : _GEN6850;
wire  _GEN11272 = io_x[41] ? _GEN6836 : _GEN11271;
wire  _GEN11273 = io_x[14] ? _GEN11272 : _GEN6843;
wire  _GEN11274 = io_x[0] ? _GEN6845 : _GEN11273;
wire  _GEN11275 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11276 = io_x[14] ? _GEN11275 : _GEN6843;
wire  _GEN11277 = io_x[0] ? _GEN11276 : _GEN6845;
wire  _GEN11278 = io_x[76] ? _GEN11277 : _GEN11274;
wire  _GEN11279 = io_x[42] ? _GEN6874 : _GEN11278;
wire  _GEN11280 = io_x[38] ? _GEN11279 : _GEN6871;
wire  _GEN11281 = io_x[10] ? _GEN11280 : _GEN7094;
wire  _GEN11282 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN11283 = io_x[42] ? _GEN6874 : _GEN11282;
wire  _GEN11284 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN11285 = io_x[76] ? _GEN11284 : _GEN6834;
wire  _GEN11286 = io_x[42] ? _GEN11285 : _GEN6863;
wire  _GEN11287 = io_x[38] ? _GEN11286 : _GEN11283;
wire  _GEN11288 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11289 = io_x[14] ? _GEN11288 : _GEN6856;
wire  _GEN11290 = io_x[0] ? _GEN11289 : _GEN6845;
wire  _GEN11291 = io_x[76] ? _GEN11290 : _GEN6834;
wire  _GEN11292 = io_x[42] ? _GEN11291 : _GEN6874;
wire  _GEN11293 = io_x[38] ? _GEN11292 : _GEN6871;
wire  _GEN11294 = io_x[10] ? _GEN11293 : _GEN11287;
wire  _GEN11295 = io_x[71] ? _GEN11294 : _GEN11281;
wire  _GEN11296 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11297 = io_x[0] ? _GEN6845 : _GEN11296;
wire  _GEN11298 = io_x[76] ? _GEN11297 : _GEN6834;
wire  _GEN11299 = io_x[42] ? _GEN11298 : _GEN6863;
wire  _GEN11300 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN11301 = io_x[42] ? _GEN11300 : _GEN6863;
wire  _GEN11302 = io_x[38] ? _GEN11301 : _GEN11299;
wire  _GEN11303 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11304 = io_x[14] ? _GEN11303 : _GEN6843;
wire  _GEN11305 = io_x[0] ? _GEN11304 : _GEN6845;
wire  _GEN11306 = io_x[76] ? _GEN6833 : _GEN11305;
wire  _GEN11307 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11308 = io_x[0] ? _GEN11307 : _GEN6845;
wire  _GEN11309 = io_x[76] ? _GEN11308 : _GEN6833;
wire  _GEN11310 = io_x[42] ? _GEN11309 : _GEN11306;
wire  _GEN11311 = io_x[38] ? _GEN7036 : _GEN11310;
wire  _GEN11312 = io_x[10] ? _GEN11311 : _GEN11302;
wire  _GEN11313 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11314 = io_x[2] ? _GEN6837 : _GEN11313;
wire  _GEN11315 = io_x[6] ? _GEN6850 : _GEN11314;
wire  _GEN11316 = io_x[41] ? _GEN6836 : _GEN11315;
wire  _GEN11317 = io_x[14] ? _GEN6843 : _GEN11316;
wire  _GEN11318 = io_x[0] ? _GEN6845 : _GEN11317;
wire  _GEN11319 = io_x[76] ? _GEN11318 : _GEN6834;
wire  _GEN11320 = io_x[42] ? _GEN6874 : _GEN11319;
wire  _GEN11321 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11322 = io_x[41] ? _GEN6836 : _GEN11321;
wire  _GEN11323 = io_x[14] ? _GEN6843 : _GEN11322;
wire  _GEN11324 = io_x[0] ? _GEN6845 : _GEN11323;
wire  _GEN11325 = io_x[76] ? _GEN11324 : _GEN6834;
wire  _GEN11326 = io_x[42] ? _GEN11325 : _GEN6874;
wire  _GEN11327 = io_x[38] ? _GEN11326 : _GEN11320;
wire  _GEN11328 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN11329 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN11330 = io_x[42] ? _GEN11329 : _GEN11328;
wire  _GEN11331 = io_x[38] ? _GEN11330 : _GEN6871;
wire  _GEN11332 = io_x[10] ? _GEN11331 : _GEN11327;
wire  _GEN11333 = io_x[71] ? _GEN11332 : _GEN11312;
wire  _GEN11334 = io_x[70] ? _GEN11333 : _GEN11295;
wire  _GEN11335 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11336 = io_x[41] ? _GEN6836 : _GEN11335;
wire  _GEN11337 = io_x[14] ? _GEN6843 : _GEN11336;
wire  _GEN11338 = io_x[0] ? _GEN6845 : _GEN11337;
wire  _GEN11339 = io_x[76] ? _GEN11338 : _GEN6834;
wire  _GEN11340 = io_x[42] ? _GEN11339 : _GEN6874;
wire  _GEN11341 = io_x[38] ? _GEN11340 : _GEN6871;
wire  _GEN11342 = io_x[10] ? _GEN7044 : _GEN11341;
wire  _GEN11343 = io_x[71] ? _GEN11342 : _GEN7196;
wire  _GEN11344 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11345 = io_x[0] ? _GEN11344 : _GEN6845;
wire  _GEN11346 = io_x[76] ? _GEN11345 : _GEN6834;
wire  _GEN11347 = io_x[42] ? _GEN6874 : _GEN11346;
wire  _GEN11348 = io_x[38] ? _GEN11347 : _GEN6871;
wire  _GEN11349 = io_x[10] ? _GEN11348 : _GEN7044;
wire  _GEN11350 = io_x[71] ? _GEN11349 : _GEN7196;
wire  _GEN11351 = io_x[70] ? _GEN11350 : _GEN11343;
wire  _GEN11352 = io_x[33] ? _GEN11351 : _GEN11334;
wire  _GEN11353 = io_x[21] ? _GEN11352 : _GEN11269;
wire  _GEN11354 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN11355 = io_x[76] ? _GEN6833 : _GEN11354;
wire  _GEN11356 = io_x[42] ? _GEN6863 : _GEN11355;
wire  _GEN11357 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN11358 = io_x[38] ? _GEN11357 : _GEN11356;
wire  _GEN11359 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11360 = io_x[41] ? _GEN6836 : _GEN11359;
wire  _GEN11361 = io_x[14] ? _GEN11360 : _GEN6843;
wire  _GEN11362 = io_x[0] ? _GEN11361 : _GEN6858;
wire  _GEN11363 = io_x[76] ? _GEN6834 : _GEN11362;
wire  _GEN11364 = io_x[42] ? _GEN6874 : _GEN11363;
wire  _GEN11365 = io_x[38] ? _GEN7036 : _GEN11364;
wire  _GEN11366 = io_x[10] ? _GEN11365 : _GEN11358;
wire  _GEN11367 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11368 = io_x[0] ? _GEN6845 : _GEN11367;
wire  _GEN11369 = io_x[76] ? _GEN6834 : _GEN11368;
wire  _GEN11370 = io_x[42] ? _GEN11369 : _GEN6874;
wire  _GEN11371 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11372 = io_x[6] ? _GEN6840 : _GEN11371;
wire  _GEN11373 = io_x[41] ? _GEN11372 : _GEN6836;
wire  _GEN11374 = io_x[14] ? _GEN6856 : _GEN11373;
wire  _GEN11375 = io_x[0] ? _GEN6845 : _GEN11374;
wire  _GEN11376 = io_x[76] ? _GEN11375 : _GEN6833;
wire  _GEN11377 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11378 = io_x[6] ? _GEN11377 : _GEN6840;
wire  _GEN11379 = io_x[41] ? _GEN6836 : _GEN11378;
wire  _GEN11380 = io_x[14] ? _GEN11379 : _GEN6856;
wire  _GEN11381 = io_x[0] ? _GEN6845 : _GEN11380;
wire  _GEN11382 = io_x[76] ? _GEN11381 : _GEN6834;
wire  _GEN11383 = io_x[42] ? _GEN11382 : _GEN11376;
wire  _GEN11384 = io_x[38] ? _GEN11383 : _GEN11370;
wire  _GEN11385 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN11386 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11387 = io_x[6] ? _GEN11386 : _GEN6840;
wire  _GEN11388 = io_x[41] ? _GEN11387 : _GEN6836;
wire  _GEN11389 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11390 = io_x[6] ? _GEN11389 : _GEN6850;
wire  _GEN11391 = io_x[41] ? _GEN11390 : _GEN6836;
wire  _GEN11392 = io_x[14] ? _GEN11391 : _GEN11388;
wire  _GEN11393 = io_x[0] ? _GEN6845 : _GEN11392;
wire  _GEN11394 = io_x[76] ? _GEN11393 : _GEN11385;
wire  _GEN11395 = io_x[42] ? _GEN6874 : _GEN11394;
wire  _GEN11396 = io_x[38] ? _GEN11395 : _GEN6871;
wire  _GEN11397 = io_x[10] ? _GEN11396 : _GEN11384;
wire  _GEN11398 = io_x[71] ? _GEN11397 : _GEN11366;
wire  _GEN11399 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11400 = io_x[0] ? _GEN11399 : _GEN6858;
wire  _GEN11401 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11402 = io_x[41] ? _GEN11401 : _GEN6836;
wire  _GEN11403 = io_x[14] ? _GEN11402 : _GEN6843;
wire  _GEN11404 = io_x[0] ? _GEN11403 : _GEN6858;
wire  _GEN11405 = io_x[76] ? _GEN11404 : _GEN11400;
wire  _GEN11406 = io_x[42] ? _GEN6874 : _GEN11405;
wire  _GEN11407 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11408 = io_x[6] ? _GEN11407 : _GEN6850;
wire  _GEN11409 = io_x[41] ? _GEN11408 : _GEN6836;
wire  _GEN11410 = io_x[14] ? _GEN6843 : _GEN11409;
wire  _GEN11411 = io_x[0] ? _GEN6845 : _GEN11410;
wire  _GEN11412 = io_x[76] ? _GEN6834 : _GEN11411;
wire  _GEN11413 = io_x[42] ? _GEN6863 : _GEN11412;
wire  _GEN11414 = io_x[38] ? _GEN11413 : _GEN11406;
wire  _GEN11415 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11416 = io_x[14] ? _GEN11415 : _GEN6843;
wire  _GEN11417 = io_x[0] ? _GEN11416 : _GEN6845;
wire  _GEN11418 = io_x[76] ? _GEN6834 : _GEN11417;
wire  _GEN11419 = io_x[42] ? _GEN6863 : _GEN11418;
wire  _GEN11420 = io_x[38] ? _GEN6871 : _GEN11419;
wire  _GEN11421 = io_x[10] ? _GEN11420 : _GEN11414;
wire  _GEN11422 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11423 = io_x[0] ? _GEN6845 : _GEN11422;
wire  _GEN11424 = io_x[76] ? _GEN6833 : _GEN11423;
wire  _GEN11425 = io_x[42] ? _GEN6863 : _GEN11424;
wire  _GEN11426 = io_x[38] ? _GEN11425 : _GEN6871;
wire  _GEN11427 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11428 = io_x[41] ? _GEN11427 : _GEN6836;
wire  _GEN11429 = io_x[14] ? _GEN11428 : _GEN6843;
wire  _GEN11430 = io_x[0] ? _GEN6845 : _GEN11429;
wire  _GEN11431 = io_x[76] ? _GEN6834 : _GEN11430;
wire  _GEN11432 = io_x[42] ? _GEN6874 : _GEN11431;
wire  _GEN11433 = io_x[38] ? _GEN11432 : _GEN6871;
wire  _GEN11434 = io_x[10] ? _GEN11433 : _GEN11426;
wire  _GEN11435 = io_x[71] ? _GEN11434 : _GEN11421;
wire  _GEN11436 = io_x[70] ? _GEN11435 : _GEN11398;
wire  _GEN11437 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN11438 = io_x[42] ? _GEN6863 : _GEN11437;
wire  _GEN11439 = io_x[38] ? _GEN6871 : _GEN11438;
wire  _GEN11440 = io_x[10] ? _GEN7044 : _GEN11439;
wire  _GEN11441 = io_x[71] ? _GEN11440 : _GEN7196;
wire  _GEN11442 = io_x[70] ? _GEN11441 : _GEN7020;
wire  _GEN11443 = io_x[33] ? _GEN11442 : _GEN11436;
wire  _GEN11444 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11445 = io_x[2] ? _GEN6837 : _GEN11444;
wire  _GEN11446 = io_x[6] ? _GEN6850 : _GEN11445;
wire  _GEN11447 = io_x[41] ? _GEN11446 : _GEN6836;
wire  _GEN11448 = io_x[14] ? _GEN6843 : _GEN11447;
wire  _GEN11449 = io_x[0] ? _GEN6845 : _GEN11448;
wire  _GEN11450 = io_x[76] ? _GEN6834 : _GEN11449;
wire  _GEN11451 = io_x[42] ? _GEN11450 : _GEN6874;
wire  _GEN11452 = io_x[38] ? _GEN11451 : _GEN7036;
wire  _GEN11453 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11454 = io_x[41] ? _GEN6836 : _GEN11453;
wire  _GEN11455 = io_x[14] ? _GEN11454 : _GEN6856;
wire  _GEN11456 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11457 = io_x[6] ? _GEN11456 : _GEN6850;
wire  _GEN11458 = io_x[41] ? _GEN6836 : _GEN11457;
wire  _GEN11459 = io_x[14] ? _GEN11458 : _GEN6856;
wire  _GEN11460 = io_x[0] ? _GEN11459 : _GEN11455;
wire  _GEN11461 = io_x[76] ? _GEN6834 : _GEN11460;
wire  _GEN11462 = io_x[42] ? _GEN6874 : _GEN11461;
wire  _GEN11463 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN11464 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11465 = io_x[14] ? _GEN11464 : _GEN11463;
wire  _GEN11466 = io_x[0] ? _GEN11465 : _GEN6845;
wire  _GEN11467 = io_x[76] ? _GEN11466 : _GEN6834;
wire  _GEN11468 = io_x[42] ? _GEN6874 : _GEN11467;
wire  _GEN11469 = io_x[38] ? _GEN11468 : _GEN11462;
wire  _GEN11470 = io_x[10] ? _GEN11469 : _GEN11452;
wire  _GEN11471 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11472 = io_x[6] ? _GEN11471 : _GEN6850;
wire  _GEN11473 = io_x[41] ? _GEN11472 : _GEN6836;
wire  _GEN11474 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11475 = io_x[41] ? _GEN11474 : _GEN6836;
wire  _GEN11476 = io_x[14] ? _GEN11475 : _GEN11473;
wire  _GEN11477 = io_x[0] ? _GEN6845 : _GEN11476;
wire  _GEN11478 = io_x[76] ? _GEN11477 : _GEN6833;
wire  _GEN11479 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11480 = io_x[0] ? _GEN6845 : _GEN11479;
wire  _GEN11481 = io_x[76] ? _GEN11480 : _GEN6834;
wire  _GEN11482 = io_x[42] ? _GEN11481 : _GEN11478;
wire  _GEN11483 = io_x[38] ? _GEN11482 : _GEN6871;
wire  _GEN11484 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN11485 = io_x[42] ? _GEN6874 : _GEN11484;
wire  _GEN11486 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11487 = io_x[6] ? _GEN6850 : _GEN11486;
wire  _GEN11488 = io_x[41] ? _GEN11487 : _GEN6836;
wire  _GEN11489 = io_x[14] ? _GEN11488 : _GEN6843;
wire  _GEN11490 = io_x[0] ? _GEN6845 : _GEN11489;
wire  _GEN11491 = io_x[76] ? _GEN11490 : _GEN6833;
wire  _GEN11492 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11493 = io_x[0] ? _GEN11492 : _GEN6858;
wire  _GEN11494 = io_x[76] ? _GEN11493 : _GEN6834;
wire  _GEN11495 = io_x[42] ? _GEN11494 : _GEN11491;
wire  _GEN11496 = io_x[38] ? _GEN11495 : _GEN11485;
wire  _GEN11497 = io_x[10] ? _GEN11496 : _GEN11483;
wire  _GEN11498 = io_x[71] ? _GEN11497 : _GEN11470;
wire  _GEN11499 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN11500 = io_x[38] ? _GEN11499 : _GEN7036;
wire  _GEN11501 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11502 = io_x[6] ? _GEN11501 : _GEN6850;
wire  _GEN11503 = io_x[41] ? _GEN11502 : _GEN6836;
wire  _GEN11504 = io_x[14] ? _GEN11503 : _GEN6856;
wire  _GEN11505 = io_x[0] ? _GEN11504 : _GEN6845;
wire  _GEN11506 = io_x[76] ? _GEN6834 : _GEN11505;
wire  _GEN11507 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11508 = io_x[2] ? _GEN11507 : _GEN6837;
wire  _GEN11509 = io_x[6] ? _GEN11508 : _GEN6850;
wire  _GEN11510 = io_x[41] ? _GEN11509 : _GEN6836;
wire  _GEN11511 = io_x[14] ? _GEN11510 : _GEN6843;
wire  _GEN11512 = io_x[0] ? _GEN11511 : _GEN6845;
wire  _GEN11513 = io_x[76] ? _GEN11512 : _GEN6834;
wire  _GEN11514 = io_x[42] ? _GEN11513 : _GEN11506;
wire  _GEN11515 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11516 = io_x[2] ? _GEN11515 : _GEN6837;
wire  _GEN11517 = io_x[6] ? _GEN11516 : _GEN6850;
wire  _GEN11518 = io_x[41] ? _GEN6836 : _GEN11517;
wire  _GEN11519 = io_x[14] ? _GEN11518 : _GEN6856;
wire  _GEN11520 = io_x[0] ? _GEN11519 : _GEN6845;
wire  _GEN11521 = io_x[76] ? _GEN11520 : _GEN6834;
wire  _GEN11522 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN11523 = io_x[76] ? _GEN11522 : _GEN6833;
wire  _GEN11524 = io_x[42] ? _GEN11523 : _GEN11521;
wire  _GEN11525 = io_x[38] ? _GEN11524 : _GEN11514;
wire  _GEN11526 = io_x[10] ? _GEN11525 : _GEN11500;
wire  _GEN11527 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11528 = io_x[2] ? _GEN6837 : _GEN11527;
wire  _GEN11529 = io_x[6] ? _GEN6850 : _GEN11528;
wire  _GEN11530 = io_x[41] ? _GEN6836 : _GEN11529;
wire  _GEN11531 = io_x[14] ? _GEN6843 : _GEN11530;
wire  _GEN11532 = io_x[0] ? _GEN6845 : _GEN11531;
wire  _GEN11533 = io_x[76] ? _GEN11532 : _GEN6834;
wire  _GEN11534 = io_x[42] ? _GEN6874 : _GEN11533;
wire  _GEN11535 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN11536 = io_x[76] ? _GEN11535 : _GEN6834;
wire  _GEN11537 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11538 = io_x[0] ? _GEN6845 : _GEN11537;
wire  _GEN11539 = io_x[76] ? _GEN11538 : _GEN6834;
wire  _GEN11540 = io_x[42] ? _GEN11539 : _GEN11536;
wire  _GEN11541 = io_x[38] ? _GEN11540 : _GEN11534;
wire  _GEN11542 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11543 = io_x[6] ? _GEN11542 : _GEN6850;
wire  _GEN11544 = io_x[41] ? _GEN6924 : _GEN11543;
wire  _GEN11545 = io_x[14] ? _GEN11544 : _GEN6843;
wire  _GEN11546 = io_x[0] ? _GEN11545 : _GEN6845;
wire  _GEN11547 = io_x[76] ? _GEN6834 : _GEN11546;
wire  _GEN11548 = io_x[42] ? _GEN6874 : _GEN11547;
wire  _GEN11549 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN11550 = io_x[14] ? _GEN6843 : _GEN11549;
wire  _GEN11551 = io_x[0] ? _GEN11550 : _GEN6858;
wire  _GEN11552 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11553 = io_x[0] ? _GEN11552 : _GEN6845;
wire  _GEN11554 = io_x[76] ? _GEN11553 : _GEN11551;
wire  _GEN11555 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN11556 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11557 = io_x[41] ? _GEN6836 : _GEN11556;
wire  _GEN11558 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11559 = io_x[41] ? _GEN6924 : _GEN11558;
wire  _GEN11560 = io_x[14] ? _GEN11559 : _GEN11557;
wire  _GEN11561 = io_x[0] ? _GEN6845 : _GEN11560;
wire  _GEN11562 = io_x[76] ? _GEN11561 : _GEN11555;
wire  _GEN11563 = io_x[42] ? _GEN11562 : _GEN11554;
wire  _GEN11564 = io_x[38] ? _GEN11563 : _GEN11548;
wire  _GEN11565 = io_x[10] ? _GEN11564 : _GEN11541;
wire  _GEN11566 = io_x[71] ? _GEN11565 : _GEN11526;
wire  _GEN11567 = io_x[70] ? _GEN11566 : _GEN11498;
wire  _GEN11568 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11569 = io_x[41] ? _GEN6836 : _GEN11568;
wire  _GEN11570 = io_x[14] ? _GEN11569 : _GEN6843;
wire  _GEN11571 = io_x[0] ? _GEN11570 : _GEN6845;
wire  _GEN11572 = io_x[76] ? _GEN11571 : _GEN6834;
wire  _GEN11573 = io_x[42] ? _GEN6874 : _GEN11572;
wire  _GEN11574 = io_x[38] ? _GEN7036 : _GEN11573;
wire  _GEN11575 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11576 = io_x[41] ? _GEN6836 : _GEN11575;
wire  _GEN11577 = io_x[14] ? _GEN11576 : _GEN6843;
wire  _GEN11578 = io_x[0] ? _GEN11577 : _GEN6845;
wire  _GEN11579 = io_x[76] ? _GEN11578 : _GEN6834;
wire  _GEN11580 = io_x[42] ? _GEN6874 : _GEN11579;
wire  _GEN11581 = io_x[38] ? _GEN6871 : _GEN11580;
wire  _GEN11582 = io_x[10] ? _GEN11581 : _GEN11574;
wire  _GEN11583 = io_x[71] ? _GEN11582 : _GEN7203;
wire  _GEN11584 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN11585 = io_x[42] ? _GEN6874 : _GEN11584;
wire  _GEN11586 = io_x[38] ? _GEN6871 : _GEN11585;
wire  _GEN11587 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN11588 = io_x[38] ? _GEN11587 : _GEN6871;
wire  _GEN11589 = io_x[10] ? _GEN11588 : _GEN11586;
wire  _GEN11590 = io_x[71] ? _GEN11589 : _GEN7203;
wire  _GEN11591 = io_x[70] ? _GEN11590 : _GEN11583;
wire  _GEN11592 = io_x[33] ? _GEN11591 : _GEN11567;
wire  _GEN11593 = io_x[21] ? _GEN11592 : _GEN11443;
wire  _GEN11594 = io_x[18] ? _GEN11593 : _GEN11353;
wire  _GEN11595 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11596 = io_x[6] ? _GEN11595 : _GEN6850;
wire  _GEN11597 = io_x[41] ? _GEN6836 : _GEN11596;
wire  _GEN11598 = io_x[14] ? _GEN11597 : _GEN6843;
wire  _GEN11599 = io_x[0] ? _GEN11598 : _GEN6845;
wire  _GEN11600 = io_x[76] ? _GEN6834 : _GEN11599;
wire  _GEN11601 = io_x[42] ? _GEN6874 : _GEN11600;
wire  _GEN11602 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN11603 = io_x[76] ? _GEN6834 : _GEN11602;
wire  _GEN11604 = io_x[42] ? _GEN11603 : _GEN6874;
wire  _GEN11605 = io_x[38] ? _GEN11604 : _GEN11601;
wire  _GEN11606 = io_x[10] ? _GEN11605 : _GEN7094;
wire  _GEN11607 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN11608 = io_x[76] ? _GEN11607 : _GEN6834;
wire  _GEN11609 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11610 = io_x[41] ? _GEN6836 : _GEN11609;
wire  _GEN11611 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11612 = io_x[41] ? _GEN6836 : _GEN11611;
wire  _GEN11613 = io_x[14] ? _GEN11612 : _GEN11610;
wire  _GEN11614 = io_x[0] ? _GEN6845 : _GEN11613;
wire  _GEN11615 = io_x[76] ? _GEN11614 : _GEN6834;
wire  _GEN11616 = io_x[42] ? _GEN11615 : _GEN11608;
wire  _GEN11617 = io_x[38] ? _GEN11616 : _GEN6871;
wire  _GEN11618 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN11619 = io_x[10] ? _GEN11618 : _GEN11617;
wire  _GEN11620 = io_x[71] ? _GEN11619 : _GEN11606;
wire  _GEN11621 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN11622 = io_x[42] ? _GEN6874 : _GEN11621;
wire  _GEN11623 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11624 = io_x[41] ? _GEN6836 : _GEN11623;
wire  _GEN11625 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11626 = io_x[41] ? _GEN6836 : _GEN11625;
wire  _GEN11627 = io_x[14] ? _GEN11626 : _GEN11624;
wire  _GEN11628 = io_x[0] ? _GEN6845 : _GEN11627;
wire  _GEN11629 = io_x[76] ? _GEN11628 : _GEN6833;
wire  _GEN11630 = io_x[42] ? _GEN11629 : _GEN6863;
wire  _GEN11631 = io_x[38] ? _GEN11630 : _GEN11622;
wire  _GEN11632 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN11633 = io_x[76] ? _GEN6834 : _GEN11632;
wire  _GEN11634 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN11635 = io_x[42] ? _GEN11634 : _GEN11633;
wire  _GEN11636 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11637 = io_x[6] ? _GEN11636 : _GEN6850;
wire  _GEN11638 = io_x[41] ? _GEN6836 : _GEN11637;
wire  _GEN11639 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11640 = io_x[6] ? _GEN11639 : _GEN6850;
wire  _GEN11641 = io_x[41] ? _GEN6836 : _GEN11640;
wire  _GEN11642 = io_x[14] ? _GEN11641 : _GEN11638;
wire  _GEN11643 = io_x[0] ? _GEN11642 : _GEN6845;
wire  _GEN11644 = io_x[76] ? _GEN6833 : _GEN11643;
wire  _GEN11645 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11646 = io_x[41] ? _GEN6836 : _GEN11645;
wire  _GEN11647 = io_x[14] ? _GEN6856 : _GEN11646;
wire  _GEN11648 = io_x[0] ? _GEN6845 : _GEN11647;
wire  _GEN11649 = io_x[76] ? _GEN11648 : _GEN6834;
wire  _GEN11650 = io_x[42] ? _GEN11649 : _GEN11644;
wire  _GEN11651 = io_x[38] ? _GEN11650 : _GEN11635;
wire  _GEN11652 = io_x[10] ? _GEN11651 : _GEN11631;
wire  _GEN11653 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11654 = io_x[0] ? _GEN6845 : _GEN11653;
wire  _GEN11655 = io_x[76] ? _GEN11654 : _GEN6834;
wire  _GEN11656 = io_x[42] ? _GEN11655 : _GEN6874;
wire  _GEN11657 = io_x[38] ? _GEN11656 : _GEN6871;
wire  _GEN11658 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN11659 = io_x[42] ? _GEN11658 : _GEN6874;
wire  _GEN11660 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11661 = io_x[0] ? _GEN6845 : _GEN11660;
wire  _GEN11662 = io_x[76] ? _GEN11661 : _GEN6834;
wire  _GEN11663 = io_x[42] ? _GEN11662 : _GEN6874;
wire  _GEN11664 = io_x[38] ? _GEN11663 : _GEN11659;
wire  _GEN11665 = io_x[10] ? _GEN11664 : _GEN11657;
wire  _GEN11666 = io_x[71] ? _GEN11665 : _GEN11652;
wire  _GEN11667 = io_x[70] ? _GEN11666 : _GEN11620;
wire  _GEN11668 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11669 = io_x[41] ? _GEN6836 : _GEN11668;
wire  _GEN11670 = io_x[14] ? _GEN6843 : _GEN11669;
wire  _GEN11671 = io_x[0] ? _GEN6845 : _GEN11670;
wire  _GEN11672 = io_x[76] ? _GEN11671 : _GEN6834;
wire  _GEN11673 = io_x[42] ? _GEN11672 : _GEN6874;
wire  _GEN11674 = io_x[38] ? _GEN11673 : _GEN6871;
wire  _GEN11675 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN11676 = io_x[10] ? _GEN11675 : _GEN11674;
wire  _GEN11677 = io_x[71] ? _GEN11676 : _GEN7196;
wire  _GEN11678 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN11679 = io_x[71] ? _GEN11678 : _GEN7196;
wire  _GEN11680 = io_x[70] ? _GEN11679 : _GEN11677;
wire  _GEN11681 = io_x[33] ? _GEN11680 : _GEN11667;
wire  _GEN11682 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11683 = io_x[0] ? _GEN6845 : _GEN11682;
wire  _GEN11684 = io_x[76] ? _GEN6833 : _GEN11683;
wire  _GEN11685 = io_x[42] ? _GEN6874 : _GEN11684;
wire  _GEN11686 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11687 = io_x[14] ? _GEN6843 : _GEN11686;
wire  _GEN11688 = io_x[0] ? _GEN6845 : _GEN11687;
wire  _GEN11689 = io_x[76] ? _GEN6834 : _GEN11688;
wire  _GEN11690 = io_x[42] ? _GEN11689 : _GEN6874;
wire  _GEN11691 = io_x[38] ? _GEN11690 : _GEN11685;
wire  _GEN11692 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN11693 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11694 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11695 = io_x[0] ? _GEN11694 : _GEN11693;
wire  _GEN11696 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11697 = io_x[14] ? _GEN11696 : _GEN6843;
wire  _GEN11698 = io_x[0] ? _GEN11697 : _GEN6845;
wire  _GEN11699 = io_x[76] ? _GEN11698 : _GEN11695;
wire  _GEN11700 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN11701 = io_x[76] ? _GEN6834 : _GEN11700;
wire  _GEN11702 = io_x[42] ? _GEN11701 : _GEN11699;
wire  _GEN11703 = io_x[38] ? _GEN11702 : _GEN11692;
wire  _GEN11704 = io_x[10] ? _GEN11703 : _GEN11691;
wire  _GEN11705 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11706 = io_x[14] ? _GEN6843 : _GEN11705;
wire  _GEN11707 = io_x[0] ? _GEN6845 : _GEN11706;
wire  _GEN11708 = io_x[76] ? _GEN6834 : _GEN11707;
wire  _GEN11709 = io_x[42] ? _GEN6874 : _GEN11708;
wire  _GEN11710 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN11711 = io_x[38] ? _GEN11710 : _GEN11709;
wire  _GEN11712 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11713 = io_x[6] ? _GEN11712 : _GEN6850;
wire  _GEN11714 = io_x[41] ? _GEN6836 : _GEN11713;
wire  _GEN11715 = io_x[14] ? _GEN11714 : _GEN6843;
wire  _GEN11716 = io_x[0] ? _GEN11715 : _GEN6845;
wire  _GEN11717 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11718 = io_x[0] ? _GEN6845 : _GEN11717;
wire  _GEN11719 = io_x[76] ? _GEN11718 : _GEN11716;
wire  _GEN11720 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11721 = io_x[0] ? _GEN11720 : _GEN6845;
wire  _GEN11722 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11723 = io_x[6] ? _GEN11722 : _GEN6850;
wire  _GEN11724 = io_x[41] ? _GEN6836 : _GEN11723;
wire  _GEN11725 = io_x[14] ? _GEN11724 : _GEN6843;
wire  _GEN11726 = io_x[0] ? _GEN11725 : _GEN6845;
wire  _GEN11727 = io_x[76] ? _GEN11726 : _GEN11721;
wire  _GEN11728 = io_x[42] ? _GEN11727 : _GEN11719;
wire  _GEN11729 = io_x[38] ? _GEN11728 : _GEN7036;
wire  _GEN11730 = io_x[10] ? _GEN11729 : _GEN11711;
wire  _GEN11731 = io_x[71] ? _GEN11730 : _GEN11704;
wire  _GEN11732 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11733 = io_x[2] ? _GEN6837 : _GEN11732;
wire  _GEN11734 = io_x[6] ? _GEN6850 : _GEN11733;
wire  _GEN11735 = io_x[41] ? _GEN6924 : _GEN11734;
wire  _GEN11736 = io_x[14] ? _GEN6843 : _GEN11735;
wire  _GEN11737 = io_x[0] ? _GEN6845 : _GEN11736;
wire  _GEN11738 = io_x[76] ? _GEN11737 : _GEN6833;
wire  _GEN11739 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11740 = io_x[2] ? _GEN6837 : _GEN11739;
wire  _GEN11741 = io_x[6] ? _GEN11740 : _GEN6850;
wire  _GEN11742 = io_x[41] ? _GEN6836 : _GEN11741;
wire  _GEN11743 = io_x[14] ? _GEN11742 : _GEN6843;
wire  _GEN11744 = io_x[0] ? _GEN6858 : _GEN11743;
wire  _GEN11745 = io_x[76] ? _GEN11744 : _GEN6833;
wire  _GEN11746 = io_x[42] ? _GEN11745 : _GEN11738;
wire  _GEN11747 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11748 = io_x[14] ? _GEN6843 : _GEN11747;
wire  _GEN11749 = io_x[0] ? _GEN6845 : _GEN11748;
wire  _GEN11750 = io_x[76] ? _GEN11749 : _GEN6834;
wire  _GEN11751 = io_x[42] ? _GEN6874 : _GEN11750;
wire  _GEN11752 = io_x[38] ? _GEN11751 : _GEN11746;
wire  _GEN11753 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11754 = io_x[2] ? _GEN11753 : _GEN6837;
wire  _GEN11755 = io_x[6] ? _GEN11754 : _GEN6840;
wire  _GEN11756 = io_x[41] ? _GEN6924 : _GEN11755;
wire  _GEN11757 = io_x[14] ? _GEN11756 : _GEN6843;
wire  _GEN11758 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11759 = io_x[6] ? _GEN11758 : _GEN6840;
wire  _GEN11760 = io_x[41] ? _GEN11759 : _GEN6836;
wire  _GEN11761 = io_x[14] ? _GEN11760 : _GEN6843;
wire  _GEN11762 = io_x[0] ? _GEN11761 : _GEN11757;
wire  _GEN11763 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11764 = io_x[6] ? _GEN11763 : _GEN6850;
wire  _GEN11765 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11766 = io_x[6] ? _GEN11765 : _GEN6850;
wire  _GEN11767 = io_x[41] ? _GEN11766 : _GEN11764;
wire  _GEN11768 = io_x[14] ? _GEN11767 : _GEN6843;
wire  _GEN11769 = io_x[0] ? _GEN6858 : _GEN11768;
wire  _GEN11770 = io_x[76] ? _GEN11769 : _GEN11762;
wire  _GEN11771 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11772 = io_x[41] ? _GEN6836 : _GEN11771;
wire  _GEN11773 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN11774 = io_x[2] ? _GEN6837 : _GEN11773;
wire  _GEN11775 = io_x[6] ? _GEN11774 : _GEN6850;
wire  _GEN11776 = io_x[41] ? _GEN6924 : _GEN11775;
wire  _GEN11777 = io_x[14] ? _GEN11776 : _GEN11772;
wire  _GEN11778 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11779 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11780 = io_x[41] ? _GEN6924 : _GEN11779;
wire  _GEN11781 = io_x[14] ? _GEN11780 : _GEN11778;
wire  _GEN11782 = io_x[0] ? _GEN11781 : _GEN11777;
wire  _GEN11783 = io_x[76] ? _GEN11782 : _GEN6833;
wire  _GEN11784 = io_x[42] ? _GEN11783 : _GEN11770;
wire  _GEN11785 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11786 = io_x[0] ? _GEN11785 : _GEN6845;
wire  _GEN11787 = io_x[76] ? _GEN11786 : _GEN6833;
wire  _GEN11788 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11789 = io_x[0] ? _GEN6845 : _GEN11788;
wire  _GEN11790 = io_x[76] ? _GEN11789 : _GEN6833;
wire  _GEN11791 = io_x[42] ? _GEN11790 : _GEN11787;
wire  _GEN11792 = io_x[38] ? _GEN11791 : _GEN11784;
wire  _GEN11793 = io_x[10] ? _GEN11792 : _GEN11752;
wire  _GEN11794 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11795 = io_x[2] ? _GEN6837 : _GEN11794;
wire  _GEN11796 = io_x[6] ? _GEN6850 : _GEN11795;
wire  _GEN11797 = io_x[41] ? _GEN6836 : _GEN11796;
wire  _GEN11798 = io_x[14] ? _GEN6843 : _GEN11797;
wire  _GEN11799 = io_x[0] ? _GEN6845 : _GEN11798;
wire  _GEN11800 = io_x[76] ? _GEN11799 : _GEN6834;
wire  _GEN11801 = io_x[42] ? _GEN6874 : _GEN11800;
wire  _GEN11802 = io_x[38] ? _GEN6871 : _GEN11801;
wire  _GEN11803 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN11804 = io_x[42] ? _GEN6863 : _GEN11803;
wire  _GEN11805 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN11806 = io_x[38] ? _GEN11805 : _GEN11804;
wire  _GEN11807 = io_x[10] ? _GEN11806 : _GEN11802;
wire  _GEN11808 = io_x[71] ? _GEN11807 : _GEN11793;
wire  _GEN11809 = io_x[70] ? _GEN11808 : _GEN11731;
wire  _GEN11810 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11811 = io_x[41] ? _GEN11810 : _GEN6836;
wire  _GEN11812 = io_x[14] ? _GEN11811 : _GEN6843;
wire  _GEN11813 = io_x[0] ? _GEN11812 : _GEN6845;
wire  _GEN11814 = io_x[76] ? _GEN11813 : _GEN6834;
wire  _GEN11815 = io_x[42] ? _GEN11814 : _GEN6863;
wire  _GEN11816 = io_x[38] ? _GEN11815 : _GEN6871;
wire  _GEN11817 = io_x[10] ? _GEN11816 : _GEN7044;
wire  _GEN11818 = io_x[71] ? _GEN11817 : _GEN7196;
wire  _GEN11819 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN11820 = io_x[38] ? _GEN11819 : _GEN6871;
wire  _GEN11821 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11822 = io_x[41] ? _GEN6836 : _GEN11821;
wire  _GEN11823 = io_x[14] ? _GEN11822 : _GEN6843;
wire  _GEN11824 = io_x[0] ? _GEN11823 : _GEN6845;
wire  _GEN11825 = io_x[76] ? _GEN11824 : _GEN6834;
wire  _GEN11826 = io_x[42] ? _GEN6874 : _GEN11825;
wire  _GEN11827 = io_x[38] ? _GEN11826 : _GEN7036;
wire  _GEN11828 = io_x[10] ? _GEN11827 : _GEN11820;
wire  _GEN11829 = io_x[71] ? _GEN11828 : _GEN7196;
wire  _GEN11830 = io_x[70] ? _GEN11829 : _GEN11818;
wire  _GEN11831 = io_x[33] ? _GEN11830 : _GEN11809;
wire  _GEN11832 = io_x[21] ? _GEN11831 : _GEN11681;
wire  _GEN11833 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11834 = io_x[6] ? _GEN6850 : _GEN11833;
wire  _GEN11835 = io_x[41] ? _GEN6836 : _GEN11834;
wire  _GEN11836 = io_x[14] ? _GEN6856 : _GEN11835;
wire  _GEN11837 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11838 = io_x[0] ? _GEN11837 : _GEN11836;
wire  _GEN11839 = io_x[76] ? _GEN6833 : _GEN11838;
wire  _GEN11840 = io_x[42] ? _GEN6874 : _GEN11839;
wire  _GEN11841 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11842 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN11843 = io_x[14] ? _GEN11842 : _GEN11841;
wire  _GEN11844 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN11845 = io_x[14] ? _GEN11844 : _GEN6843;
wire  _GEN11846 = io_x[0] ? _GEN11845 : _GEN11843;
wire  _GEN11847 = io_x[76] ? _GEN11846 : _GEN6833;
wire  _GEN11848 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN11849 = io_x[42] ? _GEN11848 : _GEN11847;
wire  _GEN11850 = io_x[38] ? _GEN11849 : _GEN11840;
wire  _GEN11851 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11852 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11853 = io_x[41] ? _GEN11852 : _GEN11851;
wire  _GEN11854 = io_x[14] ? _GEN11853 : _GEN6856;
wire  _GEN11855 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11856 = io_x[0] ? _GEN11855 : _GEN11854;
wire  _GEN11857 = io_x[76] ? _GEN6834 : _GEN11856;
wire  _GEN11858 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11859 = io_x[0] ? _GEN11858 : _GEN6845;
wire  _GEN11860 = io_x[76] ? _GEN11859 : _GEN6834;
wire  _GEN11861 = io_x[42] ? _GEN11860 : _GEN11857;
wire  _GEN11862 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11863 = io_x[14] ? _GEN11862 : _GEN6843;
wire  _GEN11864 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11865 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11866 = io_x[6] ? _GEN11865 : _GEN6850;
wire  _GEN11867 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11868 = io_x[6] ? _GEN11867 : _GEN6850;
wire  _GEN11869 = io_x[41] ? _GEN11868 : _GEN11866;
wire  _GEN11870 = io_x[14] ? _GEN11869 : _GEN11864;
wire  _GEN11871 = io_x[0] ? _GEN11870 : _GEN11863;
wire  _GEN11872 = io_x[76] ? _GEN11871 : _GEN6833;
wire  _GEN11873 = io_x[42] ? _GEN6874 : _GEN11872;
wire  _GEN11874 = io_x[38] ? _GEN11873 : _GEN11861;
wire  _GEN11875 = io_x[10] ? _GEN11874 : _GEN11850;
wire  _GEN11876 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN11877 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN11878 = io_x[41] ? _GEN6836 : _GEN11877;
wire  _GEN11879 = io_x[14] ? _GEN11878 : _GEN6843;
wire  _GEN11880 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11881 = io_x[6] ? _GEN11880 : _GEN6850;
wire  _GEN11882 = io_x[41] ? _GEN11881 : _GEN6836;
wire  _GEN11883 = io_x[14] ? _GEN11882 : _GEN6843;
wire  _GEN11884 = io_x[0] ? _GEN11883 : _GEN11879;
wire  _GEN11885 = io_x[76] ? _GEN11884 : _GEN6834;
wire  _GEN11886 = io_x[42] ? _GEN11885 : _GEN6863;
wire  _GEN11887 = io_x[38] ? _GEN11886 : _GEN11876;
wire  _GEN11888 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN11889 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN11890 = io_x[42] ? _GEN11889 : _GEN11888;
wire  _GEN11891 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN11892 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11893 = io_x[6] ? _GEN11892 : _GEN6850;
wire  _GEN11894 = io_x[41] ? _GEN11893 : _GEN6836;
wire  _GEN11895 = io_x[14] ? _GEN11894 : _GEN6843;
wire  _GEN11896 = io_x[0] ? _GEN11895 : _GEN6845;
wire  _GEN11897 = io_x[76] ? _GEN11896 : _GEN6834;
wire  _GEN11898 = io_x[42] ? _GEN11897 : _GEN11891;
wire  _GEN11899 = io_x[38] ? _GEN11898 : _GEN11890;
wire  _GEN11900 = io_x[10] ? _GEN11899 : _GEN11887;
wire  _GEN11901 = io_x[71] ? _GEN11900 : _GEN11875;
wire  _GEN11902 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11903 = io_x[2] ? _GEN6837 : _GEN11902;
wire  _GEN11904 = io_x[6] ? _GEN6850 : _GEN11903;
wire  _GEN11905 = io_x[41] ? _GEN6924 : _GEN11904;
wire  _GEN11906 = io_x[14] ? _GEN6843 : _GEN11905;
wire  _GEN11907 = io_x[0] ? _GEN6845 : _GEN11906;
wire  _GEN11908 = io_x[76] ? _GEN11907 : _GEN6833;
wire  _GEN11909 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11910 = io_x[2] ? _GEN6837 : _GEN11909;
wire  _GEN11911 = io_x[6] ? _GEN6850 : _GEN11910;
wire  _GEN11912 = io_x[41] ? _GEN6836 : _GEN11911;
wire  _GEN11913 = io_x[14] ? _GEN6843 : _GEN11912;
wire  _GEN11914 = io_x[0] ? _GEN6858 : _GEN11913;
wire  _GEN11915 = io_x[76] ? _GEN11914 : _GEN6834;
wire  _GEN11916 = io_x[42] ? _GEN11915 : _GEN11908;
wire  _GEN11917 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11918 = io_x[14] ? _GEN11917 : _GEN6843;
wire  _GEN11919 = io_x[0] ? _GEN11918 : _GEN6858;
wire  _GEN11920 = io_x[76] ? _GEN11919 : _GEN6834;
wire  _GEN11921 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11922 = io_x[0] ? _GEN6845 : _GEN11921;
wire  _GEN11923 = io_x[76] ? _GEN11922 : _GEN6834;
wire  _GEN11924 = io_x[42] ? _GEN11923 : _GEN11920;
wire  _GEN11925 = io_x[38] ? _GEN11924 : _GEN11916;
wire  _GEN11926 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN11927 = io_x[14] ? _GEN11926 : _GEN6843;
wire  _GEN11928 = io_x[0] ? _GEN11927 : _GEN6845;
wire  _GEN11929 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11930 = io_x[6] ? _GEN11929 : _GEN6840;
wire  _GEN11931 = io_x[41] ? _GEN6836 : _GEN11930;
wire  _GEN11932 = io_x[14] ? _GEN11931 : _GEN6856;
wire  _GEN11933 = io_x[0] ? _GEN11932 : _GEN6845;
wire  _GEN11934 = io_x[76] ? _GEN11933 : _GEN11928;
wire  _GEN11935 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11936 = io_x[0] ? _GEN11935 : _GEN6845;
wire  _GEN11937 = io_x[76] ? _GEN11936 : _GEN6833;
wire  _GEN11938 = io_x[42] ? _GEN11937 : _GEN11934;
wire  _GEN11939 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11940 = io_x[2] ? _GEN11939 : _GEN6838;
wire  _GEN11941 = io_x[6] ? _GEN11940 : _GEN6850;
wire  _GEN11942 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN11943 = io_x[41] ? _GEN11942 : _GEN11941;
wire  _GEN11944 = io_x[14] ? _GEN11943 : _GEN6843;
wire  _GEN11945 = io_x[0] ? _GEN11944 : _GEN6845;
wire  _GEN11946 = io_x[76] ? _GEN11945 : _GEN6834;
wire  _GEN11947 = io_x[42] ? _GEN6874 : _GEN11946;
wire  _GEN11948 = io_x[38] ? _GEN11947 : _GEN11938;
wire  _GEN11949 = io_x[10] ? _GEN11948 : _GEN11925;
wire  _GEN11950 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN11951 = io_x[0] ? _GEN6845 : _GEN11950;
wire  _GEN11952 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11953 = io_x[2] ? _GEN6837 : _GEN11952;
wire  _GEN11954 = io_x[6] ? _GEN6850 : _GEN11953;
wire  _GEN11955 = io_x[41] ? _GEN6836 : _GEN11954;
wire  _GEN11956 = io_x[14] ? _GEN6843 : _GEN11955;
wire  _GEN11957 = io_x[0] ? _GEN6845 : _GEN11956;
wire  _GEN11958 = io_x[76] ? _GEN11957 : _GEN11951;
wire  _GEN11959 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN11960 = io_x[42] ? _GEN11959 : _GEN11958;
wire  _GEN11961 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN11962 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN11963 = io_x[14] ? _GEN6843 : _GEN11962;
wire  _GEN11964 = io_x[0] ? _GEN11963 : _GEN11961;
wire  _GEN11965 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN11966 = io_x[14] ? _GEN6843 : _GEN11965;
wire  _GEN11967 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN11968 = io_x[6] ? _GEN11967 : _GEN6850;
wire  _GEN11969 = io_x[41] ? _GEN6836 : _GEN11968;
wire  _GEN11970 = io_x[14] ? _GEN11969 : _GEN6843;
wire  _GEN11971 = io_x[0] ? _GEN11970 : _GEN11966;
wire  _GEN11972 = io_x[76] ? _GEN11971 : _GEN11964;
wire  _GEN11973 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11974 = io_x[2] ? _GEN6837 : _GEN11973;
wire  _GEN11975 = io_x[6] ? _GEN6850 : _GEN11974;
wire  _GEN11976 = io_x[41] ? _GEN11975 : _GEN6836;
wire  _GEN11977 = io_x[14] ? _GEN6843 : _GEN11976;
wire  _GEN11978 = io_x[0] ? _GEN6845 : _GEN11977;
wire  _GEN11979 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11980 = io_x[6] ? _GEN6850 : _GEN11979;
wire  _GEN11981 = io_x[41] ? _GEN11980 : _GEN6924;
wire  _GEN11982 = io_x[14] ? _GEN6843 : _GEN11981;
wire  _GEN11983 = io_x[0] ? _GEN6858 : _GEN11982;
wire  _GEN11984 = io_x[76] ? _GEN11983 : _GEN11978;
wire  _GEN11985 = io_x[42] ? _GEN11984 : _GEN11972;
wire  _GEN11986 = io_x[38] ? _GEN11985 : _GEN11960;
wire  _GEN11987 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN11988 = io_x[42] ? _GEN6863 : _GEN11987;
wire  _GEN11989 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN11990 = io_x[6] ? _GEN11989 : _GEN6840;
wire  _GEN11991 = io_x[41] ? _GEN6836 : _GEN11990;
wire  _GEN11992 = io_x[14] ? _GEN11991 : _GEN6843;
wire  _GEN11993 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN11994 = io_x[2] ? _GEN11993 : _GEN6838;
wire  _GEN11995 = io_x[6] ? _GEN11994 : _GEN6840;
wire  _GEN11996 = io_x[41] ? _GEN6836 : _GEN11995;
wire  _GEN11997 = io_x[14] ? _GEN11996 : _GEN6843;
wire  _GEN11998 = io_x[0] ? _GEN11997 : _GEN11992;
wire  _GEN11999 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12000 = io_x[6] ? _GEN11999 : _GEN6850;
wire  _GEN12001 = io_x[41] ? _GEN6836 : _GEN12000;
wire  _GEN12002 = io_x[14] ? _GEN12001 : _GEN6843;
wire  _GEN12003 = io_x[0] ? _GEN12002 : _GEN6845;
wire  _GEN12004 = io_x[76] ? _GEN12003 : _GEN11998;
wire  _GEN12005 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12006 = io_x[6] ? _GEN12005 : _GEN6840;
wire  _GEN12007 = io_x[41] ? _GEN12006 : _GEN6836;
wire  _GEN12008 = io_x[14] ? _GEN12007 : _GEN6843;
wire  _GEN12009 = io_x[0] ? _GEN6845 : _GEN12008;
wire  _GEN12010 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12011 = io_x[41] ? _GEN6836 : _GEN12010;
wire  _GEN12012 = io_x[14] ? _GEN12011 : _GEN6843;
wire  _GEN12013 = io_x[0] ? _GEN6845 : _GEN12012;
wire  _GEN12014 = io_x[76] ? _GEN12013 : _GEN12009;
wire  _GEN12015 = io_x[42] ? _GEN12014 : _GEN12004;
wire  _GEN12016 = io_x[38] ? _GEN12015 : _GEN11988;
wire  _GEN12017 = io_x[10] ? _GEN12016 : _GEN11986;
wire  _GEN12018 = io_x[71] ? _GEN12017 : _GEN11949;
wire  _GEN12019 = io_x[70] ? _GEN12018 : _GEN11901;
wire  _GEN12020 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12021 = io_x[41] ? _GEN6836 : _GEN12020;
wire  _GEN12022 = io_x[14] ? _GEN12021 : _GEN6843;
wire  _GEN12023 = io_x[0] ? _GEN12022 : _GEN6845;
wire  _GEN12024 = io_x[76] ? _GEN12023 : _GEN6834;
wire  _GEN12025 = io_x[42] ? _GEN6874 : _GEN12024;
wire  _GEN12026 = io_x[38] ? _GEN12025 : _GEN6871;
wire  _GEN12027 = io_x[10] ? _GEN12026 : _GEN7044;
wire  _GEN12028 = io_x[71] ? _GEN12027 : _GEN7196;
wire  _GEN12029 = io_x[70] ? _GEN12028 : _GEN7020;
wire  _GEN12030 = io_x[33] ? _GEN12029 : _GEN12019;
wire  _GEN12031 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN12032 = io_x[76] ? _GEN6833 : _GEN12031;
wire  _GEN12033 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN12034 = io_x[42] ? _GEN12033 : _GEN12032;
wire  _GEN12035 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12036 = io_x[41] ? _GEN12035 : _GEN6924;
wire  _GEN12037 = io_x[14] ? _GEN6843 : _GEN12036;
wire  _GEN12038 = io_x[0] ? _GEN6858 : _GEN12037;
wire  _GEN12039 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12040 = io_x[2] ? _GEN6837 : _GEN12039;
wire  _GEN12041 = io_x[6] ? _GEN6850 : _GEN12040;
wire  _GEN12042 = io_x[41] ? _GEN6836 : _GEN12041;
wire  _GEN12043 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12044 = io_x[6] ? _GEN12043 : _GEN6850;
wire  _GEN12045 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12046 = io_x[6] ? _GEN12045 : _GEN6850;
wire  _GEN12047 = io_x[41] ? _GEN12046 : _GEN12044;
wire  _GEN12048 = io_x[14] ? _GEN12047 : _GEN12042;
wire  _GEN12049 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN12050 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12051 = io_x[6] ? _GEN12050 : _GEN6840;
wire  _GEN12052 = io_x[41] ? _GEN12051 : _GEN6836;
wire  _GEN12053 = io_x[14] ? _GEN12052 : _GEN12049;
wire  _GEN12054 = io_x[0] ? _GEN12053 : _GEN12048;
wire  _GEN12055 = io_x[76] ? _GEN12054 : _GEN12038;
wire  _GEN12056 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12057 = io_x[2] ? _GEN6837 : _GEN12056;
wire  _GEN12058 = io_x[6] ? _GEN6850 : _GEN12057;
wire  _GEN12059 = io_x[41] ? _GEN12058 : _GEN6924;
wire  _GEN12060 = io_x[14] ? _GEN6843 : _GEN12059;
wire  _GEN12061 = io_x[0] ? _GEN6845 : _GEN12060;
wire  _GEN12062 = io_x[76] ? _GEN6834 : _GEN12061;
wire  _GEN12063 = io_x[42] ? _GEN12062 : _GEN12055;
wire  _GEN12064 = io_x[38] ? _GEN12063 : _GEN12034;
wire  _GEN12065 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12066 = io_x[41] ? _GEN6924 : _GEN12065;
wire  _GEN12067 = io_x[14] ? _GEN12066 : _GEN6843;
wire  _GEN12068 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12069 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12070 = io_x[41] ? _GEN12069 : _GEN12068;
wire  _GEN12071 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN12072 = io_x[2] ? _GEN12071 : _GEN6837;
wire  _GEN12073 = io_x[6] ? _GEN6840 : _GEN12072;
wire  _GEN12074 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12075 = io_x[41] ? _GEN12074 : _GEN12073;
wire  _GEN12076 = io_x[14] ? _GEN12075 : _GEN12070;
wire  _GEN12077 = io_x[0] ? _GEN12076 : _GEN12067;
wire  _GEN12078 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN12079 = io_x[0] ? _GEN6858 : _GEN12078;
wire  _GEN12080 = io_x[76] ? _GEN12079 : _GEN12077;
wire  _GEN12081 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN12082 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12083 = io_x[6] ? _GEN12082 : _GEN6850;
wire  _GEN12084 = io_x[41] ? _GEN12083 : _GEN6836;
wire  _GEN12085 = io_x[14] ? _GEN12084 : _GEN6856;
wire  _GEN12086 = io_x[0] ? _GEN12085 : _GEN12081;
wire  _GEN12087 = io_x[76] ? _GEN12086 : _GEN6834;
wire  _GEN12088 = io_x[42] ? _GEN12087 : _GEN12080;
wire  _GEN12089 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12090 = io_x[6] ? _GEN12089 : _GEN6850;
wire  _GEN12091 = io_x[41] ? _GEN6836 : _GEN12090;
wire  _GEN12092 = io_x[14] ? _GEN12091 : _GEN6843;
wire  _GEN12093 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN12094 = io_x[0] ? _GEN12093 : _GEN12092;
wire  _GEN12095 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12096 = io_x[41] ? _GEN12095 : _GEN6836;
wire  _GEN12097 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12098 = io_x[2] ? _GEN12097 : _GEN6837;
wire  _GEN12099 = io_x[6] ? _GEN12098 : _GEN6850;
wire  _GEN12100 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12101 = io_x[6] ? _GEN12100 : _GEN6840;
wire  _GEN12102 = io_x[41] ? _GEN12101 : _GEN12099;
wire  _GEN12103 = io_x[14] ? _GEN12102 : _GEN12096;
wire  _GEN12104 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12105 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12106 = io_x[6] ? _GEN12105 : _GEN12104;
wire  _GEN12107 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12108 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12109 = io_x[6] ? _GEN12108 : _GEN12107;
wire  _GEN12110 = io_x[41] ? _GEN12109 : _GEN12106;
wire  _GEN12111 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12112 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12113 = io_x[6] ? _GEN12112 : _GEN12111;
wire  _GEN12114 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12115 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12116 = io_x[6] ? _GEN12115 : _GEN12114;
wire  _GEN12117 = io_x[41] ? _GEN12116 : _GEN12113;
wire  _GEN12118 = io_x[14] ? _GEN12117 : _GEN12110;
wire  _GEN12119 = io_x[0] ? _GEN12118 : _GEN12103;
wire  _GEN12120 = io_x[76] ? _GEN12119 : _GEN12094;
wire  _GEN12121 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12122 = io_x[6] ? _GEN12121 : _GEN6850;
wire  _GEN12123 = io_x[41] ? _GEN12122 : _GEN6836;
wire  _GEN12124 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12125 = io_x[2] ? _GEN12124 : _GEN6837;
wire  _GEN12126 = io_x[6] ? _GEN12125 : _GEN6840;
wire  _GEN12127 = io_x[41] ? _GEN6924 : _GEN12126;
wire  _GEN12128 = io_x[14] ? _GEN12127 : _GEN12123;
wire  _GEN12129 = io_x[0] ? _GEN12128 : _GEN6858;
wire  _GEN12130 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12131 = io_x[2] ? _GEN12130 : _GEN6837;
wire  _GEN12132 = io_x[6] ? _GEN12131 : _GEN6850;
wire  _GEN12133 = io_x[41] ? _GEN12132 : _GEN6836;
wire  _GEN12134 = io_x[14] ? _GEN12133 : _GEN6843;
wire  _GEN12135 = io_x[0] ? _GEN6858 : _GEN12134;
wire  _GEN12136 = io_x[76] ? _GEN12135 : _GEN12129;
wire  _GEN12137 = io_x[42] ? _GEN12136 : _GEN12120;
wire  _GEN12138 = io_x[38] ? _GEN12137 : _GEN12088;
wire  _GEN12139 = io_x[10] ? _GEN12138 : _GEN12064;
wire  _GEN12140 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12141 = io_x[41] ? _GEN6836 : _GEN12140;
wire  _GEN12142 = io_x[14] ? _GEN12141 : _GEN6856;
wire  _GEN12143 = io_x[0] ? _GEN12142 : _GEN6858;
wire  _GEN12144 = io_x[76] ? _GEN12143 : _GEN6833;
wire  _GEN12145 = io_x[42] ? _GEN6874 : _GEN12144;
wire  _GEN12146 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12147 = io_x[2] ? _GEN6837 : _GEN12146;
wire  _GEN12148 = io_x[6] ? _GEN6850 : _GEN12147;
wire  _GEN12149 = io_x[41] ? _GEN6924 : _GEN12148;
wire  _GEN12150 = io_x[14] ? _GEN6843 : _GEN12149;
wire  _GEN12151 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12152 = io_x[41] ? _GEN12151 : _GEN6836;
wire  _GEN12153 = io_x[14] ? _GEN6843 : _GEN12152;
wire  _GEN12154 = io_x[0] ? _GEN12153 : _GEN12150;
wire  _GEN12155 = io_x[76] ? _GEN12154 : _GEN6833;
wire  _GEN12156 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN12157 = io_x[14] ? _GEN6843 : _GEN12156;
wire  _GEN12158 = io_x[0] ? _GEN6858 : _GEN12157;
wire  _GEN12159 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12160 = io_x[6] ? _GEN12159 : _GEN6850;
wire  _GEN12161 = io_x[41] ? _GEN12160 : _GEN6836;
wire  _GEN12162 = io_x[14] ? _GEN12161 : _GEN6843;
wire  _GEN12163 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12164 = io_x[6] ? _GEN12163 : _GEN6850;
wire  _GEN12165 = io_x[41] ? _GEN12164 : _GEN6836;
wire  _GEN12166 = io_x[14] ? _GEN12165 : _GEN6843;
wire  _GEN12167 = io_x[0] ? _GEN12166 : _GEN12162;
wire  _GEN12168 = io_x[76] ? _GEN12167 : _GEN12158;
wire  _GEN12169 = io_x[42] ? _GEN12168 : _GEN12155;
wire  _GEN12170 = io_x[38] ? _GEN12169 : _GEN12145;
wire  _GEN12171 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12172 = io_x[2] ? _GEN12171 : _GEN6837;
wire  _GEN12173 = io_x[6] ? _GEN12172 : _GEN6840;
wire  _GEN12174 = io_x[41] ? _GEN6924 : _GEN12173;
wire  _GEN12175 = io_x[14] ? _GEN12174 : _GEN6843;
wire  _GEN12176 = io_x[0] ? _GEN12175 : _GEN6845;
wire  _GEN12177 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12178 = io_x[41] ? _GEN12177 : _GEN6836;
wire  _GEN12179 = io_x[14] ? _GEN12178 : _GEN6843;
wire  _GEN12180 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN12181 = io_x[0] ? _GEN12180 : _GEN12179;
wire  _GEN12182 = io_x[76] ? _GEN12181 : _GEN12176;
wire  _GEN12183 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12184 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12185 = io_x[41] ? _GEN12184 : _GEN12183;
wire  _GEN12186 = io_x[14] ? _GEN12185 : _GEN6843;
wire  _GEN12187 = io_x[0] ? _GEN12186 : _GEN6845;
wire  _GEN12188 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12189 = io_x[41] ? _GEN12188 : _GEN6836;
wire  _GEN12190 = io_x[14] ? _GEN12189 : _GEN6856;
wire  _GEN12191 = io_x[0] ? _GEN12190 : _GEN6845;
wire  _GEN12192 = io_x[76] ? _GEN12191 : _GEN12187;
wire  _GEN12193 = io_x[42] ? _GEN12192 : _GEN12182;
wire  _GEN12194 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12195 = io_x[41] ? _GEN6836 : _GEN12194;
wire  _GEN12196 = io_x[14] ? _GEN12195 : _GEN6843;
wire  _GEN12197 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN12198 = io_x[0] ? _GEN12197 : _GEN12196;
wire  _GEN12199 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN12200 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN12201 = io_x[2] ? _GEN12200 : _GEN6837;
wire  _GEN12202 = io_x[6] ? _GEN12201 : _GEN6840;
wire  _GEN12203 = io_x[41] ? _GEN12202 : _GEN6836;
wire  _GEN12204 = io_x[14] ? _GEN6856 : _GEN12203;
wire  _GEN12205 = io_x[0] ? _GEN12204 : _GEN12199;
wire  _GEN12206 = io_x[76] ? _GEN12205 : _GEN12198;
wire  _GEN12207 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12208 = io_x[41] ? _GEN6836 : _GEN12207;
wire  _GEN12209 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12210 = io_x[2] ? _GEN12209 : _GEN6838;
wire  _GEN12211 = io_x[6] ? _GEN12210 : _GEN6850;
wire  _GEN12212 = io_x[41] ? _GEN12211 : _GEN6836;
wire  _GEN12213 = io_x[14] ? _GEN12212 : _GEN12208;
wire  _GEN12214 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12215 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12216 = io_x[6] ? _GEN12215 : _GEN6850;
wire  _GEN12217 = io_x[41] ? _GEN12216 : _GEN12214;
wire  _GEN12218 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12219 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12220 = io_x[6] ? _GEN12219 : _GEN12218;
wire  _GEN12221 = io_x[41] ? _GEN12220 : _GEN6836;
wire  _GEN12222 = io_x[14] ? _GEN12221 : _GEN12217;
wire  _GEN12223 = io_x[0] ? _GEN12222 : _GEN12213;
wire  _GEN12224 = io_x[76] ? _GEN12223 : _GEN6833;
wire  _GEN12225 = io_x[42] ? _GEN12224 : _GEN12206;
wire  _GEN12226 = io_x[38] ? _GEN12225 : _GEN12193;
wire  _GEN12227 = io_x[10] ? _GEN12226 : _GEN12170;
wire  _GEN12228 = io_x[71] ? _GEN12227 : _GEN12139;
wire  _GEN12229 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12230 = io_x[41] ? _GEN6836 : _GEN12229;
wire  _GEN12231 = io_x[14] ? _GEN12230 : _GEN6856;
wire  _GEN12232 = io_x[0] ? _GEN12231 : _GEN6858;
wire  _GEN12233 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12234 = io_x[2] ? _GEN6837 : _GEN12233;
wire  _GEN12235 = io_x[6] ? _GEN6850 : _GEN12234;
wire  _GEN12236 = io_x[41] ? _GEN6924 : _GEN12235;
wire  _GEN12237 = io_x[14] ? _GEN6843 : _GEN12236;
wire  _GEN12238 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12239 = io_x[41] ? _GEN12238 : _GEN6836;
wire  _GEN12240 = io_x[14] ? _GEN12239 : _GEN6843;
wire  _GEN12241 = io_x[0] ? _GEN12240 : _GEN12237;
wire  _GEN12242 = io_x[76] ? _GEN12241 : _GEN12232;
wire  _GEN12243 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN12244 = io_x[0] ? _GEN12243 : _GEN6858;
wire  _GEN12245 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN12246 = io_x[0] ? _GEN12245 : _GEN6858;
wire  _GEN12247 = io_x[76] ? _GEN12246 : _GEN12244;
wire  _GEN12248 = io_x[42] ? _GEN12247 : _GEN12242;
wire  _GEN12249 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12250 = io_x[2] ? _GEN6837 : _GEN12249;
wire  _GEN12251 = io_x[6] ? _GEN6850 : _GEN12250;
wire  _GEN12252 = io_x[41] ? _GEN6924 : _GEN12251;
wire  _GEN12253 = io_x[14] ? _GEN6843 : _GEN12252;
wire  _GEN12254 = io_x[0] ? _GEN6845 : _GEN12253;
wire  _GEN12255 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12256 = io_x[41] ? _GEN12255 : _GEN6924;
wire  _GEN12257 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN12258 = io_x[2] ? _GEN12257 : _GEN6837;
wire  _GEN12259 = io_x[6] ? _GEN12258 : _GEN6850;
wire  _GEN12260 = io_x[41] ? _GEN6924 : _GEN12259;
wire  _GEN12261 = io_x[14] ? _GEN12260 : _GEN12256;
wire  _GEN12262 = io_x[0] ? _GEN12261 : _GEN6858;
wire  _GEN12263 = io_x[76] ? _GEN12262 : _GEN12254;
wire  _GEN12264 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN12265 = io_x[42] ? _GEN12264 : _GEN12263;
wire  _GEN12266 = io_x[38] ? _GEN12265 : _GEN12248;
wire  _GEN12267 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12268 = io_x[41] ? _GEN6924 : _GEN12267;
wire  _GEN12269 = io_x[14] ? _GEN12268 : _GEN6843;
wire  _GEN12270 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12271 = io_x[6] ? _GEN12270 : _GEN6850;
wire  _GEN12272 = io_x[41] ? _GEN6836 : _GEN12271;
wire  _GEN12273 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12274 = io_x[6] ? _GEN12273 : _GEN6850;
wire  _GEN12275 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12276 = io_x[6] ? _GEN12275 : _GEN6850;
wire  _GEN12277 = io_x[41] ? _GEN12276 : _GEN12274;
wire  _GEN12278 = io_x[14] ? _GEN12277 : _GEN12272;
wire  _GEN12279 = io_x[0] ? _GEN12278 : _GEN12269;
wire  _GEN12280 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12281 = io_x[6] ? _GEN12280 : _GEN6840;
wire  _GEN12282 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12283 = io_x[2] ? _GEN12282 : _GEN6837;
wire  _GEN12284 = io_x[6] ? _GEN12283 : _GEN6850;
wire  _GEN12285 = io_x[41] ? _GEN12284 : _GEN12281;
wire  _GEN12286 = io_x[14] ? _GEN12285 : _GEN6856;
wire  _GEN12287 = io_x[0] ? _GEN12286 : _GEN6845;
wire  _GEN12288 = io_x[76] ? _GEN12287 : _GEN12279;
wire  _GEN12289 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12290 = io_x[41] ? _GEN12289 : _GEN6836;
wire  _GEN12291 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12292 = io_x[2] ? _GEN12291 : _GEN6837;
wire  _GEN12293 = io_x[6] ? _GEN12292 : _GEN6850;
wire  _GEN12294 = io_x[41] ? _GEN12293 : _GEN6924;
wire  _GEN12295 = io_x[14] ? _GEN12294 : _GEN12290;
wire  _GEN12296 = io_x[0] ? _GEN12295 : _GEN6858;
wire  _GEN12297 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12298 = io_x[2] ? _GEN12297 : _GEN6837;
wire  _GEN12299 = io_x[6] ? _GEN12298 : _GEN6840;
wire  _GEN12300 = io_x[41] ? _GEN12299 : _GEN6836;
wire  _GEN12301 = io_x[14] ? _GEN12300 : _GEN6856;
wire  _GEN12302 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN12303 = io_x[2] ? _GEN12302 : _GEN6837;
wire  _GEN12304 = io_x[6] ? _GEN12303 : _GEN6850;
wire  _GEN12305 = io_x[41] ? _GEN12304 : _GEN6924;
wire  _GEN12306 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12307 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12308 = io_x[2] ? _GEN12307 : _GEN6837;
wire  _GEN12309 = io_x[6] ? _GEN12308 : _GEN6850;
wire  _GEN12310 = io_x[41] ? _GEN12309 : _GEN12306;
wire  _GEN12311 = io_x[14] ? _GEN12310 : _GEN12305;
wire  _GEN12312 = io_x[0] ? _GEN12311 : _GEN12301;
wire  _GEN12313 = io_x[76] ? _GEN12312 : _GEN12296;
wire  _GEN12314 = io_x[42] ? _GEN12313 : _GEN12288;
wire  _GEN12315 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12316 = io_x[41] ? _GEN6924 : _GEN12315;
wire  _GEN12317 = io_x[14] ? _GEN12316 : _GEN6856;
wire  _GEN12318 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN12319 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12320 = io_x[2] ? _GEN12319 : _GEN6838;
wire  _GEN12321 = io_x[6] ? _GEN12320 : _GEN6840;
wire  _GEN12322 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12323 = io_x[6] ? _GEN12322 : _GEN6840;
wire  _GEN12324 = io_x[41] ? _GEN12323 : _GEN12321;
wire  _GEN12325 = io_x[14] ? _GEN12324 : _GEN12318;
wire  _GEN12326 = io_x[0] ? _GEN12325 : _GEN12317;
wire  _GEN12327 = io_x[76] ? _GEN12326 : _GEN6833;
wire  _GEN12328 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN12329 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12330 = io_x[41] ? _GEN12329 : _GEN6924;
wire  _GEN12331 = io_x[14] ? _GEN12330 : _GEN12328;
wire  _GEN12332 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN12333 = io_x[2] ? _GEN12332 : _GEN6837;
wire  _GEN12334 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12335 = io_x[2] ? _GEN12334 : _GEN6837;
wire  _GEN12336 = io_x[6] ? _GEN12335 : _GEN12333;
wire  _GEN12337 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12338 = io_x[6] ? _GEN12337 : _GEN6840;
wire  _GEN12339 = io_x[41] ? _GEN12338 : _GEN12336;
wire  _GEN12340 = io_x[14] ? _GEN12339 : _GEN6843;
wire  _GEN12341 = io_x[0] ? _GEN12340 : _GEN12331;
wire  _GEN12342 = io_x[76] ? _GEN12341 : _GEN6833;
wire  _GEN12343 = io_x[42] ? _GEN12342 : _GEN12327;
wire  _GEN12344 = io_x[38] ? _GEN12343 : _GEN12314;
wire  _GEN12345 = io_x[10] ? _GEN12344 : _GEN12266;
wire  _GEN12346 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12347 = io_x[41] ? _GEN6924 : _GEN12346;
wire  _GEN12348 = io_x[14] ? _GEN12347 : _GEN6856;
wire  _GEN12349 = io_x[0] ? _GEN12348 : _GEN6845;
wire  _GEN12350 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12351 = io_x[2] ? _GEN6837 : _GEN12350;
wire  _GEN12352 = io_x[6] ? _GEN6850 : _GEN12351;
wire  _GEN12353 = io_x[41] ? _GEN6836 : _GEN12352;
wire  _GEN12354 = io_x[14] ? _GEN6843 : _GEN12353;
wire  _GEN12355 = io_x[0] ? _GEN6858 : _GEN12354;
wire  _GEN12356 = io_x[76] ? _GEN12355 : _GEN12349;
wire  _GEN12357 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12358 = io_x[2] ? _GEN6837 : _GEN12357;
wire  _GEN12359 = io_x[6] ? _GEN6850 : _GEN12358;
wire  _GEN12360 = io_x[41] ? _GEN6836 : _GEN12359;
wire  _GEN12361 = io_x[14] ? _GEN6843 : _GEN12360;
wire  _GEN12362 = io_x[0] ? _GEN6845 : _GEN12361;
wire  _GEN12363 = io_x[76] ? _GEN12362 : _GEN6834;
wire  _GEN12364 = io_x[42] ? _GEN12363 : _GEN12356;
wire  _GEN12365 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12366 = io_x[41] ? _GEN6836 : _GEN12365;
wire  _GEN12367 = io_x[14] ? _GEN12366 : _GEN6843;
wire  _GEN12368 = io_x[0] ? _GEN6858 : _GEN12367;
wire  _GEN12369 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12370 = io_x[6] ? _GEN12369 : _GEN6850;
wire  _GEN12371 = io_x[41] ? _GEN6836 : _GEN12370;
wire  _GEN12372 = io_x[14] ? _GEN12371 : _GEN6856;
wire  _GEN12373 = io_x[0] ? _GEN6845 : _GEN12372;
wire  _GEN12374 = io_x[76] ? _GEN12373 : _GEN12368;
wire  _GEN12375 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12376 = io_x[41] ? _GEN12375 : _GEN6836;
wire  _GEN12377 = io_x[14] ? _GEN12376 : _GEN6843;
wire  _GEN12378 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN12379 = io_x[0] ? _GEN12378 : _GEN12377;
wire  _GEN12380 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN12381 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12382 = io_x[41] ? _GEN6836 : _GEN12381;
wire  _GEN12383 = io_x[14] ? _GEN12382 : _GEN12380;
wire  _GEN12384 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12385 = io_x[6] ? _GEN12384 : _GEN6850;
wire  _GEN12386 = io_x[41] ? _GEN12385 : _GEN6836;
wire  _GEN12387 = io_x[14] ? _GEN12386 : _GEN6843;
wire  _GEN12388 = io_x[0] ? _GEN12387 : _GEN12383;
wire  _GEN12389 = io_x[76] ? _GEN12388 : _GEN12379;
wire  _GEN12390 = io_x[42] ? _GEN12389 : _GEN12374;
wire  _GEN12391 = io_x[38] ? _GEN12390 : _GEN12364;
wire  _GEN12392 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN12393 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12394 = io_x[41] ? _GEN6924 : _GEN12393;
wire  _GEN12395 = io_x[14] ? _GEN12394 : _GEN12392;
wire  _GEN12396 = io_x[0] ? _GEN12395 : _GEN6858;
wire  _GEN12397 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12398 = io_x[6] ? _GEN12397 : _GEN6850;
wire  _GEN12399 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12400 = io_x[2] ? _GEN12399 : _GEN6837;
wire  _GEN12401 = io_x[6] ? _GEN12400 : _GEN6850;
wire  _GEN12402 = io_x[41] ? _GEN12401 : _GEN12398;
wire  _GEN12403 = io_x[14] ? _GEN12402 : _GEN6843;
wire  _GEN12404 = io_x[0] ? _GEN12403 : _GEN6845;
wire  _GEN12405 = io_x[76] ? _GEN12404 : _GEN12396;
wire  _GEN12406 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12407 = io_x[6] ? _GEN12406 : _GEN6850;
wire  _GEN12408 = io_x[41] ? _GEN12407 : _GEN6836;
wire  _GEN12409 = io_x[14] ? _GEN12408 : _GEN6843;
wire  _GEN12410 = io_x[0] ? _GEN12409 : _GEN6858;
wire  _GEN12411 = io_x[76] ? _GEN6833 : _GEN12410;
wire  _GEN12412 = io_x[42] ? _GEN12411 : _GEN12405;
wire  _GEN12413 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12414 = io_x[41] ? _GEN6924 : _GEN12413;
wire  _GEN12415 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12416 = io_x[2] ? _GEN12415 : _GEN6837;
wire  _GEN12417 = io_x[6] ? _GEN12416 : _GEN6850;
wire  _GEN12418 = io_x[41] ? _GEN6924 : _GEN12417;
wire  _GEN12419 = io_x[14] ? _GEN12418 : _GEN12414;
wire  _GEN12420 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12421 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12422 = io_x[41] ? _GEN12421 : _GEN12420;
wire  _GEN12423 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN12424 = io_x[2] ? _GEN12423 : _GEN6837;
wire  _GEN12425 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12426 = io_x[2] ? _GEN12425 : _GEN6837;
wire  _GEN12427 = io_x[6] ? _GEN12426 : _GEN12424;
wire  _GEN12428 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12429 = io_x[2] ? _GEN12428 : _GEN6837;
wire  _GEN12430 = io_x[6] ? _GEN12429 : _GEN6840;
wire  _GEN12431 = io_x[41] ? _GEN12430 : _GEN12427;
wire  _GEN12432 = io_x[14] ? _GEN12431 : _GEN12422;
wire  _GEN12433 = io_x[0] ? _GEN12432 : _GEN12419;
wire  _GEN12434 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12435 = io_x[6] ? _GEN12434 : _GEN6850;
wire  _GEN12436 = io_x[41] ? _GEN6836 : _GEN12435;
wire  _GEN12437 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12438 = io_x[6] ? _GEN12437 : _GEN6850;
wire  _GEN12439 = io_x[41] ? _GEN6836 : _GEN12438;
wire  _GEN12440 = io_x[14] ? _GEN12439 : _GEN12436;
wire  _GEN12441 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12442 = io_x[6] ? _GEN12441 : _GEN6840;
wire  _GEN12443 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12444 = io_x[41] ? _GEN12443 : _GEN12442;
wire  _GEN12445 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12446 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12447 = io_x[6] ? _GEN12446 : _GEN12445;
wire  _GEN12448 = io_x[41] ? _GEN6924 : _GEN12447;
wire  _GEN12449 = io_x[14] ? _GEN12448 : _GEN12444;
wire  _GEN12450 = io_x[0] ? _GEN12449 : _GEN12440;
wire  _GEN12451 = io_x[76] ? _GEN12450 : _GEN12433;
wire  _GEN12452 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12453 = io_x[41] ? _GEN12452 : _GEN6836;
wire  _GEN12454 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12455 = io_x[41] ? _GEN12454 : _GEN6836;
wire  _GEN12456 = io_x[14] ? _GEN12455 : _GEN12453;
wire  _GEN12457 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12458 = io_x[6] ? _GEN12457 : _GEN6850;
wire  _GEN12459 = io_x[41] ? _GEN6924 : _GEN12458;
wire  _GEN12460 = io_x[14] ? _GEN12459 : _GEN6843;
wire  _GEN12461 = io_x[0] ? _GEN12460 : _GEN12456;
wire  _GEN12462 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12463 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12464 = io_x[6] ? _GEN12463 : _GEN6850;
wire  _GEN12465 = io_x[41] ? _GEN12464 : _GEN12462;
wire  _GEN12466 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12467 = io_x[6] ? _GEN12466 : _GEN6850;
wire  _GEN12468 = io_x[41] ? _GEN12467 : _GEN6924;
wire  _GEN12469 = io_x[14] ? _GEN12468 : _GEN12465;
wire  _GEN12470 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12471 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12472 = io_x[6] ? _GEN12471 : _GEN6850;
wire  _GEN12473 = io_x[41] ? _GEN12472 : _GEN12470;
wire  _GEN12474 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12475 = io_x[6] ? _GEN12474 : _GEN6840;
wire  _GEN12476 = io_x[41] ? _GEN12475 : _GEN6836;
wire  _GEN12477 = io_x[14] ? _GEN12476 : _GEN12473;
wire  _GEN12478 = io_x[0] ? _GEN12477 : _GEN12469;
wire  _GEN12479 = io_x[76] ? _GEN12478 : _GEN12461;
wire  _GEN12480 = io_x[42] ? _GEN12479 : _GEN12451;
wire  _GEN12481 = io_x[38] ? _GEN12480 : _GEN12412;
wire  _GEN12482 = io_x[10] ? _GEN12481 : _GEN12391;
wire  _GEN12483 = io_x[71] ? _GEN12482 : _GEN12345;
wire  _GEN12484 = io_x[70] ? _GEN12483 : _GEN12228;
wire  _GEN12485 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12486 = io_x[41] ? _GEN6924 : _GEN12485;
wire  _GEN12487 = io_x[14] ? _GEN12486 : _GEN6843;
wire  _GEN12488 = io_x[0] ? _GEN12487 : _GEN6845;
wire  _GEN12489 = io_x[76] ? _GEN6834 : _GEN12488;
wire  _GEN12490 = io_x[42] ? _GEN6874 : _GEN12489;
wire  _GEN12491 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12492 = io_x[41] ? _GEN6836 : _GEN12491;
wire  _GEN12493 = io_x[14] ? _GEN12492 : _GEN6843;
wire  _GEN12494 = io_x[0] ? _GEN12493 : _GEN6858;
wire  _GEN12495 = io_x[76] ? _GEN12494 : _GEN6833;
wire  _GEN12496 = io_x[42] ? _GEN6874 : _GEN12495;
wire  _GEN12497 = io_x[38] ? _GEN12496 : _GEN12490;
wire  _GEN12498 = io_x[10] ? _GEN12497 : _GEN7094;
wire  _GEN12499 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12500 = io_x[41] ? _GEN6836 : _GEN12499;
wire  _GEN12501 = io_x[14] ? _GEN12500 : _GEN6843;
wire  _GEN12502 = io_x[0] ? _GEN12501 : _GEN6845;
wire  _GEN12503 = io_x[76] ? _GEN12502 : _GEN6834;
wire  _GEN12504 = io_x[42] ? _GEN6874 : _GEN12503;
wire  _GEN12505 = io_x[38] ? _GEN7036 : _GEN12504;
wire  _GEN12506 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12507 = io_x[41] ? _GEN6836 : _GEN12506;
wire  _GEN12508 = io_x[14] ? _GEN12507 : _GEN6843;
wire  _GEN12509 = io_x[0] ? _GEN12508 : _GEN6845;
wire  _GEN12510 = io_x[76] ? _GEN12509 : _GEN6834;
wire  _GEN12511 = io_x[42] ? _GEN6874 : _GEN12510;
wire  _GEN12512 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12513 = io_x[6] ? _GEN12512 : _GEN6850;
wire  _GEN12514 = io_x[41] ? _GEN12513 : _GEN6924;
wire  _GEN12515 = io_x[14] ? _GEN12514 : _GEN6843;
wire  _GEN12516 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12517 = io_x[6] ? _GEN12516 : _GEN6840;
wire  _GEN12518 = io_x[41] ? _GEN12517 : _GEN6836;
wire  _GEN12519 = io_x[14] ? _GEN12518 : _GEN6856;
wire  _GEN12520 = io_x[0] ? _GEN12519 : _GEN12515;
wire  _GEN12521 = io_x[76] ? _GEN12520 : _GEN6834;
wire  _GEN12522 = io_x[42] ? _GEN12521 : _GEN6874;
wire  _GEN12523 = io_x[38] ? _GEN12522 : _GEN12511;
wire  _GEN12524 = io_x[10] ? _GEN12523 : _GEN12505;
wire  _GEN12525 = io_x[71] ? _GEN12524 : _GEN12498;
wire  _GEN12526 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12527 = io_x[41] ? _GEN6836 : _GEN12526;
wire  _GEN12528 = io_x[14] ? _GEN12527 : _GEN6843;
wire  _GEN12529 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12530 = io_x[6] ? _GEN12529 : _GEN6850;
wire  _GEN12531 = io_x[41] ? _GEN6836 : _GEN12530;
wire  _GEN12532 = io_x[14] ? _GEN12531 : _GEN6843;
wire  _GEN12533 = io_x[0] ? _GEN12532 : _GEN12528;
wire  _GEN12534 = io_x[76] ? _GEN12533 : _GEN6834;
wire  _GEN12535 = io_x[42] ? _GEN6874 : _GEN12534;
wire  _GEN12536 = io_x[38] ? _GEN12535 : _GEN6871;
wire  _GEN12537 = io_x[10] ? _GEN12536 : _GEN7044;
wire  _GEN12538 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12539 = io_x[6] ? _GEN12538 : _GEN6850;
wire  _GEN12540 = io_x[41] ? _GEN6836 : _GEN12539;
wire  _GEN12541 = io_x[14] ? _GEN12540 : _GEN6856;
wire  _GEN12542 = io_x[0] ? _GEN12541 : _GEN6845;
wire  _GEN12543 = io_x[76] ? _GEN12542 : _GEN6834;
wire  _GEN12544 = io_x[42] ? _GEN6863 : _GEN12543;
wire  _GEN12545 = io_x[38] ? _GEN12544 : _GEN6871;
wire  _GEN12546 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12547 = io_x[41] ? _GEN6836 : _GEN12546;
wire  _GEN12548 = io_x[14] ? _GEN12547 : _GEN6843;
wire  _GEN12549 = io_x[0] ? _GEN6845 : _GEN12548;
wire  _GEN12550 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12551 = io_x[6] ? _GEN12550 : _GEN6840;
wire  _GEN12552 = io_x[41] ? _GEN6836 : _GEN12551;
wire  _GEN12553 = io_x[14] ? _GEN12552 : _GEN6856;
wire  _GEN12554 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12555 = io_x[6] ? _GEN12554 : _GEN6840;
wire  _GEN12556 = io_x[41] ? _GEN6836 : _GEN12555;
wire  _GEN12557 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12558 = io_x[6] ? _GEN12557 : _GEN6850;
wire  _GEN12559 = io_x[41] ? _GEN6836 : _GEN12558;
wire  _GEN12560 = io_x[14] ? _GEN12559 : _GEN12556;
wire  _GEN12561 = io_x[0] ? _GEN12560 : _GEN12553;
wire  _GEN12562 = io_x[76] ? _GEN12561 : _GEN12549;
wire  _GEN12563 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12564 = io_x[41] ? _GEN12563 : _GEN6836;
wire  _GEN12565 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN12566 = io_x[6] ? _GEN12565 : _GEN6850;
wire  _GEN12567 = io_x[41] ? _GEN12566 : _GEN6836;
wire  _GEN12568 = io_x[14] ? _GEN12567 : _GEN12564;
wire  _GEN12569 = io_x[0] ? _GEN12568 : _GEN6845;
wire  _GEN12570 = io_x[76] ? _GEN12569 : _GEN6834;
wire  _GEN12571 = io_x[42] ? _GEN12570 : _GEN12562;
wire  _GEN12572 = io_x[38] ? _GEN12571 : _GEN6871;
wire  _GEN12573 = io_x[10] ? _GEN12572 : _GEN12545;
wire  _GEN12574 = io_x[71] ? _GEN12573 : _GEN12537;
wire  _GEN12575 = io_x[70] ? _GEN12574 : _GEN12525;
wire  _GEN12576 = io_x[33] ? _GEN12575 : _GEN12484;
wire  _GEN12577 = io_x[21] ? _GEN12576 : _GEN12030;
wire  _GEN12578 = io_x[18] ? _GEN12577 : _GEN11832;
wire  _GEN12579 = io_x[20] ? _GEN12578 : _GEN11594;
wire  _GEN12580 = io_x[45] ? _GEN12579 : _GEN11204;
wire  _GEN12581 = io_x[28] ? _GEN12580 : _GEN9291;
wire  _GEN12582 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN12583 = io_x[14] ? _GEN6843 : _GEN12582;
wire  _GEN12584 = io_x[0] ? _GEN6845 : _GEN12583;
wire  _GEN12585 = io_x[76] ? _GEN6834 : _GEN12584;
wire  _GEN12586 = io_x[42] ? _GEN6874 : _GEN12585;
wire  _GEN12587 = io_x[38] ? _GEN12586 : _GEN6871;
wire  _GEN12588 = io_x[10] ? _GEN7044 : _GEN12587;
wire  _GEN12589 = io_x[71] ? _GEN7203 : _GEN12588;
wire  _GEN12590 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN12591 = io_x[14] ? _GEN6856 : _GEN12590;
wire  _GEN12592 = io_x[0] ? _GEN6845 : _GEN12591;
wire  _GEN12593 = io_x[76] ? _GEN6834 : _GEN12592;
wire  _GEN12594 = io_x[42] ? _GEN6874 : _GEN12593;
wire  _GEN12595 = io_x[38] ? _GEN12594 : _GEN6871;
wire  _GEN12596 = io_x[10] ? _GEN7094 : _GEN12595;
wire  _GEN12597 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN12598 = io_x[76] ? _GEN6834 : _GEN12597;
wire  _GEN12599 = io_x[42] ? _GEN6874 : _GEN12598;
wire  _GEN12600 = io_x[38] ? _GEN6871 : _GEN12599;
wire  _GEN12601 = io_x[10] ? _GEN7044 : _GEN12600;
wire  _GEN12602 = io_x[71] ? _GEN12601 : _GEN12596;
wire  _GEN12603 = io_x[70] ? _GEN12602 : _GEN12589;
wire  _GEN12604 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN12605 = io_x[76] ? _GEN6834 : _GEN12604;
wire  _GEN12606 = io_x[42] ? _GEN6874 : _GEN12605;
wire  _GEN12607 = io_x[38] ? _GEN12606 : _GEN6871;
wire  _GEN12608 = io_x[10] ? _GEN7044 : _GEN12607;
wire  _GEN12609 = io_x[71] ? _GEN12608 : _GEN7196;
wire  _GEN12610 = io_x[70] ? _GEN8474 : _GEN12609;
wire  _GEN12611 = io_x[33] ? _GEN12610 : _GEN12603;
wire  _GEN12612 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN12613 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN12614 = io_x[10] ? _GEN7044 : _GEN12613;
wire  _GEN12615 = io_x[71] ? _GEN12614 : _GEN12612;
wire  _GEN12616 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12617 = io_x[6] ? _GEN6850 : _GEN12616;
wire  _GEN12618 = io_x[41] ? _GEN6836 : _GEN12617;
wire  _GEN12619 = io_x[14] ? _GEN6856 : _GEN12618;
wire  _GEN12620 = io_x[0] ? _GEN6845 : _GEN12619;
wire  _GEN12621 = io_x[76] ? _GEN6834 : _GEN12620;
wire  _GEN12622 = io_x[42] ? _GEN6874 : _GEN12621;
wire  _GEN12623 = io_x[38] ? _GEN12622 : _GEN6871;
wire  _GEN12624 = io_x[10] ? _GEN7044 : _GEN12623;
wire  _GEN12625 = io_x[71] ? _GEN7196 : _GEN12624;
wire  _GEN12626 = io_x[70] ? _GEN12625 : _GEN12615;
wire  _GEN12627 = 1'b1;
wire  _GEN12628 = io_x[33] ? _GEN12627 : _GEN12626;
wire  _GEN12629 = io_x[21] ? _GEN12628 : _GEN12611;
wire  _GEN12630 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN12631 = io_x[14] ? _GEN6856 : _GEN12630;
wire  _GEN12632 = io_x[0] ? _GEN6845 : _GEN12631;
wire  _GEN12633 = io_x[76] ? _GEN6834 : _GEN12632;
wire  _GEN12634 = io_x[42] ? _GEN6874 : _GEN12633;
wire  _GEN12635 = io_x[38] ? _GEN12634 : _GEN6871;
wire  _GEN12636 = io_x[10] ? _GEN7044 : _GEN12635;
wire  _GEN12637 = io_x[71] ? _GEN7196 : _GEN12636;
wire  _GEN12638 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN12639 = io_x[71] ? _GEN12638 : _GEN7203;
wire  _GEN12640 = io_x[70] ? _GEN12639 : _GEN12637;
wire  _GEN12641 = 1'b0;
wire  _GEN12642 = io_x[33] ? _GEN12641 : _GEN12640;
wire  _GEN12643 = 1'b1;
wire  _GEN12644 = io_x[21] ? _GEN12643 : _GEN12642;
wire  _GEN12645 = io_x[18] ? _GEN12644 : _GEN12629;
wire  _GEN12646 = io_x[33] ? _GEN12627 : _GEN12641;
wire  _GEN12647 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN12648 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN12649 = io_x[42] ? _GEN6874 : _GEN12648;
wire  _GEN12650 = io_x[38] ? _GEN12649 : _GEN6871;
wire  _GEN12651 = io_x[10] ? _GEN7044 : _GEN12650;
wire  _GEN12652 = io_x[71] ? _GEN12651 : _GEN12647;
wire  _GEN12653 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN12654 = io_x[71] ? _GEN7196 : _GEN12653;
wire  _GEN12655 = io_x[70] ? _GEN12654 : _GEN12652;
wire  _GEN12656 = io_x[33] ? _GEN12627 : _GEN12655;
wire  _GEN12657 = io_x[21] ? _GEN12656 : _GEN12646;
wire  _GEN12658 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN12659 = io_x[0] ? _GEN6845 : _GEN12658;
wire  _GEN12660 = io_x[76] ? _GEN6834 : _GEN12659;
wire  _GEN12661 = io_x[42] ? _GEN6874 : _GEN12660;
wire  _GEN12662 = io_x[38] ? _GEN12661 : _GEN6871;
wire  _GEN12663 = io_x[10] ? _GEN7044 : _GEN12662;
wire  _GEN12664 = io_x[71] ? _GEN7196 : _GEN12663;
wire  _GEN12665 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN12666 = io_x[14] ? _GEN6843 : _GEN12665;
wire  _GEN12667 = io_x[0] ? _GEN6845 : _GEN12666;
wire  _GEN12668 = io_x[76] ? _GEN6834 : _GEN12667;
wire  _GEN12669 = io_x[42] ? _GEN6874 : _GEN12668;
wire  _GEN12670 = io_x[38] ? _GEN12669 : _GEN6871;
wire  _GEN12671 = io_x[10] ? _GEN7044 : _GEN12670;
wire  _GEN12672 = io_x[71] ? _GEN7196 : _GEN12671;
wire  _GEN12673 = io_x[70] ? _GEN12672 : _GEN12664;
wire  _GEN12674 = io_x[33] ? _GEN12627 : _GEN12673;
wire  _GEN12675 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12676 = io_x[6] ? _GEN6850 : _GEN12675;
wire  _GEN12677 = io_x[41] ? _GEN6924 : _GEN12676;
wire  _GEN12678 = io_x[14] ? _GEN6843 : _GEN12677;
wire  _GEN12679 = io_x[0] ? _GEN6845 : _GEN12678;
wire  _GEN12680 = io_x[76] ? _GEN6834 : _GEN12679;
wire  _GEN12681 = io_x[42] ? _GEN6863 : _GEN12680;
wire  _GEN12682 = io_x[38] ? _GEN12681 : _GEN6871;
wire  _GEN12683 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN12684 = io_x[10] ? _GEN12683 : _GEN12682;
wire  _GEN12685 = io_x[71] ? _GEN7196 : _GEN12684;
wire  _GEN12686 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN12687 = io_x[14] ? _GEN6843 : _GEN12686;
wire  _GEN12688 = io_x[0] ? _GEN6845 : _GEN12687;
wire  _GEN12689 = io_x[76] ? _GEN6834 : _GEN12688;
wire  _GEN12690 = io_x[42] ? _GEN6874 : _GEN12689;
wire  _GEN12691 = io_x[38] ? _GEN12690 : _GEN6871;
wire  _GEN12692 = io_x[10] ? _GEN7094 : _GEN12691;
wire  _GEN12693 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN12694 = io_x[38] ? _GEN6871 : _GEN12693;
wire  _GEN12695 = io_x[10] ? _GEN7044 : _GEN12694;
wire  _GEN12696 = io_x[71] ? _GEN12695 : _GEN12692;
wire  _GEN12697 = io_x[70] ? _GEN12696 : _GEN12685;
wire  _GEN12698 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN12699 = io_x[10] ? _GEN7044 : _GEN12698;
wire  _GEN12700 = io_x[71] ? _GEN12699 : _GEN7203;
wire  _GEN12701 = io_x[70] ? _GEN8474 : _GEN12700;
wire  _GEN12702 = io_x[33] ? _GEN12701 : _GEN12697;
wire  _GEN12703 = io_x[21] ? _GEN12702 : _GEN12674;
wire  _GEN12704 = io_x[18] ? _GEN12703 : _GEN12657;
wire  _GEN12705 = io_x[20] ? _GEN12704 : _GEN12645;
wire  _GEN12706 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN12707 = io_x[42] ? _GEN6863 : _GEN12706;
wire  _GEN12708 = io_x[38] ? _GEN12707 : _GEN7036;
wire  _GEN12709 = io_x[10] ? _GEN7044 : _GEN12708;
wire  _GEN12710 = io_x[71] ? _GEN12709 : _GEN7196;
wire  _GEN12711 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN12712 = io_x[10] ? _GEN7044 : _GEN12711;
wire  _GEN12713 = io_x[71] ? _GEN12712 : _GEN7196;
wire  _GEN12714 = io_x[70] ? _GEN12713 : _GEN12710;
wire  _GEN12715 = io_x[33] ? _GEN12641 : _GEN12714;
wire  _GEN12716 = io_x[71] ? _GEN7203 : _GEN7196;
wire  _GEN12717 = io_x[70] ? _GEN7020 : _GEN12716;
wire  _GEN12718 = io_x[33] ? _GEN12627 : _GEN12717;
wire  _GEN12719 = io_x[21] ? _GEN12718 : _GEN12715;
wire  _GEN12720 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN12721 = io_x[42] ? _GEN6863 : _GEN12720;
wire  _GEN12722 = io_x[38] ? _GEN12721 : _GEN6871;
wire  _GEN12723 = io_x[10] ? _GEN7044 : _GEN12722;
wire  _GEN12724 = io_x[71] ? _GEN12723 : _GEN7196;
wire  _GEN12725 = io_x[70] ? _GEN8474 : _GEN12724;
wire  _GEN12726 = io_x[33] ? _GEN12627 : _GEN12725;
wire  _GEN12727 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN12728 = io_x[71] ? _GEN12727 : _GEN7196;
wire  _GEN12729 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN12730 = io_x[38] ? _GEN6871 : _GEN12729;
wire  _GEN12731 = io_x[10] ? _GEN7044 : _GEN12730;
wire  _GEN12732 = io_x[71] ? _GEN12731 : _GEN7196;
wire  _GEN12733 = io_x[70] ? _GEN12732 : _GEN12728;
wire  _GEN12734 = io_x[33] ? _GEN12627 : _GEN12733;
wire  _GEN12735 = io_x[21] ? _GEN12734 : _GEN12726;
wire  _GEN12736 = io_x[18] ? _GEN12735 : _GEN12719;
wire  _GEN12737 = io_x[70] ? _GEN8474 : _GEN7020;
wire  _GEN12738 = io_x[33] ? _GEN12627 : _GEN12737;
wire  _GEN12739 = io_x[71] ? _GEN7203 : _GEN7196;
wire  _GEN12740 = io_x[70] ? _GEN8474 : _GEN12739;
wire  _GEN12741 = io_x[33] ? _GEN12627 : _GEN12740;
wire  _GEN12742 = io_x[21] ? _GEN12741 : _GEN12738;
wire  _GEN12743 = io_x[70] ? _GEN8474 : _GEN7020;
wire  _GEN12744 = io_x[33] ? _GEN12627 : _GEN12743;
wire  _GEN12745 = io_x[21] ? _GEN12744 : _GEN12643;
wire  _GEN12746 = io_x[18] ? _GEN12745 : _GEN12742;
wire  _GEN12747 = io_x[20] ? _GEN12746 : _GEN12736;
wire  _GEN12748 = io_x[45] ? _GEN12747 : _GEN12705;
wire  _GEN12749 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN12750 = io_x[71] ? _GEN7196 : _GEN12749;
wire  _GEN12751 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN12752 = io_x[10] ? _GEN12751 : _GEN7044;
wire  _GEN12753 = io_x[71] ? _GEN7203 : _GEN12752;
wire  _GEN12754 = io_x[70] ? _GEN12753 : _GEN12750;
wire  _GEN12755 = io_x[33] ? _GEN12627 : _GEN12754;
wire  _GEN12756 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN12757 = io_x[71] ? _GEN12756 : _GEN7203;
wire  _GEN12758 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN12759 = io_x[10] ? _GEN12758 : _GEN7094;
wire  _GEN12760 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN12761 = io_x[38] ? _GEN6871 : _GEN12760;
wire  _GEN12762 = io_x[10] ? _GEN7044 : _GEN12761;
wire  _GEN12763 = io_x[71] ? _GEN12762 : _GEN12759;
wire  _GEN12764 = io_x[70] ? _GEN12763 : _GEN12757;
wire  _GEN12765 = io_x[33] ? _GEN12627 : _GEN12764;
wire  _GEN12766 = io_x[21] ? _GEN12765 : _GEN12755;
wire  _GEN12767 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN12768 = io_x[14] ? _GEN6856 : _GEN12767;
wire  _GEN12769 = io_x[0] ? _GEN6845 : _GEN12768;
wire  _GEN12770 = io_x[76] ? _GEN6834 : _GEN12769;
wire  _GEN12771 = io_x[42] ? _GEN6874 : _GEN12770;
wire  _GEN12772 = io_x[38] ? _GEN12771 : _GEN6871;
wire  _GEN12773 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN12774 = io_x[0] ? _GEN6845 : _GEN12773;
wire  _GEN12775 = io_x[76] ? _GEN6834 : _GEN12774;
wire  _GEN12776 = io_x[42] ? _GEN6874 : _GEN12775;
wire  _GEN12777 = io_x[38] ? _GEN12776 : _GEN6871;
wire  _GEN12778 = io_x[10] ? _GEN12777 : _GEN12772;
wire  _GEN12779 = io_x[71] ? _GEN7203 : _GEN12778;
wire  _GEN12780 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN12781 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN12782 = io_x[71] ? _GEN12781 : _GEN12780;
wire  _GEN12783 = io_x[70] ? _GEN12782 : _GEN12779;
wire  _GEN12784 = io_x[33] ? _GEN12641 : _GEN12783;
wire  _GEN12785 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN12786 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN12787 = io_x[38] ? _GEN6871 : _GEN12786;
wire  _GEN12788 = io_x[10] ? _GEN12787 : _GEN12785;
wire  _GEN12789 = io_x[71] ? _GEN7203 : _GEN12788;
wire  _GEN12790 = io_x[70] ? _GEN7020 : _GEN12789;
wire  _GEN12791 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN12792 = io_x[71] ? _GEN12791 : _GEN7203;
wire  _GEN12793 = io_x[70] ? _GEN7020 : _GEN12792;
wire  _GEN12794 = io_x[33] ? _GEN12793 : _GEN12790;
wire  _GEN12795 = io_x[21] ? _GEN12794 : _GEN12784;
wire  _GEN12796 = io_x[18] ? _GEN12795 : _GEN12766;
wire  _GEN12797 = io_x[33] ? _GEN12627 : _GEN12641;
wire  _GEN12798 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12799 = io_x[2] ? _GEN6837 : _GEN12798;
wire  _GEN12800 = io_x[6] ? _GEN6850 : _GEN12799;
wire  _GEN12801 = io_x[41] ? _GEN12800 : _GEN6836;
wire  _GEN12802 = io_x[14] ? _GEN6843 : _GEN12801;
wire  _GEN12803 = io_x[0] ? _GEN6845 : _GEN12802;
wire  _GEN12804 = io_x[76] ? _GEN6834 : _GEN12803;
wire  _GEN12805 = io_x[42] ? _GEN6874 : _GEN12804;
wire  _GEN12806 = io_x[38] ? _GEN7036 : _GEN12805;
wire  _GEN12807 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN12808 = io_x[10] ? _GEN12807 : _GEN12806;
wire  _GEN12809 = io_x[71] ? _GEN7203 : _GEN12808;
wire  _GEN12810 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12811 = io_x[41] ? _GEN12810 : _GEN6836;
wire  _GEN12812 = io_x[14] ? _GEN12811 : _GEN6843;
wire  _GEN12813 = io_x[0] ? _GEN6845 : _GEN12812;
wire  _GEN12814 = io_x[76] ? _GEN12813 : _GEN6834;
wire  _GEN12815 = io_x[42] ? _GEN6874 : _GEN12814;
wire  _GEN12816 = io_x[38] ? _GEN12815 : _GEN6871;
wire  _GEN12817 = io_x[10] ? _GEN12816 : _GEN7044;
wire  _GEN12818 = io_x[71] ? _GEN7196 : _GEN12817;
wire  _GEN12819 = io_x[70] ? _GEN12818 : _GEN12809;
wire  _GEN12820 = io_x[33] ? _GEN12641 : _GEN12819;
wire  _GEN12821 = io_x[21] ? _GEN12820 : _GEN12797;
wire  _GEN12822 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12823 = io_x[2] ? _GEN6837 : _GEN12822;
wire  _GEN12824 = io_x[6] ? _GEN6850 : _GEN12823;
wire  _GEN12825 = io_x[41] ? _GEN12824 : _GEN6836;
wire  _GEN12826 = io_x[14] ? _GEN6843 : _GEN12825;
wire  _GEN12827 = io_x[0] ? _GEN6845 : _GEN12826;
wire  _GEN12828 = io_x[76] ? _GEN6834 : _GEN12827;
wire  _GEN12829 = io_x[42] ? _GEN6874 : _GEN12828;
wire  _GEN12830 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN12831 = io_x[14] ? _GEN6843 : _GEN12830;
wire  _GEN12832 = io_x[0] ? _GEN6845 : _GEN12831;
wire  _GEN12833 = io_x[76] ? _GEN6834 : _GEN12832;
wire  _GEN12834 = io_x[42] ? _GEN6863 : _GEN12833;
wire  _GEN12835 = io_x[38] ? _GEN12834 : _GEN12829;
wire  _GEN12836 = io_x[10] ? _GEN7094 : _GEN12835;
wire  _GEN12837 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN12838 = io_x[38] ? _GEN12837 : _GEN6871;
wire  _GEN12839 = io_x[10] ? _GEN7094 : _GEN12838;
wire  _GEN12840 = io_x[71] ? _GEN12839 : _GEN12836;
wire  _GEN12841 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN12842 = io_x[14] ? _GEN6843 : _GEN12841;
wire  _GEN12843 = io_x[0] ? _GEN6845 : _GEN12842;
wire  _GEN12844 = io_x[76] ? _GEN6834 : _GEN12843;
wire  _GEN12845 = io_x[42] ? _GEN6874 : _GEN12844;
wire  _GEN12846 = io_x[38] ? _GEN12845 : _GEN6871;
wire  _GEN12847 = io_x[10] ? _GEN7094 : _GEN12846;
wire  _GEN12848 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN12849 = io_x[10] ? _GEN12848 : _GEN7044;
wire  _GEN12850 = io_x[71] ? _GEN12849 : _GEN12847;
wire  _GEN12851 = io_x[70] ? _GEN12850 : _GEN12840;
wire  _GEN12852 = io_x[33] ? _GEN12627 : _GEN12851;
wire  _GEN12853 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN12854 = io_x[2] ? _GEN6837 : _GEN12853;
wire  _GEN12855 = io_x[6] ? _GEN6850 : _GEN12854;
wire  _GEN12856 = io_x[41] ? _GEN12855 : _GEN6836;
wire  _GEN12857 = io_x[14] ? _GEN6843 : _GEN12856;
wire  _GEN12858 = io_x[0] ? _GEN6845 : _GEN12857;
wire  _GEN12859 = io_x[76] ? _GEN6834 : _GEN12858;
wire  _GEN12860 = io_x[42] ? _GEN6874 : _GEN12859;
wire  _GEN12861 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN12862 = io_x[14] ? _GEN6843 : _GEN12861;
wire  _GEN12863 = io_x[0] ? _GEN6845 : _GEN12862;
wire  _GEN12864 = io_x[76] ? _GEN6834 : _GEN12863;
wire  _GEN12865 = io_x[42] ? _GEN6874 : _GEN12864;
wire  _GEN12866 = io_x[38] ? _GEN12865 : _GEN12860;
wire  _GEN12867 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12868 = io_x[41] ? _GEN6836 : _GEN12867;
wire  _GEN12869 = io_x[14] ? _GEN12868 : _GEN6843;
wire  _GEN12870 = io_x[0] ? _GEN12869 : _GEN6845;
wire  _GEN12871 = io_x[76] ? _GEN6834 : _GEN12870;
wire  _GEN12872 = io_x[42] ? _GEN12871 : _GEN6874;
wire  _GEN12873 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN12874 = io_x[0] ? _GEN12873 : _GEN6845;
wire  _GEN12875 = io_x[76] ? _GEN6834 : _GEN12874;
wire  _GEN12876 = io_x[42] ? _GEN12875 : _GEN6874;
wire  _GEN12877 = io_x[38] ? _GEN12876 : _GEN12872;
wire  _GEN12878 = io_x[10] ? _GEN12877 : _GEN12866;
wire  _GEN12879 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN12880 = io_x[0] ? _GEN12879 : _GEN6845;
wire  _GEN12881 = io_x[76] ? _GEN6834 : _GEN12880;
wire  _GEN12882 = io_x[42] ? _GEN6874 : _GEN12881;
wire  _GEN12883 = io_x[38] ? _GEN12882 : _GEN7036;
wire  _GEN12884 = io_x[10] ? _GEN12883 : _GEN7094;
wire  _GEN12885 = io_x[71] ? _GEN12884 : _GEN12878;
wire  _GEN12886 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN12887 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN12888 = io_x[76] ? _GEN12887 : _GEN12886;
wire  _GEN12889 = io_x[42] ? _GEN6874 : _GEN12888;
wire  _GEN12890 = io_x[38] ? _GEN12889 : _GEN6871;
wire  _GEN12891 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12892 = io_x[41] ? _GEN12891 : _GEN6836;
wire  _GEN12893 = io_x[14] ? _GEN12892 : _GEN6843;
wire  _GEN12894 = io_x[0] ? _GEN6858 : _GEN12893;
wire  _GEN12895 = io_x[76] ? _GEN12894 : _GEN6834;
wire  _GEN12896 = io_x[42] ? _GEN6874 : _GEN12895;
wire  _GEN12897 = io_x[38] ? _GEN12896 : _GEN6871;
wire  _GEN12898 = io_x[10] ? _GEN12897 : _GEN12890;
wire  _GEN12899 = io_x[71] ? _GEN7196 : _GEN12898;
wire  _GEN12900 = io_x[70] ? _GEN12899 : _GEN12885;
wire  _GEN12901 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN12902 = io_x[41] ? _GEN12901 : _GEN6836;
wire  _GEN12903 = io_x[14] ? _GEN12902 : _GEN6843;
wire  _GEN12904 = io_x[0] ? _GEN12903 : _GEN6845;
wire  _GEN12905 = io_x[76] ? _GEN6834 : _GEN12904;
wire  _GEN12906 = io_x[42] ? _GEN6874 : _GEN12905;
wire  _GEN12907 = io_x[38] ? _GEN12906 : _GEN6871;
wire  _GEN12908 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN12909 = io_x[0] ? _GEN12908 : _GEN6845;
wire  _GEN12910 = io_x[76] ? _GEN6834 : _GEN12909;
wire  _GEN12911 = io_x[42] ? _GEN6874 : _GEN12910;
wire  _GEN12912 = io_x[38] ? _GEN12911 : _GEN6871;
wire  _GEN12913 = io_x[10] ? _GEN12912 : _GEN12907;
wire  _GEN12914 = io_x[71] ? _GEN12913 : _GEN7203;
wire  _GEN12915 = io_x[70] ? _GEN8474 : _GEN12914;
wire  _GEN12916 = io_x[33] ? _GEN12915 : _GEN12900;
wire  _GEN12917 = io_x[21] ? _GEN12916 : _GEN12852;
wire  _GEN12918 = io_x[18] ? _GEN12917 : _GEN12821;
wire  _GEN12919 = io_x[20] ? _GEN12918 : _GEN12796;
wire  _GEN12920 = 1'b0;
wire  _GEN12921 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN12922 = io_x[71] ? _GEN12921 : _GEN7196;
wire  _GEN12923 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN12924 = io_x[42] ? _GEN12923 : _GEN6874;
wire  _GEN12925 = io_x[38] ? _GEN6871 : _GEN12924;
wire  _GEN12926 = io_x[10] ? _GEN7044 : _GEN12925;
wire  _GEN12927 = io_x[71] ? _GEN12926 : _GEN7203;
wire  _GEN12928 = io_x[70] ? _GEN12927 : _GEN12922;
wire  _GEN12929 = io_x[33] ? _GEN12627 : _GEN12928;
wire  _GEN12930 = io_x[33] ? _GEN12627 : _GEN12641;
wire  _GEN12931 = io_x[21] ? _GEN12930 : _GEN12929;
wire  _GEN12932 = io_x[18] ? _GEN12931 : _GEN12920;
wire  _GEN12933 = 1'b0;
wire  _GEN12934 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN12935 = io_x[10] ? _GEN12934 : _GEN7094;
wire  _GEN12936 = io_x[71] ? _GEN7203 : _GEN12935;
wire  _GEN12937 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN12938 = io_x[0] ? _GEN6845 : _GEN12937;
wire  _GEN12939 = io_x[76] ? _GEN12938 : _GEN6834;
wire  _GEN12940 = io_x[42] ? _GEN6874 : _GEN12939;
wire  _GEN12941 = io_x[38] ? _GEN12940 : _GEN6871;
wire  _GEN12942 = io_x[10] ? _GEN12941 : _GEN7094;
wire  _GEN12943 = io_x[71] ? _GEN12942 : _GEN7203;
wire  _GEN12944 = io_x[70] ? _GEN12943 : _GEN12936;
wire  _GEN12945 = io_x[33] ? _GEN12627 : _GEN12944;
wire  _GEN12946 = io_x[21] ? _GEN12945 : _GEN12933;
wire  _GEN12947 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN12948 = io_x[38] ? _GEN7036 : _GEN12947;
wire  _GEN12949 = io_x[10] ? _GEN7044 : _GEN12948;
wire  _GEN12950 = io_x[71] ? _GEN7196 : _GEN12949;
wire  _GEN12951 = io_x[70] ? _GEN12950 : _GEN7020;
wire  _GEN12952 = io_x[33] ? _GEN12627 : _GEN12951;
wire  _GEN12953 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN12954 = io_x[41] ? _GEN12953 : _GEN6836;
wire  _GEN12955 = io_x[14] ? _GEN12954 : _GEN6843;
wire  _GEN12956 = io_x[0] ? _GEN12955 : _GEN6858;
wire  _GEN12957 = io_x[76] ? _GEN6834 : _GEN12956;
wire  _GEN12958 = io_x[42] ? _GEN6874 : _GEN12957;
wire  _GEN12959 = io_x[38] ? _GEN12958 : _GEN6871;
wire  _GEN12960 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN12961 = io_x[0] ? _GEN12960 : _GEN6845;
wire  _GEN12962 = io_x[76] ? _GEN6834 : _GEN12961;
wire  _GEN12963 = io_x[42] ? _GEN6874 : _GEN12962;
wire  _GEN12964 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN12965 = io_x[42] ? _GEN6874 : _GEN12964;
wire  _GEN12966 = io_x[38] ? _GEN12965 : _GEN12963;
wire  _GEN12967 = io_x[10] ? _GEN12966 : _GEN12959;
wire  _GEN12968 = io_x[71] ? _GEN12967 : _GEN7196;
wire  _GEN12969 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN12970 = io_x[42] ? _GEN6874 : _GEN12969;
wire  _GEN12971 = io_x[38] ? _GEN7036 : _GEN12970;
wire  _GEN12972 = io_x[10] ? _GEN7044 : _GEN12971;
wire  _GEN12973 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN12974 = io_x[71] ? _GEN12973 : _GEN12972;
wire  _GEN12975 = io_x[70] ? _GEN12974 : _GEN12968;
wire  _GEN12976 = io_x[33] ? _GEN12641 : _GEN12975;
wire  _GEN12977 = io_x[21] ? _GEN12976 : _GEN12952;
wire  _GEN12978 = io_x[18] ? _GEN12977 : _GEN12946;
wire  _GEN12979 = io_x[20] ? _GEN12978 : _GEN12932;
wire  _GEN12980 = io_x[45] ? _GEN12979 : _GEN12919;
wire  _GEN12981 = io_x[28] ? _GEN12980 : _GEN12748;
wire  _GEN12982 = io_x[79] ? _GEN12981 : _GEN12581;
wire  _GEN12983 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN12984 = io_x[0] ? _GEN6845 : _GEN12983;
wire  _GEN12985 = io_x[76] ? _GEN6833 : _GEN12984;
wire  _GEN12986 = io_x[42] ? _GEN12985 : _GEN6874;
wire  _GEN12987 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN12988 = io_x[42] ? _GEN12987 : _GEN6874;
wire  _GEN12989 = io_x[38] ? _GEN12988 : _GEN12986;
wire  _GEN12990 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN12991 = io_x[0] ? _GEN12990 : _GEN6845;
wire  _GEN12992 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN12993 = io_x[0] ? _GEN12992 : _GEN6845;
wire  _GEN12994 = io_x[76] ? _GEN12993 : _GEN12991;
wire  _GEN12995 = io_x[42] ? _GEN12994 : _GEN6874;
wire  _GEN12996 = io_x[38] ? _GEN7036 : _GEN12995;
wire  _GEN12997 = io_x[10] ? _GEN12996 : _GEN12989;
wire  _GEN12998 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN12999 = io_x[6] ? _GEN12998 : _GEN6850;
wire  _GEN13000 = io_x[41] ? _GEN6836 : _GEN12999;
wire  _GEN13001 = io_x[14] ? _GEN6843 : _GEN13000;
wire  _GEN13002 = io_x[0] ? _GEN13001 : _GEN6845;
wire  _GEN13003 = io_x[76] ? _GEN6834 : _GEN13002;
wire  _GEN13004 = io_x[42] ? _GEN13003 : _GEN6874;
wire  _GEN13005 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13006 = io_x[0] ? _GEN6845 : _GEN13005;
wire  _GEN13007 = io_x[76] ? _GEN13006 : _GEN6833;
wire  _GEN13008 = io_x[42] ? _GEN13007 : _GEN6874;
wire  _GEN13009 = io_x[38] ? _GEN13008 : _GEN13004;
wire  _GEN13010 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13011 = io_x[0] ? _GEN6845 : _GEN13010;
wire  _GEN13012 = io_x[76] ? _GEN6834 : _GEN13011;
wire  _GEN13013 = io_x[42] ? _GEN13012 : _GEN6874;
wire  _GEN13014 = io_x[38] ? _GEN13013 : _GEN6871;
wire  _GEN13015 = io_x[10] ? _GEN13014 : _GEN13009;
wire  _GEN13016 = io_x[71] ? _GEN13015 : _GEN12997;
wire  _GEN13017 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13018 = io_x[0] ? _GEN6845 : _GEN13017;
wire  _GEN13019 = io_x[76] ? _GEN13018 : _GEN6834;
wire  _GEN13020 = io_x[42] ? _GEN13019 : _GEN6863;
wire  _GEN13021 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13022 = io_x[6] ? _GEN6850 : _GEN13021;
wire  _GEN13023 = io_x[41] ? _GEN6836 : _GEN13022;
wire  _GEN13024 = io_x[14] ? _GEN13023 : _GEN6843;
wire  _GEN13025 = io_x[0] ? _GEN13024 : _GEN6845;
wire  _GEN13026 = io_x[76] ? _GEN13025 : _GEN6834;
wire  _GEN13027 = io_x[42] ? _GEN13026 : _GEN6874;
wire  _GEN13028 = io_x[38] ? _GEN13027 : _GEN13020;
wire  _GEN13029 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13030 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13031 = io_x[0] ? _GEN13030 : _GEN13029;
wire  _GEN13032 = io_x[76] ? _GEN13031 : _GEN6834;
wire  _GEN13033 = io_x[42] ? _GEN13032 : _GEN6874;
wire  _GEN13034 = io_x[38] ? _GEN7036 : _GEN13033;
wire  _GEN13035 = io_x[10] ? _GEN13034 : _GEN13028;
wire  _GEN13036 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13037 = io_x[6] ? _GEN6850 : _GEN13036;
wire  _GEN13038 = io_x[41] ? _GEN13037 : _GEN6836;
wire  _GEN13039 = io_x[14] ? _GEN6843 : _GEN13038;
wire  _GEN13040 = io_x[0] ? _GEN13039 : _GEN6845;
wire  _GEN13041 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13042 = io_x[6] ? _GEN6850 : _GEN13041;
wire  _GEN13043 = io_x[41] ? _GEN6836 : _GEN13042;
wire  _GEN13044 = io_x[14] ? _GEN13043 : _GEN6843;
wire  _GEN13045 = io_x[0] ? _GEN13044 : _GEN6858;
wire  _GEN13046 = io_x[76] ? _GEN13045 : _GEN13040;
wire  _GEN13047 = io_x[42] ? _GEN13046 : _GEN6863;
wire  _GEN13048 = io_x[38] ? _GEN13047 : _GEN6871;
wire  _GEN13049 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13050 = io_x[0] ? _GEN13049 : _GEN6845;
wire  _GEN13051 = io_x[76] ? _GEN13050 : _GEN6834;
wire  _GEN13052 = io_x[42] ? _GEN13051 : _GEN6874;
wire  _GEN13053 = io_x[38] ? _GEN13052 : _GEN6871;
wire  _GEN13054 = io_x[10] ? _GEN13053 : _GEN13048;
wire  _GEN13055 = io_x[71] ? _GEN13054 : _GEN13035;
wire  _GEN13056 = io_x[70] ? _GEN13055 : _GEN13016;
wire  _GEN13057 = io_x[33] ? _GEN12641 : _GEN13056;
wire  _GEN13058 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13059 = io_x[0] ? _GEN6858 : _GEN13058;
wire  _GEN13060 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13061 = io_x[41] ? _GEN13060 : _GEN6836;
wire  _GEN13062 = io_x[14] ? _GEN6843 : _GEN13061;
wire  _GEN13063 = io_x[0] ? _GEN6845 : _GEN13062;
wire  _GEN13064 = io_x[76] ? _GEN13063 : _GEN13059;
wire  _GEN13065 = io_x[42] ? _GEN13064 : _GEN6874;
wire  _GEN13066 = io_x[38] ? _GEN6871 : _GEN13065;
wire  _GEN13067 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13068 = io_x[0] ? _GEN6845 : _GEN13067;
wire  _GEN13069 = io_x[76] ? _GEN6834 : _GEN13068;
wire  _GEN13070 = io_x[42] ? _GEN13069 : _GEN6874;
wire  _GEN13071 = io_x[38] ? _GEN6871 : _GEN13070;
wire  _GEN13072 = io_x[10] ? _GEN13071 : _GEN13066;
wire  _GEN13073 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13074 = io_x[41] ? _GEN6836 : _GEN13073;
wire  _GEN13075 = io_x[14] ? _GEN13074 : _GEN6843;
wire  _GEN13076 = io_x[0] ? _GEN6858 : _GEN13075;
wire  _GEN13077 = io_x[76] ? _GEN6834 : _GEN13076;
wire  _GEN13078 = io_x[42] ? _GEN13077 : _GEN6874;
wire  _GEN13079 = io_x[38] ? _GEN7036 : _GEN13078;
wire  _GEN13080 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13081 = io_x[0] ? _GEN13080 : _GEN6845;
wire  _GEN13082 = io_x[76] ? _GEN6834 : _GEN13081;
wire  _GEN13083 = io_x[42] ? _GEN13082 : _GEN6874;
wire  _GEN13084 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13085 = io_x[0] ? _GEN6845 : _GEN13084;
wire  _GEN13086 = io_x[76] ? _GEN6834 : _GEN13085;
wire  _GEN13087 = io_x[42] ? _GEN13086 : _GEN6874;
wire  _GEN13088 = io_x[38] ? _GEN13087 : _GEN13083;
wire  _GEN13089 = io_x[10] ? _GEN13088 : _GEN13079;
wire  _GEN13090 = io_x[71] ? _GEN13089 : _GEN13072;
wire  _GEN13091 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN13092 = io_x[6] ? _GEN13091 : _GEN6840;
wire  _GEN13093 = io_x[41] ? _GEN6836 : _GEN13092;
wire  _GEN13094 = io_x[14] ? _GEN6856 : _GEN13093;
wire  _GEN13095 = io_x[0] ? _GEN13094 : _GEN6858;
wire  _GEN13096 = io_x[76] ? _GEN6834 : _GEN13095;
wire  _GEN13097 = io_x[42] ? _GEN13096 : _GEN6874;
wire  _GEN13098 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN13099 = io_x[38] ? _GEN13098 : _GEN13097;
wire  _GEN13100 = io_x[10] ? _GEN7094 : _GEN13099;
wire  _GEN13101 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13102 = io_x[41] ? _GEN6836 : _GEN13101;
wire  _GEN13103 = io_x[14] ? _GEN6856 : _GEN13102;
wire  _GEN13104 = io_x[0] ? _GEN6845 : _GEN13103;
wire  _GEN13105 = io_x[76] ? _GEN6834 : _GEN13104;
wire  _GEN13106 = io_x[42] ? _GEN13105 : _GEN6874;
wire  _GEN13107 = io_x[38] ? _GEN7036 : _GEN13106;
wire  _GEN13108 = io_x[10] ? _GEN7044 : _GEN13107;
wire  _GEN13109 = io_x[71] ? _GEN13108 : _GEN13100;
wire  _GEN13110 = io_x[70] ? _GEN13109 : _GEN13090;
wire  _GEN13111 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13112 = io_x[41] ? _GEN13111 : _GEN6836;
wire  _GEN13113 = io_x[14] ? _GEN6843 : _GEN13112;
wire  _GEN13114 = io_x[0] ? _GEN6845 : _GEN13113;
wire  _GEN13115 = io_x[76] ? _GEN13114 : _GEN6834;
wire  _GEN13116 = io_x[42] ? _GEN13115 : _GEN6874;
wire  _GEN13117 = io_x[38] ? _GEN6871 : _GEN13116;
wire  _GEN13118 = io_x[10] ? _GEN7044 : _GEN13117;
wire  _GEN13119 = io_x[71] ? _GEN7196 : _GEN13118;
wire  _GEN13120 = io_x[70] ? _GEN8474 : _GEN13119;
wire  _GEN13121 = io_x[33] ? _GEN13120 : _GEN13110;
wire  _GEN13122 = io_x[21] ? _GEN13121 : _GEN13057;
wire  _GEN13123 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13124 = io_x[6] ? _GEN6850 : _GEN13123;
wire  _GEN13125 = io_x[41] ? _GEN6836 : _GEN13124;
wire  _GEN13126 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13127 = io_x[41] ? _GEN6836 : _GEN13126;
wire  _GEN13128 = io_x[14] ? _GEN13127 : _GEN13125;
wire  _GEN13129 = io_x[0] ? _GEN13128 : _GEN6858;
wire  _GEN13130 = io_x[76] ? _GEN6834 : _GEN13129;
wire  _GEN13131 = io_x[42] ? _GEN13130 : _GEN6874;
wire  _GEN13132 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13133 = io_x[0] ? _GEN13132 : _GEN6845;
wire  _GEN13134 = io_x[76] ? _GEN13133 : _GEN6834;
wire  _GEN13135 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13136 = io_x[0] ? _GEN13135 : _GEN6845;
wire  _GEN13137 = io_x[76] ? _GEN13136 : _GEN6833;
wire  _GEN13138 = io_x[42] ? _GEN13137 : _GEN13134;
wire  _GEN13139 = io_x[38] ? _GEN13138 : _GEN13131;
wire  _GEN13140 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13141 = io_x[6] ? _GEN13140 : _GEN6850;
wire  _GEN13142 = io_x[41] ? _GEN13141 : _GEN6836;
wire  _GEN13143 = io_x[14] ? _GEN13142 : _GEN6843;
wire  _GEN13144 = io_x[0] ? _GEN13143 : _GEN6845;
wire  _GEN13145 = io_x[76] ? _GEN13144 : _GEN6834;
wire  _GEN13146 = io_x[42] ? _GEN6874 : _GEN13145;
wire  _GEN13147 = io_x[38] ? _GEN13146 : _GEN6871;
wire  _GEN13148 = io_x[10] ? _GEN13147 : _GEN13139;
wire  _GEN13149 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN13150 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13151 = io_x[41] ? _GEN6836 : _GEN13150;
wire  _GEN13152 = io_x[14] ? _GEN6843 : _GEN13151;
wire  _GEN13153 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13154 = io_x[0] ? _GEN13153 : _GEN13152;
wire  _GEN13155 = io_x[76] ? _GEN6834 : _GEN13154;
wire  _GEN13156 = io_x[42] ? _GEN13155 : _GEN6874;
wire  _GEN13157 = io_x[38] ? _GEN7036 : _GEN13156;
wire  _GEN13158 = io_x[10] ? _GEN13157 : _GEN13149;
wire  _GEN13159 = io_x[71] ? _GEN13158 : _GEN13148;
wire  _GEN13160 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN13161 = io_x[14] ? _GEN6843 : _GEN13160;
wire  _GEN13162 = io_x[0] ? _GEN13161 : _GEN6845;
wire  _GEN13163 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13164 = io_x[41] ? _GEN6836 : _GEN13163;
wire  _GEN13165 = io_x[14] ? _GEN6856 : _GEN13164;
wire  _GEN13166 = io_x[0] ? _GEN13165 : _GEN6858;
wire  _GEN13167 = io_x[76] ? _GEN13166 : _GEN13162;
wire  _GEN13168 = io_x[42] ? _GEN13167 : _GEN6874;
wire  _GEN13169 = io_x[38] ? _GEN7036 : _GEN13168;
wire  _GEN13170 = io_x[10] ? _GEN7044 : _GEN13169;
wire  _GEN13171 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13172 = io_x[0] ? _GEN13171 : _GEN6845;
wire  _GEN13173 = io_x[76] ? _GEN13172 : _GEN6834;
wire  _GEN13174 = io_x[42] ? _GEN13173 : _GEN6874;
wire  _GEN13175 = io_x[38] ? _GEN13174 : _GEN6871;
wire  _GEN13176 = io_x[10] ? _GEN7044 : _GEN13175;
wire  _GEN13177 = io_x[71] ? _GEN13176 : _GEN13170;
wire  _GEN13178 = io_x[70] ? _GEN13177 : _GEN13159;
wire  _GEN13179 = io_x[33] ? _GEN12627 : _GEN13178;
wire  _GEN13180 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN13181 = io_x[6] ? _GEN13180 : _GEN6850;
wire  _GEN13182 = io_x[41] ? _GEN6836 : _GEN13181;
wire  _GEN13183 = io_x[14] ? _GEN6856 : _GEN13182;
wire  _GEN13184 = io_x[0] ? _GEN13183 : _GEN6845;
wire  _GEN13185 = io_x[76] ? _GEN6834 : _GEN13184;
wire  _GEN13186 = io_x[42] ? _GEN13185 : _GEN6874;
wire  _GEN13187 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN13188 = io_x[38] ? _GEN13187 : _GEN13186;
wire  _GEN13189 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13190 = io_x[0] ? _GEN6845 : _GEN13189;
wire  _GEN13191 = io_x[76] ? _GEN6834 : _GEN13190;
wire  _GEN13192 = io_x[42] ? _GEN6874 : _GEN13191;
wire  _GEN13193 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN13194 = io_x[38] ? _GEN13193 : _GEN13192;
wire  _GEN13195 = io_x[10] ? _GEN13194 : _GEN13188;
wire  _GEN13196 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN13197 = io_x[76] ? _GEN13196 : _GEN6833;
wire  _GEN13198 = io_x[42] ? _GEN13197 : _GEN6874;
wire  _GEN13199 = io_x[38] ? _GEN13198 : _GEN7036;
wire  _GEN13200 = io_x[10] ? _GEN7044 : _GEN13199;
wire  _GEN13201 = io_x[71] ? _GEN13200 : _GEN13195;
wire  _GEN13202 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13203 = io_x[41] ? _GEN6836 : _GEN13202;
wire  _GEN13204 = io_x[14] ? _GEN13203 : _GEN6843;
wire  _GEN13205 = io_x[0] ? _GEN13204 : _GEN6858;
wire  _GEN13206 = io_x[76] ? _GEN6833 : _GEN13205;
wire  _GEN13207 = io_x[42] ? _GEN13206 : _GEN6874;
wire  _GEN13208 = io_x[38] ? _GEN6871 : _GEN13207;
wire  _GEN13209 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13210 = io_x[0] ? _GEN6845 : _GEN13209;
wire  _GEN13211 = io_x[76] ? _GEN6833 : _GEN13210;
wire  _GEN13212 = io_x[42] ? _GEN13211 : _GEN6874;
wire  _GEN13213 = io_x[38] ? _GEN7036 : _GEN13212;
wire  _GEN13214 = io_x[10] ? _GEN13213 : _GEN13208;
wire  _GEN13215 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN13216 = io_x[42] ? _GEN13215 : _GEN6874;
wire  _GEN13217 = io_x[38] ? _GEN7036 : _GEN13216;
wire  _GEN13218 = io_x[10] ? _GEN7094 : _GEN13217;
wire  _GEN13219 = io_x[71] ? _GEN13218 : _GEN13214;
wire  _GEN13220 = io_x[70] ? _GEN13219 : _GEN13201;
wire  _GEN13221 = io_x[33] ? _GEN12627 : _GEN13220;
wire  _GEN13222 = io_x[21] ? _GEN13221 : _GEN13179;
wire  _GEN13223 = io_x[18] ? _GEN13222 : _GEN13122;
wire  _GEN13224 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN13225 = io_x[76] ? _GEN13224 : _GEN6834;
wire  _GEN13226 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN13227 = io_x[6] ? _GEN6850 : _GEN13226;
wire  _GEN13228 = io_x[41] ? _GEN6836 : _GEN13227;
wire  _GEN13229 = io_x[14] ? _GEN13228 : _GEN6856;
wire  _GEN13230 = io_x[0] ? _GEN13229 : _GEN6858;
wire  _GEN13231 = io_x[76] ? _GEN6834 : _GEN13230;
wire  _GEN13232 = io_x[42] ? _GEN13231 : _GEN13225;
wire  _GEN13233 = io_x[38] ? _GEN6871 : _GEN13232;
wire  _GEN13234 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN13235 = io_x[14] ? _GEN6843 : _GEN13234;
wire  _GEN13236 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN13237 = io_x[6] ? _GEN6850 : _GEN13236;
wire  _GEN13238 = io_x[41] ? _GEN6836 : _GEN13237;
wire  _GEN13239 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13240 = io_x[41] ? _GEN6836 : _GEN13239;
wire  _GEN13241 = io_x[14] ? _GEN13240 : _GEN13238;
wire  _GEN13242 = io_x[0] ? _GEN13241 : _GEN13235;
wire  _GEN13243 = io_x[76] ? _GEN6834 : _GEN13242;
wire  _GEN13244 = io_x[42] ? _GEN13243 : _GEN6874;
wire  _GEN13245 = io_x[38] ? _GEN6871 : _GEN13244;
wire  _GEN13246 = io_x[10] ? _GEN13245 : _GEN13233;
wire  _GEN13247 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13248 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13249 = io_x[41] ? _GEN6924 : _GEN13248;
wire  _GEN13250 = io_x[14] ? _GEN6856 : _GEN13249;
wire  _GEN13251 = io_x[0] ? _GEN13250 : _GEN13247;
wire  _GEN13252 = io_x[76] ? _GEN6834 : _GEN13251;
wire  _GEN13253 = io_x[42] ? _GEN13252 : _GEN6874;
wire  _GEN13254 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13255 = io_x[0] ? _GEN6845 : _GEN13254;
wire  _GEN13256 = io_x[76] ? _GEN13255 : _GEN6834;
wire  _GEN13257 = io_x[42] ? _GEN13256 : _GEN6874;
wire  _GEN13258 = io_x[38] ? _GEN13257 : _GEN13253;
wire  _GEN13259 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13260 = io_x[0] ? _GEN6845 : _GEN13259;
wire  _GEN13261 = io_x[76] ? _GEN6833 : _GEN13260;
wire  _GEN13262 = io_x[42] ? _GEN6874 : _GEN13261;
wire  _GEN13263 = io_x[38] ? _GEN7036 : _GEN13262;
wire  _GEN13264 = io_x[10] ? _GEN13263 : _GEN13258;
wire  _GEN13265 = io_x[71] ? _GEN13264 : _GEN13246;
wire  _GEN13266 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13267 = io_x[41] ? _GEN6836 : _GEN13266;
wire  _GEN13268 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN13269 = io_x[6] ? _GEN13268 : _GEN6850;
wire  _GEN13270 = io_x[41] ? _GEN6836 : _GEN13269;
wire  _GEN13271 = io_x[14] ? _GEN13270 : _GEN13267;
wire  _GEN13272 = io_x[0] ? _GEN6845 : _GEN13271;
wire  _GEN13273 = io_x[76] ? _GEN13272 : _GEN6834;
wire  _GEN13274 = io_x[42] ? _GEN13273 : _GEN6874;
wire  _GEN13275 = io_x[38] ? _GEN13274 : _GEN6871;
wire  _GEN13276 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN13277 = io_x[38] ? _GEN7036 : _GEN13276;
wire  _GEN13278 = io_x[10] ? _GEN13277 : _GEN13275;
wire  _GEN13279 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN13280 = io_x[14] ? _GEN6843 : _GEN13279;
wire  _GEN13281 = io_x[0] ? _GEN6845 : _GEN13280;
wire  _GEN13282 = io_x[76] ? _GEN13281 : _GEN6834;
wire  _GEN13283 = io_x[42] ? _GEN13282 : _GEN6874;
wire  _GEN13284 = io_x[38] ? _GEN13283 : _GEN7036;
wire  _GEN13285 = io_x[10] ? _GEN7094 : _GEN13284;
wire  _GEN13286 = io_x[71] ? _GEN13285 : _GEN13278;
wire  _GEN13287 = io_x[70] ? _GEN13286 : _GEN13265;
wire  _GEN13288 = io_x[33] ? _GEN12627 : _GEN13287;
wire  _GEN13289 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13290 = io_x[41] ? _GEN13289 : _GEN6924;
wire  _GEN13291 = io_x[14] ? _GEN6843 : _GEN13290;
wire  _GEN13292 = io_x[0] ? _GEN6845 : _GEN13291;
wire  _GEN13293 = io_x[76] ? _GEN6833 : _GEN13292;
wire  _GEN13294 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13295 = io_x[6] ? _GEN6850 : _GEN13294;
wire  _GEN13296 = io_x[41] ? _GEN6836 : _GEN13295;
wire  _GEN13297 = io_x[14] ? _GEN6843 : _GEN13296;
wire  _GEN13298 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13299 = io_x[6] ? _GEN13298 : _GEN6850;
wire  _GEN13300 = io_x[41] ? _GEN6836 : _GEN13299;
wire  _GEN13301 = io_x[14] ? _GEN13300 : _GEN6856;
wire  _GEN13302 = io_x[0] ? _GEN13301 : _GEN13297;
wire  _GEN13303 = io_x[76] ? _GEN6833 : _GEN13302;
wire  _GEN13304 = io_x[42] ? _GEN13303 : _GEN13293;
wire  _GEN13305 = io_x[38] ? _GEN7036 : _GEN13304;
wire  _GEN13306 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13307 = io_x[41] ? _GEN6836 : _GEN13306;
wire  _GEN13308 = io_x[14] ? _GEN13307 : _GEN6843;
wire  _GEN13309 = io_x[0] ? _GEN13308 : _GEN6845;
wire  _GEN13310 = io_x[76] ? _GEN6834 : _GEN13309;
wire  _GEN13311 = io_x[42] ? _GEN13310 : _GEN6874;
wire  _GEN13312 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13313 = io_x[0] ? _GEN13312 : _GEN6845;
wire  _GEN13314 = io_x[76] ? _GEN13313 : _GEN6834;
wire  _GEN13315 = io_x[42] ? _GEN6874 : _GEN13314;
wire  _GEN13316 = io_x[38] ? _GEN13315 : _GEN13311;
wire  _GEN13317 = io_x[10] ? _GEN13316 : _GEN13305;
wire  _GEN13318 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13319 = io_x[0] ? _GEN6845 : _GEN13318;
wire  _GEN13320 = io_x[76] ? _GEN13319 : _GEN6834;
wire  _GEN13321 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13322 = io_x[41] ? _GEN6836 : _GEN13321;
wire  _GEN13323 = io_x[14] ? _GEN6843 : _GEN13322;
wire  _GEN13324 = io_x[0] ? _GEN6845 : _GEN13323;
wire  _GEN13325 = io_x[76] ? _GEN6834 : _GEN13324;
wire  _GEN13326 = io_x[42] ? _GEN13325 : _GEN13320;
wire  _GEN13327 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13328 = io_x[41] ? _GEN13327 : _GEN6836;
wire  _GEN13329 = io_x[14] ? _GEN6843 : _GEN13328;
wire  _GEN13330 = io_x[0] ? _GEN6845 : _GEN13329;
wire  _GEN13331 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13332 = io_x[0] ? _GEN6845 : _GEN13331;
wire  _GEN13333 = io_x[76] ? _GEN13332 : _GEN13330;
wire  _GEN13334 = io_x[42] ? _GEN13333 : _GEN6874;
wire  _GEN13335 = io_x[38] ? _GEN13334 : _GEN13326;
wire  _GEN13336 = io_x[10] ? _GEN7094 : _GEN13335;
wire  _GEN13337 = io_x[71] ? _GEN13336 : _GEN13317;
wire  _GEN13338 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN13339 = io_x[42] ? _GEN13338 : _GEN6874;
wire  _GEN13340 = io_x[38] ? _GEN7036 : _GEN13339;
wire  _GEN13341 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13342 = io_x[0] ? _GEN6845 : _GEN13341;
wire  _GEN13343 = io_x[76] ? _GEN13342 : _GEN6834;
wire  _GEN13344 = io_x[42] ? _GEN6874 : _GEN13343;
wire  _GEN13345 = io_x[38] ? _GEN7036 : _GEN13344;
wire  _GEN13346 = io_x[10] ? _GEN13345 : _GEN13340;
wire  _GEN13347 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN13348 = io_x[38] ? _GEN13347 : _GEN6871;
wire  _GEN13349 = io_x[10] ? _GEN7044 : _GEN13348;
wire  _GEN13350 = io_x[71] ? _GEN13349 : _GEN13346;
wire  _GEN13351 = io_x[70] ? _GEN13350 : _GEN13337;
wire  _GEN13352 = io_x[33] ? _GEN12627 : _GEN13351;
wire  _GEN13353 = io_x[21] ? _GEN13352 : _GEN13288;
wire  _GEN13354 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13355 = io_x[41] ? _GEN13354 : _GEN6924;
wire  _GEN13356 = io_x[14] ? _GEN6843 : _GEN13355;
wire  _GEN13357 = io_x[0] ? _GEN13356 : _GEN6858;
wire  _GEN13358 = io_x[76] ? _GEN6833 : _GEN13357;
wire  _GEN13359 = io_x[42] ? _GEN13358 : _GEN6874;
wire  _GEN13360 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13361 = io_x[6] ? _GEN6850 : _GEN13360;
wire  _GEN13362 = io_x[41] ? _GEN13361 : _GEN6836;
wire  _GEN13363 = io_x[14] ? _GEN6843 : _GEN13362;
wire  _GEN13364 = io_x[0] ? _GEN13363 : _GEN6845;
wire  _GEN13365 = io_x[76] ? _GEN6834 : _GEN13364;
wire  _GEN13366 = io_x[42] ? _GEN13365 : _GEN6874;
wire  _GEN13367 = io_x[38] ? _GEN13366 : _GEN13359;
wire  _GEN13368 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13369 = io_x[0] ? _GEN13368 : _GEN6845;
wire  _GEN13370 = io_x[76] ? _GEN13369 : _GEN6834;
wire  _GEN13371 = io_x[42] ? _GEN6874 : _GEN13370;
wire  _GEN13372 = io_x[38] ? _GEN13371 : _GEN6871;
wire  _GEN13373 = io_x[10] ? _GEN13372 : _GEN13367;
wire  _GEN13374 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13375 = io_x[0] ? _GEN13374 : _GEN6858;
wire  _GEN13376 = io_x[76] ? _GEN6834 : _GEN13375;
wire  _GEN13377 = io_x[42] ? _GEN13376 : _GEN6874;
wire  _GEN13378 = io_x[38] ? _GEN6871 : _GEN13377;
wire  _GEN13379 = io_x[10] ? _GEN7044 : _GEN13378;
wire  _GEN13380 = io_x[71] ? _GEN13379 : _GEN13373;
wire  _GEN13381 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13382 = io_x[0] ? _GEN13381 : _GEN6845;
wire  _GEN13383 = io_x[76] ? _GEN13382 : _GEN6834;
wire  _GEN13384 = io_x[42] ? _GEN13383 : _GEN6874;
wire  _GEN13385 = io_x[38] ? _GEN6871 : _GEN13384;
wire  _GEN13386 = io_x[10] ? _GEN7094 : _GEN13385;
wire  _GEN13387 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13388 = io_x[6] ? _GEN6850 : _GEN13387;
wire  _GEN13389 = io_x[41] ? _GEN6836 : _GEN13388;
wire  _GEN13390 = io_x[14] ? _GEN13389 : _GEN6843;
wire  _GEN13391 = io_x[0] ? _GEN13390 : _GEN6845;
wire  _GEN13392 = io_x[76] ? _GEN13391 : _GEN6834;
wire  _GEN13393 = io_x[42] ? _GEN13392 : _GEN6874;
wire  _GEN13394 = io_x[38] ? _GEN13393 : _GEN6871;
wire  _GEN13395 = io_x[10] ? _GEN7044 : _GEN13394;
wire  _GEN13396 = io_x[71] ? _GEN13395 : _GEN13386;
wire  _GEN13397 = io_x[70] ? _GEN13396 : _GEN13380;
wire  _GEN13398 = io_x[33] ? _GEN12641 : _GEN13397;
wire  _GEN13399 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN13400 = io_x[6] ? _GEN13399 : _GEN6850;
wire  _GEN13401 = io_x[41] ? _GEN6836 : _GEN13400;
wire  _GEN13402 = io_x[14] ? _GEN6856 : _GEN13401;
wire  _GEN13403 = io_x[0] ? _GEN13402 : _GEN6845;
wire  _GEN13404 = io_x[76] ? _GEN6834 : _GEN13403;
wire  _GEN13405 = io_x[42] ? _GEN13404 : _GEN6874;
wire  _GEN13406 = io_x[38] ? _GEN7036 : _GEN13405;
wire  _GEN13407 = io_x[10] ? _GEN7094 : _GEN13406;
wire  _GEN13408 = io_x[71] ? _GEN7203 : _GEN13407;
wire  _GEN13409 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN13410 = io_x[14] ? _GEN6843 : _GEN13409;
wire  _GEN13411 = io_x[0] ? _GEN6845 : _GEN13410;
wire  _GEN13412 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13413 = io_x[0] ? _GEN6845 : _GEN13412;
wire  _GEN13414 = io_x[76] ? _GEN13413 : _GEN13411;
wire  _GEN13415 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13416 = io_x[0] ? _GEN13415 : _GEN6845;
wire  _GEN13417 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13418 = io_x[41] ? _GEN6836 : _GEN13417;
wire  _GEN13419 = io_x[14] ? _GEN13418 : _GEN6843;
wire  _GEN13420 = io_x[0] ? _GEN13419 : _GEN6845;
wire  _GEN13421 = io_x[76] ? _GEN13420 : _GEN13416;
wire  _GEN13422 = io_x[42] ? _GEN13421 : _GEN13414;
wire  _GEN13423 = io_x[38] ? _GEN6871 : _GEN13422;
wire  _GEN13424 = io_x[10] ? _GEN7044 : _GEN13423;
wire  _GEN13425 = io_x[71] ? _GEN7196 : _GEN13424;
wire  _GEN13426 = io_x[70] ? _GEN13425 : _GEN13408;
wire  _GEN13427 = io_x[33] ? _GEN12627 : _GEN13426;
wire  _GEN13428 = io_x[21] ? _GEN13427 : _GEN13398;
wire  _GEN13429 = io_x[18] ? _GEN13428 : _GEN13353;
wire  _GEN13430 = io_x[20] ? _GEN13429 : _GEN13223;
wire  _GEN13431 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN13432 = io_x[14] ? _GEN6843 : _GEN13431;
wire  _GEN13433 = io_x[0] ? _GEN6845 : _GEN13432;
wire  _GEN13434 = io_x[76] ? _GEN6834 : _GEN13433;
wire  _GEN13435 = io_x[42] ? _GEN6874 : _GEN13434;
wire  _GEN13436 = io_x[38] ? _GEN13435 : _GEN6871;
wire  _GEN13437 = io_x[10] ? _GEN7044 : _GEN13436;
wire  _GEN13438 = io_x[71] ? _GEN7196 : _GEN13437;
wire  _GEN13439 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN13440 = io_x[10] ? _GEN7044 : _GEN13439;
wire  _GEN13441 = io_x[71] ? _GEN7203 : _GEN13440;
wire  _GEN13442 = io_x[70] ? _GEN13441 : _GEN13438;
wire  _GEN13443 = io_x[33] ? _GEN12627 : _GEN13442;
wire  _GEN13444 = io_x[21] ? _GEN12643 : _GEN13443;
wire  _GEN13445 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN13446 = io_x[76] ? _GEN13445 : _GEN6834;
wire  _GEN13447 = io_x[42] ? _GEN6874 : _GEN13446;
wire  _GEN13448 = io_x[38] ? _GEN6871 : _GEN13447;
wire  _GEN13449 = io_x[10] ? _GEN7094 : _GEN13448;
wire  _GEN13450 = io_x[71] ? _GEN7196 : _GEN13449;
wire  _GEN13451 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN13452 = io_x[38] ? _GEN6871 : _GEN13451;
wire  _GEN13453 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN13454 = io_x[10] ? _GEN13453 : _GEN13452;
wire  _GEN13455 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN13456 = io_x[10] ? _GEN7044 : _GEN13455;
wire  _GEN13457 = io_x[71] ? _GEN13456 : _GEN13454;
wire  _GEN13458 = io_x[70] ? _GEN13457 : _GEN13450;
wire  _GEN13459 = io_x[33] ? _GEN12627 : _GEN13458;
wire  _GEN13460 = io_x[21] ? _GEN12643 : _GEN13459;
wire  _GEN13461 = io_x[18] ? _GEN13460 : _GEN13444;
wire  _GEN13462 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13463 = io_x[41] ? _GEN6836 : _GEN13462;
wire  _GEN13464 = io_x[14] ? _GEN13463 : _GEN6843;
wire  _GEN13465 = io_x[0] ? _GEN13464 : _GEN6845;
wire  _GEN13466 = io_x[76] ? _GEN13465 : _GEN6834;
wire  _GEN13467 = io_x[42] ? _GEN6863 : _GEN13466;
wire  _GEN13468 = io_x[38] ? _GEN6871 : _GEN13467;
wire  _GEN13469 = io_x[10] ? _GEN13468 : _GEN7094;
wire  _GEN13470 = io_x[71] ? _GEN7196 : _GEN13469;
wire  _GEN13471 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN13472 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13473 = io_x[41] ? _GEN13472 : _GEN6836;
wire  _GEN13474 = io_x[14] ? _GEN13473 : _GEN6843;
wire  _GEN13475 = io_x[0] ? _GEN6845 : _GEN13474;
wire  _GEN13476 = io_x[76] ? _GEN13475 : _GEN6834;
wire  _GEN13477 = io_x[42] ? _GEN6874 : _GEN13476;
wire  _GEN13478 = io_x[38] ? _GEN6871 : _GEN13477;
wire  _GEN13479 = io_x[10] ? _GEN7044 : _GEN13478;
wire  _GEN13480 = io_x[71] ? _GEN13479 : _GEN13471;
wire  _GEN13481 = io_x[70] ? _GEN13480 : _GEN13470;
wire  _GEN13482 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13483 = io_x[41] ? _GEN13482 : _GEN6836;
wire  _GEN13484 = io_x[14] ? _GEN13483 : _GEN6843;
wire  _GEN13485 = io_x[0] ? _GEN6845 : _GEN13484;
wire  _GEN13486 = io_x[76] ? _GEN13485 : _GEN6834;
wire  _GEN13487 = io_x[42] ? _GEN6874 : _GEN13486;
wire  _GEN13488 = io_x[38] ? _GEN6871 : _GEN13487;
wire  _GEN13489 = io_x[10] ? _GEN7044 : _GEN13488;
wire  _GEN13490 = io_x[71] ? _GEN7196 : _GEN13489;
wire  _GEN13491 = io_x[70] ? _GEN8474 : _GEN13490;
wire  _GEN13492 = io_x[33] ? _GEN13491 : _GEN13481;
wire  _GEN13493 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13494 = io_x[0] ? _GEN13493 : _GEN6845;
wire  _GEN13495 = io_x[76] ? _GEN6834 : _GEN13494;
wire  _GEN13496 = io_x[42] ? _GEN6874 : _GEN13495;
wire  _GEN13497 = io_x[38] ? _GEN13496 : _GEN7036;
wire  _GEN13498 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN13499 = io_x[42] ? _GEN6874 : _GEN13498;
wire  _GEN13500 = io_x[38] ? _GEN6871 : _GEN13499;
wire  _GEN13501 = io_x[10] ? _GEN13500 : _GEN13497;
wire  _GEN13502 = io_x[71] ? _GEN7196 : _GEN13501;
wire  _GEN13503 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13504 = io_x[0] ? _GEN13503 : _GEN6845;
wire  _GEN13505 = io_x[76] ? _GEN13504 : _GEN6834;
wire  _GEN13506 = io_x[42] ? _GEN6874 : _GEN13505;
wire  _GEN13507 = io_x[38] ? _GEN6871 : _GEN13506;
wire  _GEN13508 = io_x[10] ? _GEN7044 : _GEN13507;
wire  _GEN13509 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN13510 = io_x[71] ? _GEN13509 : _GEN13508;
wire  _GEN13511 = io_x[70] ? _GEN13510 : _GEN13502;
wire  _GEN13512 = io_x[71] ? _GEN7196 : _GEN7203;
wire  _GEN13513 = io_x[70] ? _GEN13512 : _GEN8474;
wire  _GEN13514 = io_x[33] ? _GEN13513 : _GEN13511;
wire  _GEN13515 = io_x[21] ? _GEN13514 : _GEN13492;
wire  _GEN13516 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN13517 = io_x[10] ? _GEN7094 : _GEN13516;
wire  _GEN13518 = io_x[71] ? _GEN7203 : _GEN13517;
wire  _GEN13519 = io_x[70] ? _GEN8474 : _GEN13518;
wire  _GEN13520 = io_x[33] ? _GEN12627 : _GEN13519;
wire  _GEN13521 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13522 = io_x[41] ? _GEN6836 : _GEN13521;
wire  _GEN13523 = io_x[14] ? _GEN13522 : _GEN6843;
wire  _GEN13524 = io_x[0] ? _GEN13523 : _GEN6845;
wire  _GEN13525 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN13526 = io_x[14] ? _GEN6843 : _GEN13525;
wire  _GEN13527 = io_x[0] ? _GEN6845 : _GEN13526;
wire  _GEN13528 = io_x[76] ? _GEN13527 : _GEN13524;
wire  _GEN13529 = io_x[42] ? _GEN6874 : _GEN13528;
wire  _GEN13530 = io_x[38] ? _GEN13529 : _GEN7036;
wire  _GEN13531 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN13532 = io_x[14] ? _GEN13531 : _GEN6843;
wire  _GEN13533 = io_x[0] ? _GEN13532 : _GEN6845;
wire  _GEN13534 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN13535 = io_x[6] ? _GEN13534 : _GEN6850;
wire  _GEN13536 = io_x[41] ? _GEN13535 : _GEN6836;
wire  _GEN13537 = io_x[14] ? _GEN6856 : _GEN13536;
wire  _GEN13538 = io_x[0] ? _GEN13537 : _GEN6845;
wire  _GEN13539 = io_x[76] ? _GEN13538 : _GEN13533;
wire  _GEN13540 = io_x[42] ? _GEN6874 : _GEN13539;
wire  _GEN13541 = io_x[38] ? _GEN6871 : _GEN13540;
wire  _GEN13542 = io_x[10] ? _GEN13541 : _GEN13530;
wire  _GEN13543 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13544 = io_x[41] ? _GEN13543 : _GEN6836;
wire  _GEN13545 = io_x[14] ? _GEN6843 : _GEN13544;
wire  _GEN13546 = io_x[0] ? _GEN13545 : _GEN6845;
wire  _GEN13547 = io_x[76] ? _GEN6834 : _GEN13546;
wire  _GEN13548 = io_x[42] ? _GEN6874 : _GEN13547;
wire  _GEN13549 = io_x[38] ? _GEN13548 : _GEN6871;
wire  _GEN13550 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13551 = io_x[41] ? _GEN13550 : _GEN6836;
wire  _GEN13552 = io_x[14] ? _GEN13551 : _GEN6843;
wire  _GEN13553 = io_x[0] ? _GEN6845 : _GEN13552;
wire  _GEN13554 = io_x[76] ? _GEN13553 : _GEN6834;
wire  _GEN13555 = io_x[42] ? _GEN6874 : _GEN13554;
wire  _GEN13556 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN13557 = io_x[42] ? _GEN6874 : _GEN13556;
wire  _GEN13558 = io_x[38] ? _GEN13557 : _GEN13555;
wire  _GEN13559 = io_x[10] ? _GEN13558 : _GEN13549;
wire  _GEN13560 = io_x[71] ? _GEN13559 : _GEN13542;
wire  _GEN13561 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13562 = io_x[41] ? _GEN13561 : _GEN6836;
wire  _GEN13563 = io_x[14] ? _GEN6843 : _GEN13562;
wire  _GEN13564 = io_x[0] ? _GEN13563 : _GEN6845;
wire  _GEN13565 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13566 = io_x[41] ? _GEN13565 : _GEN6836;
wire  _GEN13567 = io_x[14] ? _GEN13566 : _GEN6843;
wire  _GEN13568 = io_x[0] ? _GEN13567 : _GEN6845;
wire  _GEN13569 = io_x[76] ? _GEN13568 : _GEN13564;
wire  _GEN13570 = io_x[42] ? _GEN6874 : _GEN13569;
wire  _GEN13571 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13572 = io_x[41] ? _GEN6836 : _GEN13571;
wire  _GEN13573 = io_x[14] ? _GEN13572 : _GEN6843;
wire  _GEN13574 = io_x[0] ? _GEN13573 : _GEN6845;
wire  _GEN13575 = io_x[76] ? _GEN13574 : _GEN6834;
wire  _GEN13576 = io_x[42] ? _GEN6874 : _GEN13575;
wire  _GEN13577 = io_x[38] ? _GEN13576 : _GEN13570;
wire  _GEN13578 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13579 = io_x[41] ? _GEN13578 : _GEN6836;
wire  _GEN13580 = io_x[14] ? _GEN13579 : _GEN6843;
wire  _GEN13581 = io_x[0] ? _GEN13580 : _GEN6845;
wire  _GEN13582 = io_x[76] ? _GEN13581 : _GEN6834;
wire  _GEN13583 = io_x[42] ? _GEN6874 : _GEN13582;
wire  _GEN13584 = io_x[38] ? _GEN6871 : _GEN13583;
wire  _GEN13585 = io_x[10] ? _GEN13584 : _GEN13577;
wire  _GEN13586 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN13587 = io_x[76] ? _GEN13586 : _GEN6834;
wire  _GEN13588 = io_x[42] ? _GEN6874 : _GEN13587;
wire  _GEN13589 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13590 = io_x[41] ? _GEN13589 : _GEN6836;
wire  _GEN13591 = io_x[14] ? _GEN6843 : _GEN13590;
wire  _GEN13592 = io_x[0] ? _GEN13591 : _GEN6845;
wire  _GEN13593 = io_x[76] ? _GEN6834 : _GEN13592;
wire  _GEN13594 = io_x[42] ? _GEN6874 : _GEN13593;
wire  _GEN13595 = io_x[38] ? _GEN13594 : _GEN13588;
wire  _GEN13596 = io_x[10] ? _GEN7044 : _GEN13595;
wire  _GEN13597 = io_x[71] ? _GEN13596 : _GEN13585;
wire  _GEN13598 = io_x[70] ? _GEN13597 : _GEN13560;
wire  _GEN13599 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13600 = io_x[41] ? _GEN6836 : _GEN13599;
wire  _GEN13601 = io_x[14] ? _GEN13600 : _GEN6843;
wire  _GEN13602 = io_x[0] ? _GEN13601 : _GEN6845;
wire  _GEN13603 = io_x[76] ? _GEN6833 : _GEN13602;
wire  _GEN13604 = io_x[42] ? _GEN6874 : _GEN13603;
wire  _GEN13605 = io_x[38] ? _GEN6871 : _GEN13604;
wire  _GEN13606 = io_x[10] ? _GEN7044 : _GEN13605;
wire  _GEN13607 = io_x[71] ? _GEN7196 : _GEN13606;
wire  _GEN13608 = io_x[70] ? _GEN8474 : _GEN13607;
wire  _GEN13609 = io_x[33] ? _GEN13608 : _GEN13598;
wire  _GEN13610 = io_x[21] ? _GEN13609 : _GEN13520;
wire  _GEN13611 = io_x[18] ? _GEN13610 : _GEN13515;
wire  _GEN13612 = io_x[20] ? _GEN13611 : _GEN13461;
wire  _GEN13613 = io_x[45] ? _GEN13612 : _GEN13430;
wire  _GEN13614 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13615 = io_x[6] ? _GEN6850 : _GEN13614;
wire  _GEN13616 = io_x[41] ? _GEN13615 : _GEN6836;
wire  _GEN13617 = io_x[14] ? _GEN6843 : _GEN13616;
wire  _GEN13618 = io_x[0] ? _GEN13617 : _GEN6845;
wire  _GEN13619 = io_x[76] ? _GEN13618 : _GEN6834;
wire  _GEN13620 = io_x[42] ? _GEN13619 : _GEN6874;
wire  _GEN13621 = io_x[38] ? _GEN6871 : _GEN13620;
wire  _GEN13622 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13623 = io_x[0] ? _GEN6845 : _GEN13622;
wire  _GEN13624 = io_x[76] ? _GEN13623 : _GEN6833;
wire  _GEN13625 = io_x[42] ? _GEN13624 : _GEN6874;
wire  _GEN13626 = io_x[38] ? _GEN7036 : _GEN13625;
wire  _GEN13627 = io_x[10] ? _GEN13626 : _GEN13621;
wire  _GEN13628 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN13629 = io_x[6] ? _GEN13628 : _GEN6850;
wire  _GEN13630 = io_x[41] ? _GEN13629 : _GEN6836;
wire  _GEN13631 = io_x[14] ? _GEN6843 : _GEN13630;
wire  _GEN13632 = io_x[0] ? _GEN13631 : _GEN6845;
wire  _GEN13633 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13634 = io_x[41] ? _GEN6836 : _GEN13633;
wire  _GEN13635 = io_x[14] ? _GEN13634 : _GEN6843;
wire  _GEN13636 = io_x[0] ? _GEN6845 : _GEN13635;
wire  _GEN13637 = io_x[76] ? _GEN13636 : _GEN13632;
wire  _GEN13638 = io_x[42] ? _GEN13637 : _GEN6874;
wire  _GEN13639 = io_x[38] ? _GEN13638 : _GEN6871;
wire  _GEN13640 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN13641 = io_x[14] ? _GEN13640 : _GEN6856;
wire  _GEN13642 = io_x[0] ? _GEN6845 : _GEN13641;
wire  _GEN13643 = io_x[76] ? _GEN13642 : _GEN6834;
wire  _GEN13644 = io_x[42] ? _GEN13643 : _GEN6874;
wire  _GEN13645 = io_x[38] ? _GEN13644 : _GEN7036;
wire  _GEN13646 = io_x[10] ? _GEN13645 : _GEN13639;
wire  _GEN13647 = io_x[71] ? _GEN13646 : _GEN13627;
wire  _GEN13648 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13649 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13650 = io_x[6] ? _GEN6840 : _GEN13649;
wire  _GEN13651 = io_x[41] ? _GEN6836 : _GEN13650;
wire  _GEN13652 = io_x[14] ? _GEN13651 : _GEN6843;
wire  _GEN13653 = io_x[0] ? _GEN13652 : _GEN13648;
wire  _GEN13654 = io_x[76] ? _GEN13653 : _GEN6833;
wire  _GEN13655 = io_x[42] ? _GEN13654 : _GEN6874;
wire  _GEN13656 = io_x[38] ? _GEN7036 : _GEN13655;
wire  _GEN13657 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13658 = io_x[0] ? _GEN6845 : _GEN13657;
wire  _GEN13659 = io_x[76] ? _GEN13658 : _GEN6834;
wire  _GEN13660 = io_x[42] ? _GEN13659 : _GEN6874;
wire  _GEN13661 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN13662 = io_x[76] ? _GEN13661 : _GEN6834;
wire  _GEN13663 = io_x[42] ? _GEN13662 : _GEN6874;
wire  _GEN13664 = io_x[38] ? _GEN13663 : _GEN13660;
wire  _GEN13665 = io_x[10] ? _GEN13664 : _GEN13656;
wire  _GEN13666 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN13667 = io_x[76] ? _GEN13666 : _GEN6834;
wire  _GEN13668 = io_x[42] ? _GEN13667 : _GEN6874;
wire  _GEN13669 = io_x[38] ? _GEN13668 : _GEN6871;
wire  _GEN13670 = io_x[10] ? _GEN13669 : _GEN7094;
wire  _GEN13671 = io_x[71] ? _GEN13670 : _GEN13665;
wire  _GEN13672 = io_x[70] ? _GEN13671 : _GEN13647;
wire  _GEN13673 = io_x[70] ? _GEN7020 : _GEN8474;
wire  _GEN13674 = io_x[33] ? _GEN13673 : _GEN13672;
wire  _GEN13675 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN13676 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN13677 = io_x[10] ? _GEN7044 : _GEN13676;
wire  _GEN13678 = io_x[71] ? _GEN13677 : _GEN13675;
wire  _GEN13679 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN13680 = io_x[10] ? _GEN13679 : _GEN7094;
wire  _GEN13681 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN13682 = io_x[71] ? _GEN13681 : _GEN13680;
wire  _GEN13683 = io_x[70] ? _GEN13682 : _GEN13678;
wire  _GEN13684 = io_x[33] ? _GEN12641 : _GEN13683;
wire  _GEN13685 = io_x[21] ? _GEN13684 : _GEN13674;
wire  _GEN13686 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13687 = io_x[41] ? _GEN6836 : _GEN13686;
wire  _GEN13688 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13689 = io_x[41] ? _GEN6924 : _GEN13688;
wire  _GEN13690 = io_x[14] ? _GEN13689 : _GEN13687;
wire  _GEN13691 = io_x[0] ? _GEN13690 : _GEN6845;
wire  _GEN13692 = io_x[76] ? _GEN6834 : _GEN13691;
wire  _GEN13693 = io_x[42] ? _GEN13692 : _GEN6874;
wire  _GEN13694 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13695 = io_x[6] ? _GEN6850 : _GEN13694;
wire  _GEN13696 = io_x[41] ? _GEN13695 : _GEN6836;
wire  _GEN13697 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13698 = io_x[41] ? _GEN13697 : _GEN6836;
wire  _GEN13699 = io_x[14] ? _GEN13698 : _GEN13696;
wire  _GEN13700 = io_x[0] ? _GEN13699 : _GEN6845;
wire  _GEN13701 = io_x[76] ? _GEN13700 : _GEN6834;
wire  _GEN13702 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13703 = io_x[0] ? _GEN13702 : _GEN6845;
wire  _GEN13704 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13705 = io_x[0] ? _GEN13704 : _GEN6845;
wire  _GEN13706 = io_x[76] ? _GEN13705 : _GEN13703;
wire  _GEN13707 = io_x[42] ? _GEN13706 : _GEN13701;
wire  _GEN13708 = io_x[38] ? _GEN13707 : _GEN13693;
wire  _GEN13709 = io_x[10] ? _GEN13708 : _GEN7094;
wire  _GEN13710 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13711 = io_x[6] ? _GEN6850 : _GEN13710;
wire  _GEN13712 = io_x[41] ? _GEN6836 : _GEN13711;
wire  _GEN13713 = io_x[14] ? _GEN6856 : _GEN13712;
wire  _GEN13714 = io_x[0] ? _GEN13713 : _GEN6845;
wire  _GEN13715 = io_x[76] ? _GEN6834 : _GEN13714;
wire  _GEN13716 = io_x[42] ? _GEN13715 : _GEN6874;
wire  _GEN13717 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN13718 = io_x[76] ? _GEN6834 : _GEN13717;
wire  _GEN13719 = io_x[42] ? _GEN13718 : _GEN6874;
wire  _GEN13720 = io_x[38] ? _GEN13719 : _GEN13716;
wire  _GEN13721 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN13722 = io_x[38] ? _GEN7036 : _GEN13721;
wire  _GEN13723 = io_x[10] ? _GEN13722 : _GEN13720;
wire  _GEN13724 = io_x[71] ? _GEN13723 : _GEN13709;
wire  _GEN13725 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN13726 = io_x[38] ? _GEN7036 : _GEN13725;
wire  _GEN13727 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13728 = io_x[41] ? _GEN6836 : _GEN13727;
wire  _GEN13729 = io_x[14] ? _GEN13728 : _GEN6843;
wire  _GEN13730 = io_x[0] ? _GEN13729 : _GEN6845;
wire  _GEN13731 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13732 = io_x[41] ? _GEN6836 : _GEN13731;
wire  _GEN13733 = io_x[14] ? _GEN6856 : _GEN13732;
wire  _GEN13734 = io_x[0] ? _GEN13733 : _GEN6858;
wire  _GEN13735 = io_x[76] ? _GEN13734 : _GEN13730;
wire  _GEN13736 = io_x[42] ? _GEN13735 : _GEN6874;
wire  _GEN13737 = io_x[38] ? _GEN7036 : _GEN13736;
wire  _GEN13738 = io_x[10] ? _GEN13737 : _GEN13726;
wire  _GEN13739 = io_x[71] ? _GEN7196 : _GEN13738;
wire  _GEN13740 = io_x[70] ? _GEN13739 : _GEN13724;
wire  _GEN13741 = io_x[33] ? _GEN12627 : _GEN13740;
wire  _GEN13742 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN13743 = io_x[42] ? _GEN6863 : _GEN13742;
wire  _GEN13744 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13745 = io_x[0] ? _GEN13744 : _GEN6845;
wire  _GEN13746 = io_x[76] ? _GEN13745 : _GEN6834;
wire  _GEN13747 = io_x[42] ? _GEN6874 : _GEN13746;
wire  _GEN13748 = io_x[38] ? _GEN13747 : _GEN13743;
wire  _GEN13749 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13750 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13751 = io_x[41] ? _GEN6924 : _GEN13750;
wire  _GEN13752 = io_x[14] ? _GEN13751 : _GEN6856;
wire  _GEN13753 = io_x[0] ? _GEN13752 : _GEN13749;
wire  _GEN13754 = io_x[76] ? _GEN6834 : _GEN13753;
wire  _GEN13755 = io_x[42] ? _GEN13754 : _GEN6863;
wire  _GEN13756 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN13757 = io_x[6] ? _GEN13756 : _GEN6850;
wire  _GEN13758 = io_x[41] ? _GEN13757 : _GEN6836;
wire  _GEN13759 = io_x[14] ? _GEN6843 : _GEN13758;
wire  _GEN13760 = io_x[0] ? _GEN13759 : _GEN6845;
wire  _GEN13761 = io_x[76] ? _GEN13760 : _GEN6834;
wire  _GEN13762 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13763 = io_x[0] ? _GEN13762 : _GEN6845;
wire  _GEN13764 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13765 = io_x[0] ? _GEN13764 : _GEN6845;
wire  _GEN13766 = io_x[76] ? _GEN13765 : _GEN13763;
wire  _GEN13767 = io_x[42] ? _GEN13766 : _GEN13761;
wire  _GEN13768 = io_x[38] ? _GEN13767 : _GEN13755;
wire  _GEN13769 = io_x[10] ? _GEN13768 : _GEN13748;
wire  _GEN13770 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN13771 = io_x[6] ? _GEN6850 : _GEN13770;
wire  _GEN13772 = io_x[41] ? _GEN6836 : _GEN13771;
wire  _GEN13773 = io_x[14] ? _GEN13772 : _GEN6856;
wire  _GEN13774 = io_x[0] ? _GEN6845 : _GEN13773;
wire  _GEN13775 = io_x[76] ? _GEN6834 : _GEN13774;
wire  _GEN13776 = io_x[42] ? _GEN13775 : _GEN6863;
wire  _GEN13777 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13778 = io_x[0] ? _GEN6845 : _GEN13777;
wire  _GEN13779 = io_x[76] ? _GEN6834 : _GEN13778;
wire  _GEN13780 = io_x[42] ? _GEN13779 : _GEN6874;
wire  _GEN13781 = io_x[38] ? _GEN13780 : _GEN13776;
wire  _GEN13782 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN13783 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN13784 = io_x[76] ? _GEN6834 : _GEN13783;
wire  _GEN13785 = io_x[42] ? _GEN13784 : _GEN13782;
wire  _GEN13786 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN13787 = io_x[6] ? _GEN6850 : _GEN13786;
wire  _GEN13788 = io_x[41] ? _GEN13787 : _GEN6836;
wire  _GEN13789 = io_x[14] ? _GEN6856 : _GEN13788;
wire  _GEN13790 = io_x[0] ? _GEN13789 : _GEN6845;
wire  _GEN13791 = io_x[76] ? _GEN13790 : _GEN6833;
wire  _GEN13792 = io_x[42] ? _GEN13791 : _GEN6874;
wire  _GEN13793 = io_x[38] ? _GEN13792 : _GEN13785;
wire  _GEN13794 = io_x[10] ? _GEN13793 : _GEN13781;
wire  _GEN13795 = io_x[71] ? _GEN13794 : _GEN13769;
wire  _GEN13796 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN13797 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN13798 = io_x[42] ? _GEN13797 : _GEN13796;
wire  _GEN13799 = io_x[38] ? _GEN6871 : _GEN13798;
wire  _GEN13800 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN13801 = io_x[14] ? _GEN6843 : _GEN13800;
wire  _GEN13802 = io_x[0] ? _GEN13801 : _GEN6858;
wire  _GEN13803 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13804 = io_x[41] ? _GEN6836 : _GEN13803;
wire  _GEN13805 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13806 = io_x[41] ? _GEN6836 : _GEN13805;
wire  _GEN13807 = io_x[14] ? _GEN13806 : _GEN13804;
wire  _GEN13808 = io_x[0] ? _GEN13807 : _GEN6858;
wire  _GEN13809 = io_x[76] ? _GEN13808 : _GEN13802;
wire  _GEN13810 = io_x[42] ? _GEN13809 : _GEN6874;
wire  _GEN13811 = io_x[38] ? _GEN6871 : _GEN13810;
wire  _GEN13812 = io_x[10] ? _GEN13811 : _GEN13799;
wire  _GEN13813 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN13814 = io_x[10] ? _GEN13813 : _GEN7044;
wire  _GEN13815 = io_x[71] ? _GEN13814 : _GEN13812;
wire  _GEN13816 = io_x[70] ? _GEN13815 : _GEN13795;
wire  _GEN13817 = io_x[33] ? _GEN12627 : _GEN13816;
wire  _GEN13818 = io_x[21] ? _GEN13817 : _GEN13741;
wire  _GEN13819 = io_x[18] ? _GEN13818 : _GEN13685;
wire  _GEN13820 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN13821 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13822 = io_x[41] ? _GEN13821 : _GEN6836;
wire  _GEN13823 = io_x[14] ? _GEN13822 : _GEN13820;
wire  _GEN13824 = io_x[0] ? _GEN6845 : _GEN13823;
wire  _GEN13825 = io_x[76] ? _GEN6834 : _GEN13824;
wire  _GEN13826 = io_x[42] ? _GEN13825 : _GEN6874;
wire  _GEN13827 = io_x[38] ? _GEN6871 : _GEN13826;
wire  _GEN13828 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN13829 = io_x[10] ? _GEN13828 : _GEN13827;
wire  _GEN13830 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN13831 = io_x[6] ? _GEN6850 : _GEN13830;
wire  _GEN13832 = io_x[41] ? _GEN6836 : _GEN13831;
wire  _GEN13833 = io_x[14] ? _GEN6856 : _GEN13832;
wire  _GEN13834 = io_x[0] ? _GEN13833 : _GEN6845;
wire  _GEN13835 = io_x[76] ? _GEN6834 : _GEN13834;
wire  _GEN13836 = io_x[42] ? _GEN13835 : _GEN6874;
wire  _GEN13837 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13838 = io_x[41] ? _GEN13837 : _GEN6836;
wire  _GEN13839 = io_x[14] ? _GEN6843 : _GEN13838;
wire  _GEN13840 = io_x[0] ? _GEN6845 : _GEN13839;
wire  _GEN13841 = io_x[76] ? _GEN6834 : _GEN13840;
wire  _GEN13842 = io_x[42] ? _GEN13841 : _GEN6874;
wire  _GEN13843 = io_x[38] ? _GEN13842 : _GEN13836;
wire  _GEN13844 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN13845 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13846 = io_x[41] ? _GEN6924 : _GEN13845;
wire  _GEN13847 = io_x[14] ? _GEN13846 : _GEN13844;
wire  _GEN13848 = io_x[0] ? _GEN13847 : _GEN6845;
wire  _GEN13849 = io_x[76] ? _GEN6834 : _GEN13848;
wire  _GEN13850 = io_x[42] ? _GEN13849 : _GEN6874;
wire  _GEN13851 = io_x[38] ? _GEN7036 : _GEN13850;
wire  _GEN13852 = io_x[10] ? _GEN13851 : _GEN13843;
wire  _GEN13853 = io_x[71] ? _GEN13852 : _GEN13829;
wire  _GEN13854 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN13855 = io_x[10] ? _GEN13854 : _GEN7094;
wire  _GEN13856 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN13857 = io_x[71] ? _GEN13856 : _GEN13855;
wire  _GEN13858 = io_x[70] ? _GEN13857 : _GEN13853;
wire  _GEN13859 = io_x[33] ? _GEN12627 : _GEN13858;
wire  _GEN13860 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN13861 = io_x[14] ? _GEN13860 : _GEN6843;
wire  _GEN13862 = io_x[0] ? _GEN6845 : _GEN13861;
wire  _GEN13863 = io_x[76] ? _GEN6833 : _GEN13862;
wire  _GEN13864 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13865 = io_x[0] ? _GEN6858 : _GEN13864;
wire  _GEN13866 = io_x[76] ? _GEN6834 : _GEN13865;
wire  _GEN13867 = io_x[42] ? _GEN13866 : _GEN13863;
wire  _GEN13868 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13869 = io_x[0] ? _GEN13868 : _GEN6845;
wire  _GEN13870 = io_x[76] ? _GEN13869 : _GEN6834;
wire  _GEN13871 = io_x[42] ? _GEN6874 : _GEN13870;
wire  _GEN13872 = io_x[38] ? _GEN13871 : _GEN13867;
wire  _GEN13873 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN13874 = io_x[10] ? _GEN13873 : _GEN13872;
wire  _GEN13875 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13876 = io_x[0] ? _GEN13875 : _GEN6845;
wire  _GEN13877 = io_x[76] ? _GEN6834 : _GEN13876;
wire  _GEN13878 = io_x[42] ? _GEN6863 : _GEN13877;
wire  _GEN13879 = io_x[38] ? _GEN6871 : _GEN13878;
wire  _GEN13880 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN13881 = io_x[0] ? _GEN13880 : _GEN6845;
wire  _GEN13882 = io_x[76] ? _GEN13881 : _GEN6833;
wire  _GEN13883 = io_x[42] ? _GEN6874 : _GEN13882;
wire  _GEN13884 = io_x[38] ? _GEN7036 : _GEN13883;
wire  _GEN13885 = io_x[10] ? _GEN13884 : _GEN13879;
wire  _GEN13886 = io_x[71] ? _GEN13885 : _GEN13874;
wire  _GEN13887 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN13888 = io_x[14] ? _GEN6843 : _GEN13887;
wire  _GEN13889 = io_x[0] ? _GEN6845 : _GEN13888;
wire  _GEN13890 = io_x[76] ? _GEN13889 : _GEN6834;
wire  _GEN13891 = io_x[42] ? _GEN6874 : _GEN13890;
wire  _GEN13892 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN13893 = io_x[42] ? _GEN13892 : _GEN6874;
wire  _GEN13894 = io_x[38] ? _GEN13893 : _GEN13891;
wire  _GEN13895 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN13896 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN13897 = io_x[76] ? _GEN6833 : _GEN13896;
wire  _GEN13898 = io_x[42] ? _GEN13897 : _GEN13895;
wire  _GEN13899 = io_x[38] ? _GEN6871 : _GEN13898;
wire  _GEN13900 = io_x[10] ? _GEN13899 : _GEN13894;
wire  _GEN13901 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN13902 = io_x[76] ? _GEN6834 : _GEN13901;
wire  _GEN13903 = io_x[42] ? _GEN13902 : _GEN6874;
wire  _GEN13904 = io_x[38] ? _GEN6871 : _GEN13903;
wire  _GEN13905 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN13906 = io_x[38] ? _GEN13905 : _GEN6871;
wire  _GEN13907 = io_x[10] ? _GEN13906 : _GEN13904;
wire  _GEN13908 = io_x[71] ? _GEN13907 : _GEN13900;
wire  _GEN13909 = io_x[70] ? _GEN13908 : _GEN13886;
wire  _GEN13910 = io_x[33] ? _GEN12641 : _GEN13909;
wire  _GEN13911 = io_x[21] ? _GEN13910 : _GEN13859;
wire  _GEN13912 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN13913 = io_x[42] ? _GEN13912 : _GEN6874;
wire  _GEN13914 = io_x[38] ? _GEN6871 : _GEN13913;
wire  _GEN13915 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13916 = io_x[0] ? _GEN13915 : _GEN6845;
wire  _GEN13917 = io_x[76] ? _GEN6834 : _GEN13916;
wire  _GEN13918 = io_x[42] ? _GEN13917 : _GEN6874;
wire  _GEN13919 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN13920 = io_x[42] ? _GEN13919 : _GEN6863;
wire  _GEN13921 = io_x[38] ? _GEN13920 : _GEN13918;
wire  _GEN13922 = io_x[10] ? _GEN13921 : _GEN13914;
wire  _GEN13923 = io_x[71] ? _GEN7196 : _GEN13922;
wire  _GEN13924 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN13925 = io_x[6] ? _GEN6850 : _GEN13924;
wire  _GEN13926 = io_x[41] ? _GEN6836 : _GEN13925;
wire  _GEN13927 = io_x[14] ? _GEN6843 : _GEN13926;
wire  _GEN13928 = io_x[0] ? _GEN6858 : _GEN13927;
wire  _GEN13929 = io_x[76] ? _GEN13928 : _GEN6834;
wire  _GEN13930 = io_x[42] ? _GEN13929 : _GEN6863;
wire  _GEN13931 = io_x[38] ? _GEN13930 : _GEN6871;
wire  _GEN13932 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13933 = io_x[41] ? _GEN6836 : _GEN13932;
wire  _GEN13934 = io_x[14] ? _GEN13933 : _GEN6856;
wire  _GEN13935 = io_x[0] ? _GEN13934 : _GEN6845;
wire  _GEN13936 = io_x[76] ? _GEN13935 : _GEN6834;
wire  _GEN13937 = io_x[42] ? _GEN13936 : _GEN6874;
wire  _GEN13938 = io_x[38] ? _GEN13937 : _GEN6871;
wire  _GEN13939 = io_x[10] ? _GEN13938 : _GEN13931;
wire  _GEN13940 = io_x[71] ? _GEN13939 : _GEN7196;
wire  _GEN13941 = io_x[70] ? _GEN13940 : _GEN13923;
wire  _GEN13942 = io_x[33] ? _GEN12641 : _GEN13941;
wire  _GEN13943 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13944 = io_x[41] ? _GEN13943 : _GEN6836;
wire  _GEN13945 = io_x[14] ? _GEN13944 : _GEN6843;
wire  _GEN13946 = io_x[0] ? _GEN13945 : _GEN6845;
wire  _GEN13947 = io_x[76] ? _GEN13946 : _GEN6834;
wire  _GEN13948 = io_x[42] ? _GEN6874 : _GEN13947;
wire  _GEN13949 = io_x[38] ? _GEN13948 : _GEN7036;
wire  _GEN13950 = io_x[10] ? _GEN7044 : _GEN13949;
wire  _GEN13951 = io_x[71] ? _GEN7196 : _GEN13950;
wire  _GEN13952 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN13953 = io_x[0] ? _GEN6845 : _GEN13952;
wire  _GEN13954 = io_x[76] ? _GEN13953 : _GEN6834;
wire  _GEN13955 = io_x[42] ? _GEN6874 : _GEN13954;
wire  _GEN13956 = io_x[38] ? _GEN6871 : _GEN13955;
wire  _GEN13957 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13958 = io_x[41] ? _GEN6836 : _GEN13957;
wire  _GEN13959 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN13960 = io_x[41] ? _GEN6836 : _GEN13959;
wire  _GEN13961 = io_x[14] ? _GEN13960 : _GEN13958;
wire  _GEN13962 = io_x[0] ? _GEN13961 : _GEN6845;
wire  _GEN13963 = io_x[76] ? _GEN13962 : _GEN6834;
wire  _GEN13964 = io_x[42] ? _GEN13963 : _GEN6874;
wire  _GEN13965 = io_x[38] ? _GEN7036 : _GEN13964;
wire  _GEN13966 = io_x[10] ? _GEN13965 : _GEN13956;
wire  _GEN13967 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN13968 = io_x[42] ? _GEN13967 : _GEN6874;
wire  _GEN13969 = io_x[38] ? _GEN7036 : _GEN13968;
wire  _GEN13970 = io_x[10] ? _GEN13969 : _GEN7044;
wire  _GEN13971 = io_x[71] ? _GEN13970 : _GEN13966;
wire  _GEN13972 = io_x[70] ? _GEN13971 : _GEN13951;
wire  _GEN13973 = io_x[33] ? _GEN12627 : _GEN13972;
wire  _GEN13974 = io_x[21] ? _GEN13973 : _GEN13942;
wire  _GEN13975 = io_x[18] ? _GEN13974 : _GEN13911;
wire  _GEN13976 = io_x[20] ? _GEN13975 : _GEN13819;
wire  _GEN13977 = io_x[71] ? _GEN7203 : _GEN7196;
wire  _GEN13978 = io_x[70] ? _GEN13977 : _GEN8474;
wire  _GEN13979 = io_x[33] ? _GEN12627 : _GEN13978;
wire  _GEN13980 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN13981 = io_x[10] ? _GEN7044 : _GEN13980;
wire  _GEN13982 = io_x[71] ? _GEN13981 : _GEN7196;
wire  _GEN13983 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN13984 = io_x[14] ? _GEN6843 : _GEN13983;
wire  _GEN13985 = io_x[0] ? _GEN6845 : _GEN13984;
wire  _GEN13986 = io_x[76] ? _GEN6834 : _GEN13985;
wire  _GEN13987 = io_x[42] ? _GEN6874 : _GEN13986;
wire  _GEN13988 = io_x[38] ? _GEN13987 : _GEN6871;
wire  _GEN13989 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN13990 = io_x[10] ? _GEN13989 : _GEN13988;
wire  _GEN13991 = io_x[71] ? _GEN7196 : _GEN13990;
wire  _GEN13992 = io_x[70] ? _GEN13991 : _GEN13982;
wire  _GEN13993 = io_x[33] ? _GEN12627 : _GEN13992;
wire  _GEN13994 = io_x[21] ? _GEN13993 : _GEN13979;
wire  _GEN13995 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN13996 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN13997 = io_x[41] ? _GEN6836 : _GEN13996;
wire  _GEN13998 = io_x[14] ? _GEN13997 : _GEN6843;
wire  _GEN13999 = io_x[0] ? _GEN13998 : _GEN6845;
wire  _GEN14000 = io_x[76] ? _GEN6834 : _GEN13999;
wire  _GEN14001 = io_x[42] ? _GEN6874 : _GEN14000;
wire  _GEN14002 = io_x[38] ? _GEN6871 : _GEN14001;
wire  _GEN14003 = io_x[10] ? _GEN14002 : _GEN13995;
wire  _GEN14004 = io_x[71] ? _GEN7196 : _GEN14003;
wire  _GEN14005 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN14006 = io_x[10] ? _GEN14005 : _GEN7044;
wire  _GEN14007 = io_x[71] ? _GEN7196 : _GEN14006;
wire  _GEN14008 = io_x[70] ? _GEN14007 : _GEN14004;
wire  _GEN14009 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14010 = io_x[41] ? _GEN6836 : _GEN14009;
wire  _GEN14011 = io_x[14] ? _GEN14010 : _GEN6843;
wire  _GEN14012 = io_x[0] ? _GEN14011 : _GEN6845;
wire  _GEN14013 = io_x[76] ? _GEN6834 : _GEN14012;
wire  _GEN14014 = io_x[42] ? _GEN6874 : _GEN14013;
wire  _GEN14015 = io_x[38] ? _GEN6871 : _GEN14014;
wire  _GEN14016 = io_x[10] ? _GEN14015 : _GEN7044;
wire  _GEN14017 = io_x[71] ? _GEN7196 : _GEN14016;
wire  _GEN14018 = io_x[70] ? _GEN8474 : _GEN14017;
wire  _GEN14019 = io_x[33] ? _GEN14018 : _GEN14008;
wire  _GEN14020 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14021 = io_x[41] ? _GEN14020 : _GEN6836;
wire  _GEN14022 = io_x[14] ? _GEN14021 : _GEN6843;
wire  _GEN14023 = io_x[0] ? _GEN6845 : _GEN14022;
wire  _GEN14024 = io_x[76] ? _GEN14023 : _GEN6834;
wire  _GEN14025 = io_x[42] ? _GEN6874 : _GEN14024;
wire  _GEN14026 = io_x[38] ? _GEN14025 : _GEN6871;
wire  _GEN14027 = io_x[10] ? _GEN14026 : _GEN7044;
wire  _GEN14028 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN14029 = io_x[0] ? _GEN6845 : _GEN14028;
wire  _GEN14030 = io_x[76] ? _GEN14029 : _GEN6834;
wire  _GEN14031 = io_x[42] ? _GEN6874 : _GEN14030;
wire  _GEN14032 = io_x[38] ? _GEN6871 : _GEN14031;
wire  _GEN14033 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN14034 = io_x[38] ? _GEN14033 : _GEN6871;
wire  _GEN14035 = io_x[10] ? _GEN14034 : _GEN14032;
wire  _GEN14036 = io_x[71] ? _GEN14035 : _GEN14027;
wire  _GEN14037 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN14038 = io_x[38] ? _GEN6871 : _GEN14037;
wire  _GEN14039 = io_x[10] ? _GEN14038 : _GEN7094;
wire  _GEN14040 = io_x[71] ? _GEN14039 : _GEN7196;
wire  _GEN14041 = io_x[70] ? _GEN14040 : _GEN14036;
wire  _GEN14042 = io_x[33] ? _GEN12627 : _GEN14041;
wire  _GEN14043 = io_x[21] ? _GEN14042 : _GEN14019;
wire  _GEN14044 = io_x[18] ? _GEN14043 : _GEN13994;
wire  _GEN14045 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN14046 = io_x[0] ? _GEN14045 : _GEN6845;
wire  _GEN14047 = io_x[76] ? _GEN14046 : _GEN6834;
wire  _GEN14048 = io_x[42] ? _GEN6874 : _GEN14047;
wire  _GEN14049 = io_x[38] ? _GEN6871 : _GEN14048;
wire  _GEN14050 = io_x[10] ? _GEN14049 : _GEN7044;
wire  _GEN14051 = io_x[71] ? _GEN7196 : _GEN14050;
wire  _GEN14052 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN14053 = io_x[0] ? _GEN14052 : _GEN6845;
wire  _GEN14054 = io_x[76] ? _GEN14053 : _GEN6834;
wire  _GEN14055 = io_x[42] ? _GEN14054 : _GEN6874;
wire  _GEN14056 = io_x[38] ? _GEN6871 : _GEN14055;
wire  _GEN14057 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN14058 = io_x[0] ? _GEN14057 : _GEN6845;
wire  _GEN14059 = io_x[76] ? _GEN14058 : _GEN6834;
wire  _GEN14060 = io_x[42] ? _GEN14059 : _GEN6863;
wire  _GEN14061 = io_x[38] ? _GEN6871 : _GEN14060;
wire  _GEN14062 = io_x[10] ? _GEN14061 : _GEN14056;
wire  _GEN14063 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14064 = io_x[41] ? _GEN14063 : _GEN6836;
wire  _GEN14065 = io_x[14] ? _GEN14064 : _GEN6843;
wire  _GEN14066 = io_x[0] ? _GEN6845 : _GEN14065;
wire  _GEN14067 = io_x[76] ? _GEN14066 : _GEN6834;
wire  _GEN14068 = io_x[42] ? _GEN6863 : _GEN14067;
wire  _GEN14069 = io_x[38] ? _GEN6871 : _GEN14068;
wire  _GEN14070 = io_x[10] ? _GEN14069 : _GEN7094;
wire  _GEN14071 = io_x[71] ? _GEN14070 : _GEN14062;
wire  _GEN14072 = io_x[70] ? _GEN14071 : _GEN14051;
wire  _GEN14073 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14074 = io_x[41] ? _GEN14073 : _GEN6836;
wire  _GEN14075 = io_x[14] ? _GEN14074 : _GEN6843;
wire  _GEN14076 = io_x[0] ? _GEN6845 : _GEN14075;
wire  _GEN14077 = io_x[76] ? _GEN14076 : _GEN6834;
wire  _GEN14078 = io_x[42] ? _GEN6874 : _GEN14077;
wire  _GEN14079 = io_x[38] ? _GEN6871 : _GEN14078;
wire  _GEN14080 = io_x[10] ? _GEN14079 : _GEN7044;
wire  _GEN14081 = io_x[71] ? _GEN7196 : _GEN14080;
wire  _GEN14082 = io_x[70] ? _GEN8474 : _GEN14081;
wire  _GEN14083 = io_x[33] ? _GEN14082 : _GEN14072;
wire  _GEN14084 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN14085 = io_x[0] ? _GEN14084 : _GEN6845;
wire  _GEN14086 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14087 = io_x[6] ? _GEN14086 : _GEN6850;
wire  _GEN14088 = io_x[41] ? _GEN14087 : _GEN6836;
wire  _GEN14089 = io_x[14] ? _GEN14088 : _GEN6843;
wire  _GEN14090 = io_x[0] ? _GEN14089 : _GEN6845;
wire  _GEN14091 = io_x[76] ? _GEN14090 : _GEN14085;
wire  _GEN14092 = io_x[42] ? _GEN6874 : _GEN14091;
wire  _GEN14093 = io_x[38] ? _GEN14092 : _GEN6871;
wire  _GEN14094 = io_x[10] ? _GEN14093 : _GEN7044;
wire  _GEN14095 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN14096 = io_x[71] ? _GEN14095 : _GEN14094;
wire  _GEN14097 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14098 = io_x[6] ? _GEN14097 : _GEN6850;
wire  _GEN14099 = io_x[41] ? _GEN14098 : _GEN6836;
wire  _GEN14100 = io_x[14] ? _GEN14099 : _GEN6843;
wire  _GEN14101 = io_x[0] ? _GEN6845 : _GEN14100;
wire  _GEN14102 = io_x[76] ? _GEN14101 : _GEN6834;
wire  _GEN14103 = io_x[42] ? _GEN6863 : _GEN14102;
wire  _GEN14104 = io_x[38] ? _GEN7036 : _GEN14103;
wire  _GEN14105 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN14106 = io_x[76] ? _GEN14105 : _GEN6833;
wire  _GEN14107 = io_x[42] ? _GEN6874 : _GEN14106;
wire  _GEN14108 = io_x[38] ? _GEN7036 : _GEN14107;
wire  _GEN14109 = io_x[10] ? _GEN14108 : _GEN14104;
wire  _GEN14110 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN14111 = io_x[0] ? _GEN14110 : _GEN6845;
wire  _GEN14112 = io_x[76] ? _GEN6833 : _GEN14111;
wire  _GEN14113 = io_x[42] ? _GEN6874 : _GEN14112;
wire  _GEN14114 = io_x[38] ? _GEN14113 : _GEN6871;
wire  _GEN14115 = io_x[10] ? _GEN14114 : _GEN7044;
wire  _GEN14116 = io_x[71] ? _GEN14115 : _GEN14109;
wire  _GEN14117 = io_x[70] ? _GEN14116 : _GEN14096;
wire  _GEN14118 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14119 = io_x[41] ? _GEN6836 : _GEN14118;
wire  _GEN14120 = io_x[14] ? _GEN14119 : _GEN6843;
wire  _GEN14121 = io_x[0] ? _GEN6845 : _GEN14120;
wire  _GEN14122 = io_x[76] ? _GEN6834 : _GEN14121;
wire  _GEN14123 = io_x[42] ? _GEN6874 : _GEN14122;
wire  _GEN14124 = io_x[38] ? _GEN6871 : _GEN14123;
wire  _GEN14125 = io_x[10] ? _GEN14124 : _GEN7044;
wire  _GEN14126 = io_x[71] ? _GEN7196 : _GEN14125;
wire  _GEN14127 = io_x[70] ? _GEN7020 : _GEN14126;
wire  _GEN14128 = io_x[33] ? _GEN14127 : _GEN14117;
wire  _GEN14129 = io_x[21] ? _GEN14128 : _GEN14083;
wire  _GEN14130 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN14131 = io_x[10] ? _GEN14130 : _GEN7044;
wire  _GEN14132 = io_x[71] ? _GEN7196 : _GEN14131;
wire  _GEN14133 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN14134 = io_x[71] ? _GEN14133 : _GEN7196;
wire  _GEN14135 = io_x[70] ? _GEN14134 : _GEN14132;
wire  _GEN14136 = io_x[33] ? _GEN12627 : _GEN14135;
wire  _GEN14137 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN14138 = io_x[76] ? _GEN14137 : _GEN6834;
wire  _GEN14139 = io_x[42] ? _GEN6874 : _GEN14138;
wire  _GEN14140 = io_x[38] ? _GEN14139 : _GEN6871;
wire  _GEN14141 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14142 = io_x[6] ? _GEN14141 : _GEN6850;
wire  _GEN14143 = io_x[41] ? _GEN14142 : _GEN6924;
wire  _GEN14144 = io_x[14] ? _GEN6843 : _GEN14143;
wire  _GEN14145 = io_x[0] ? _GEN14144 : _GEN6845;
wire  _GEN14146 = io_x[76] ? _GEN14145 : _GEN6834;
wire  _GEN14147 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14148 = io_x[6] ? _GEN14147 : _GEN6850;
wire  _GEN14149 = io_x[41] ? _GEN14148 : _GEN6836;
wire  _GEN14150 = io_x[14] ? _GEN14149 : _GEN6843;
wire  _GEN14151 = io_x[0] ? _GEN14150 : _GEN6845;
wire  _GEN14152 = io_x[76] ? _GEN14151 : _GEN6834;
wire  _GEN14153 = io_x[42] ? _GEN14152 : _GEN14146;
wire  _GEN14154 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN14155 = io_x[0] ? _GEN14154 : _GEN6845;
wire  _GEN14156 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14157 = io_x[41] ? _GEN14156 : _GEN6836;
wire  _GEN14158 = io_x[14] ? _GEN14157 : _GEN6843;
wire  _GEN14159 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14160 = io_x[6] ? _GEN14159 : _GEN6840;
wire  _GEN14161 = io_x[41] ? _GEN14160 : _GEN6836;
wire  _GEN14162 = io_x[14] ? _GEN14161 : _GEN6856;
wire  _GEN14163 = io_x[0] ? _GEN14162 : _GEN14158;
wire  _GEN14164 = io_x[76] ? _GEN14163 : _GEN14155;
wire  _GEN14165 = io_x[42] ? _GEN6874 : _GEN14164;
wire  _GEN14166 = io_x[38] ? _GEN14165 : _GEN14153;
wire  _GEN14167 = io_x[10] ? _GEN14166 : _GEN14140;
wire  _GEN14168 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN14169 = io_x[76] ? _GEN14168 : _GEN6834;
wire  _GEN14170 = io_x[42] ? _GEN6874 : _GEN14169;
wire  _GEN14171 = io_x[38] ? _GEN6871 : _GEN14170;
wire  _GEN14172 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN14173 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14174 = io_x[41] ? _GEN14173 : _GEN6836;
wire  _GEN14175 = io_x[14] ? _GEN14174 : _GEN6856;
wire  _GEN14176 = io_x[0] ? _GEN14175 : _GEN14172;
wire  _GEN14177 = io_x[76] ? _GEN14176 : _GEN6833;
wire  _GEN14178 = io_x[42] ? _GEN6874 : _GEN14177;
wire  _GEN14179 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN14180 = io_x[14] ? _GEN6843 : _GEN14179;
wire  _GEN14181 = io_x[0] ? _GEN14180 : _GEN6858;
wire  _GEN14182 = io_x[76] ? _GEN6833 : _GEN14181;
wire  _GEN14183 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14184 = io_x[41] ? _GEN6836 : _GEN14183;
wire  _GEN14185 = io_x[14] ? _GEN14184 : _GEN6843;
wire  _GEN14186 = io_x[0] ? _GEN14185 : _GEN6845;
wire  _GEN14187 = io_x[76] ? _GEN14186 : _GEN6834;
wire  _GEN14188 = io_x[42] ? _GEN14187 : _GEN14182;
wire  _GEN14189 = io_x[38] ? _GEN14188 : _GEN14178;
wire  _GEN14190 = io_x[10] ? _GEN14189 : _GEN14171;
wire  _GEN14191 = io_x[71] ? _GEN14190 : _GEN14167;
wire  _GEN14192 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14193 = io_x[41] ? _GEN14192 : _GEN6836;
wire  _GEN14194 = io_x[14] ? _GEN14193 : _GEN6843;
wire  _GEN14195 = io_x[0] ? _GEN14194 : _GEN6858;
wire  _GEN14196 = io_x[76] ? _GEN14195 : _GEN6834;
wire  _GEN14197 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN14198 = io_x[76] ? _GEN14197 : _GEN6834;
wire  _GEN14199 = io_x[42] ? _GEN14198 : _GEN14196;
wire  _GEN14200 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN14201 = io_x[42] ? _GEN6863 : _GEN14200;
wire  _GEN14202 = io_x[38] ? _GEN14201 : _GEN14199;
wire  _GEN14203 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN14204 = io_x[0] ? _GEN14203 : _GEN6845;
wire  _GEN14205 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14206 = io_x[6] ? _GEN14205 : _GEN6840;
wire  _GEN14207 = io_x[41] ? _GEN14206 : _GEN6836;
wire  _GEN14208 = io_x[14] ? _GEN14207 : _GEN6856;
wire  _GEN14209 = io_x[0] ? _GEN14208 : _GEN6858;
wire  _GEN14210 = io_x[76] ? _GEN14209 : _GEN14204;
wire  _GEN14211 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN14212 = io_x[76] ? _GEN14211 : _GEN6834;
wire  _GEN14213 = io_x[42] ? _GEN14212 : _GEN14210;
wire  _GEN14214 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN14215 = io_x[0] ? _GEN14214 : _GEN6845;
wire  _GEN14216 = io_x[76] ? _GEN14215 : _GEN6833;
wire  _GEN14217 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN14218 = io_x[76] ? _GEN14217 : _GEN6834;
wire  _GEN14219 = io_x[42] ? _GEN14218 : _GEN14216;
wire  _GEN14220 = io_x[38] ? _GEN14219 : _GEN14213;
wire  _GEN14221 = io_x[10] ? _GEN14220 : _GEN14202;
wire  _GEN14222 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14223 = io_x[41] ? _GEN14222 : _GEN6836;
wire  _GEN14224 = io_x[14] ? _GEN14223 : _GEN6856;
wire  _GEN14225 = io_x[0] ? _GEN14224 : _GEN6845;
wire  _GEN14226 = io_x[76] ? _GEN14225 : _GEN6834;
wire  _GEN14227 = io_x[42] ? _GEN6874 : _GEN14226;
wire  _GEN14228 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN14229 = io_x[0] ? _GEN14228 : _GEN6845;
wire  _GEN14230 = io_x[76] ? _GEN6834 : _GEN14229;
wire  _GEN14231 = io_x[42] ? _GEN6863 : _GEN14230;
wire  _GEN14232 = io_x[38] ? _GEN14231 : _GEN14227;
wire  _GEN14233 = io_x[10] ? _GEN14232 : _GEN7044;
wire  _GEN14234 = io_x[71] ? _GEN14233 : _GEN14221;
wire  _GEN14235 = io_x[70] ? _GEN14234 : _GEN14191;
wire  _GEN14236 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14237 = io_x[41] ? _GEN14236 : _GEN6836;
wire  _GEN14238 = io_x[14] ? _GEN14237 : _GEN6843;
wire  _GEN14239 = io_x[0] ? _GEN14238 : _GEN6845;
wire  _GEN14240 = io_x[76] ? _GEN14239 : _GEN6833;
wire  _GEN14241 = io_x[42] ? _GEN6874 : _GEN14240;
wire  _GEN14242 = io_x[38] ? _GEN6871 : _GEN14241;
wire  _GEN14243 = io_x[10] ? _GEN14242 : _GEN7044;
wire  _GEN14244 = io_x[71] ? _GEN7196 : _GEN14243;
wire  _GEN14245 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14246 = io_x[6] ? _GEN14245 : _GEN6850;
wire  _GEN14247 = io_x[41] ? _GEN14246 : _GEN6836;
wire  _GEN14248 = io_x[14] ? _GEN14247 : _GEN6843;
wire  _GEN14249 = io_x[0] ? _GEN14248 : _GEN6845;
wire  _GEN14250 = io_x[76] ? _GEN14249 : _GEN6834;
wire  _GEN14251 = io_x[42] ? _GEN6874 : _GEN14250;
wire  _GEN14252 = io_x[38] ? _GEN6871 : _GEN14251;
wire  _GEN14253 = io_x[10] ? _GEN14252 : _GEN7044;
wire  _GEN14254 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN14255 = io_x[71] ? _GEN14254 : _GEN14253;
wire  _GEN14256 = io_x[70] ? _GEN14255 : _GEN14244;
wire  _GEN14257 = io_x[33] ? _GEN14256 : _GEN14235;
wire  _GEN14258 = io_x[21] ? _GEN14257 : _GEN14136;
wire  _GEN14259 = io_x[18] ? _GEN14258 : _GEN14129;
wire  _GEN14260 = io_x[20] ? _GEN14259 : _GEN14044;
wire  _GEN14261 = io_x[45] ? _GEN14260 : _GEN13976;
wire  _GEN14262 = io_x[28] ? _GEN14261 : _GEN13613;
wire  _GEN14263 = 1'b1;
wire  _GEN14264 = 1'b1;
wire  _GEN14265 = io_x[18] ? _GEN12920 : _GEN14264;
wire  _GEN14266 = io_x[71] ? _GEN7196 : _GEN7203;
wire  _GEN14267 = io_x[70] ? _GEN7020 : _GEN14266;
wire  _GEN14268 = io_x[33] ? _GEN12627 : _GEN14267;
wire  _GEN14269 = io_x[21] ? _GEN14268 : _GEN12933;
wire  _GEN14270 = io_x[18] ? _GEN14269 : _GEN14264;
wire  _GEN14271 = io_x[20] ? _GEN14270 : _GEN14265;
wire  _GEN14272 = io_x[45] ? _GEN14271 : _GEN14263;
wire  _GEN14273 = 1'b1;
wire  _GEN14274 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN14275 = io_x[0] ? _GEN14274 : _GEN6845;
wire  _GEN14276 = io_x[76] ? _GEN6834 : _GEN14275;
wire  _GEN14277 = io_x[42] ? _GEN14276 : _GEN6874;
wire  _GEN14278 = io_x[38] ? _GEN6871 : _GEN14277;
wire  _GEN14279 = io_x[10] ? _GEN14278 : _GEN7094;
wire  _GEN14280 = io_x[71] ? _GEN7196 : _GEN14279;
wire  _GEN14281 = io_x[70] ? _GEN8474 : _GEN14280;
wire  _GEN14282 = io_x[33] ? _GEN12627 : _GEN14281;
wire  _GEN14283 = io_x[21] ? _GEN14282 : _GEN12643;
wire  _GEN14284 = io_x[18] ? _GEN14283 : _GEN14264;
wire  _GEN14285 = io_x[20] ? _GEN14284 : _GEN14273;
wire  _GEN14286 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN14287 = io_x[42] ? _GEN6874 : _GEN14286;
wire  _GEN14288 = io_x[38] ? _GEN6871 : _GEN14287;
wire  _GEN14289 = io_x[10] ? _GEN14288 : _GEN7044;
wire  _GEN14290 = io_x[71] ? _GEN14289 : _GEN7196;
wire  _GEN14291 = io_x[70] ? _GEN14290 : _GEN8474;
wire  _GEN14292 = io_x[33] ? _GEN12627 : _GEN14291;
wire  _GEN14293 = io_x[21] ? _GEN12643 : _GEN14292;
wire  _GEN14294 = io_x[18] ? _GEN14264 : _GEN14293;
wire  _GEN14295 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN14296 = io_x[71] ? _GEN7196 : _GEN14295;
wire  _GEN14297 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN14298 = io_x[71] ? _GEN7203 : _GEN14297;
wire  _GEN14299 = io_x[70] ? _GEN14298 : _GEN14296;
wire  _GEN14300 = io_x[33] ? _GEN12627 : _GEN14299;
wire  _GEN14301 = io_x[70] ? _GEN8474 : _GEN7020;
wire  _GEN14302 = io_x[33] ? _GEN12627 : _GEN14301;
wire  _GEN14303 = io_x[21] ? _GEN14302 : _GEN14300;
wire  _GEN14304 = io_x[18] ? _GEN14303 : _GEN14264;
wire  _GEN14305 = io_x[20] ? _GEN14304 : _GEN14294;
wire  _GEN14306 = io_x[45] ? _GEN14305 : _GEN14285;
wire  _GEN14307 = io_x[28] ? _GEN14306 : _GEN14272;
wire  _GEN14308 = io_x[79] ? _GEN14307 : _GEN14262;
wire  _GEN14309 = io_x[48] ? _GEN14308 : _GEN12982;
wire  _GEN14310 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN14311 = io_x[38] ? _GEN6871 : _GEN14310;
wire  _GEN14312 = io_x[10] ? _GEN7044 : _GEN14311;
wire  _GEN14313 = io_x[71] ? _GEN7203 : _GEN14312;
wire  _GEN14314 = io_x[70] ? _GEN14313 : _GEN7020;
wire  _GEN14315 = io_x[33] ? _GEN12627 : _GEN14314;
wire  _GEN14316 = io_x[21] ? _GEN12933 : _GEN14315;
wire  _GEN14317 = io_x[18] ? _GEN12920 : _GEN14316;
wire  _GEN14318 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN14319 = io_x[0] ? _GEN6845 : _GEN14318;
wire  _GEN14320 = io_x[76] ? _GEN6833 : _GEN14319;
wire  _GEN14321 = io_x[42] ? _GEN6874 : _GEN14320;
wire  _GEN14322 = io_x[38] ? _GEN14321 : _GEN7036;
wire  _GEN14323 = io_x[10] ? _GEN7044 : _GEN14322;
wire  _GEN14324 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN14325 = io_x[10] ? _GEN7044 : _GEN14324;
wire  _GEN14326 = io_x[71] ? _GEN14325 : _GEN14323;
wire  _GEN14327 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN14328 = io_x[38] ? _GEN6871 : _GEN14327;
wire  _GEN14329 = io_x[10] ? _GEN7044 : _GEN14328;
wire  _GEN14330 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN14331 = io_x[38] ? _GEN14330 : _GEN6871;
wire  _GEN14332 = io_x[10] ? _GEN7044 : _GEN14331;
wire  _GEN14333 = io_x[71] ? _GEN14332 : _GEN14329;
wire  _GEN14334 = io_x[70] ? _GEN14333 : _GEN14326;
wire  _GEN14335 = io_x[33] ? _GEN12627 : _GEN14334;
wire  _GEN14336 = io_x[21] ? _GEN14335 : _GEN12933;
wire  _GEN14337 = io_x[18] ? _GEN14336 : _GEN12920;
wire  _GEN14338 = io_x[20] ? _GEN14337 : _GEN14317;
wire  _GEN14339 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN14340 = io_x[10] ? _GEN7044 : _GEN14339;
wire  _GEN14341 = io_x[71] ? _GEN14340 : _GEN7203;
wire  _GEN14342 = io_x[70] ? _GEN14341 : _GEN8474;
wire  _GEN14343 = io_x[33] ? _GEN12627 : _GEN14342;
wire  _GEN14344 = io_x[21] ? _GEN12933 : _GEN14343;
wire  _GEN14345 = io_x[18] ? _GEN14344 : _GEN12920;
wire  _GEN14346 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN14347 = io_x[71] ? _GEN14346 : _GEN7196;
wire  _GEN14348 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN14349 = io_x[2] ? _GEN6837 : _GEN14348;
wire  _GEN14350 = io_x[6] ? _GEN6850 : _GEN14349;
wire  _GEN14351 = io_x[41] ? _GEN14350 : _GEN6836;
wire  _GEN14352 = io_x[14] ? _GEN6843 : _GEN14351;
wire  _GEN14353 = io_x[0] ? _GEN6845 : _GEN14352;
wire  _GEN14354 = io_x[76] ? _GEN6834 : _GEN14353;
wire  _GEN14355 = io_x[42] ? _GEN14354 : _GEN6874;
wire  _GEN14356 = io_x[38] ? _GEN6871 : _GEN14355;
wire  _GEN14357 = io_x[10] ? _GEN7044 : _GEN14356;
wire  _GEN14358 = io_x[71] ? _GEN14357 : _GEN7203;
wire  _GEN14359 = io_x[70] ? _GEN14358 : _GEN14347;
wire  _GEN14360 = io_x[33] ? _GEN12627 : _GEN14359;
wire  _GEN14361 = io_x[21] ? _GEN14360 : _GEN12933;
wire  _GEN14362 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14363 = io_x[6] ? _GEN6840 : _GEN14362;
wire  _GEN14364 = io_x[41] ? _GEN14363 : _GEN6836;
wire  _GEN14365 = io_x[14] ? _GEN6843 : _GEN14364;
wire  _GEN14366 = io_x[0] ? _GEN6845 : _GEN14365;
wire  _GEN14367 = io_x[76] ? _GEN14366 : _GEN6834;
wire  _GEN14368 = io_x[42] ? _GEN6874 : _GEN14367;
wire  _GEN14369 = io_x[38] ? _GEN14368 : _GEN6871;
wire  _GEN14370 = io_x[10] ? _GEN7044 : _GEN14369;
wire  _GEN14371 = io_x[71] ? _GEN7203 : _GEN14370;
wire  _GEN14372 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14373 = io_x[6] ? _GEN6840 : _GEN14372;
wire  _GEN14374 = io_x[41] ? _GEN14373 : _GEN6836;
wire  _GEN14375 = io_x[14] ? _GEN6843 : _GEN14374;
wire  _GEN14376 = io_x[0] ? _GEN6845 : _GEN14375;
wire  _GEN14377 = io_x[76] ? _GEN14376 : _GEN6834;
wire  _GEN14378 = io_x[42] ? _GEN6874 : _GEN14377;
wire  _GEN14379 = io_x[38] ? _GEN14378 : _GEN6871;
wire  _GEN14380 = io_x[10] ? _GEN7044 : _GEN14379;
wire  _GEN14381 = io_x[71] ? _GEN14380 : _GEN7196;
wire  _GEN14382 = io_x[70] ? _GEN14381 : _GEN14371;
wire  _GEN14383 = io_x[33] ? _GEN12627 : _GEN14382;
wire  _GEN14384 = io_x[21] ? _GEN14383 : _GEN12643;
wire  _GEN14385 = io_x[18] ? _GEN14384 : _GEN14361;
wire  _GEN14386 = io_x[20] ? _GEN14385 : _GEN14345;
wire  _GEN14387 = io_x[45] ? _GEN14386 : _GEN14338;
wire  _GEN14388 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN14389 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN14390 = io_x[0] ? _GEN6845 : _GEN14389;
wire  _GEN14391 = io_x[76] ? _GEN6834 : _GEN14390;
wire  _GEN14392 = io_x[42] ? _GEN6874 : _GEN14391;
wire  _GEN14393 = io_x[38] ? _GEN14392 : _GEN6871;
wire  _GEN14394 = io_x[10] ? _GEN7094 : _GEN14393;
wire  _GEN14395 = io_x[71] ? _GEN14394 : _GEN14388;
wire  _GEN14396 = io_x[70] ? _GEN14395 : _GEN7020;
wire  _GEN14397 = io_x[33] ? _GEN12627 : _GEN14396;
wire  _GEN14398 = io_x[21] ? _GEN14397 : _GEN12933;
wire  _GEN14399 = io_x[18] ? _GEN14398 : _GEN12920;
wire  _GEN14400 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN14401 = io_x[0] ? _GEN6845 : _GEN14400;
wire  _GEN14402 = io_x[76] ? _GEN6833 : _GEN14401;
wire  _GEN14403 = io_x[42] ? _GEN6874 : _GEN14402;
wire  _GEN14404 = io_x[38] ? _GEN14403 : _GEN6871;
wire  _GEN14405 = io_x[10] ? _GEN14404 : _GEN7094;
wire  _GEN14406 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN14407 = io_x[0] ? _GEN6845 : _GEN14406;
wire  _GEN14408 = io_x[76] ? _GEN14407 : _GEN6833;
wire  _GEN14409 = io_x[42] ? _GEN6874 : _GEN14408;
wire  _GEN14410 = io_x[38] ? _GEN14409 : _GEN6871;
wire  _GEN14411 = io_x[10] ? _GEN14410 : _GEN7094;
wire  _GEN14412 = io_x[71] ? _GEN14411 : _GEN14405;
wire  _GEN14413 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN14414 = io_x[38] ? _GEN7036 : _GEN14413;
wire  _GEN14415 = io_x[10] ? _GEN7094 : _GEN14414;
wire  _GEN14416 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN14417 = io_x[14] ? _GEN6843 : _GEN14416;
wire  _GEN14418 = io_x[0] ? _GEN6845 : _GEN14417;
wire  _GEN14419 = io_x[76] ? _GEN14418 : _GEN6833;
wire  _GEN14420 = io_x[42] ? _GEN6874 : _GEN14419;
wire  _GEN14421 = io_x[38] ? _GEN14420 : _GEN7036;
wire  _GEN14422 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN14423 = io_x[10] ? _GEN14422 : _GEN14421;
wire  _GEN14424 = io_x[71] ? _GEN14423 : _GEN14415;
wire  _GEN14425 = io_x[70] ? _GEN14424 : _GEN14412;
wire  _GEN14426 = io_x[33] ? _GEN12627 : _GEN14425;
wire  _GEN14427 = io_x[21] ? _GEN14426 : _GEN12933;
wire  _GEN14428 = io_x[18] ? _GEN14427 : _GEN12920;
wire  _GEN14429 = io_x[20] ? _GEN14428 : _GEN14399;
wire  _GEN14430 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN14431 = io_x[71] ? _GEN14430 : _GEN7196;
wire  _GEN14432 = io_x[70] ? _GEN7020 : _GEN14431;
wire  _GEN14433 = io_x[33] ? _GEN12627 : _GEN14432;
wire  _GEN14434 = io_x[21] ? _GEN14433 : _GEN12933;
wire  _GEN14435 = io_x[18] ? _GEN14434 : _GEN12920;
wire  _GEN14436 = io_x[71] ? _GEN7196 : _GEN7203;
wire  _GEN14437 = io_x[70] ? _GEN7020 : _GEN14436;
wire  _GEN14438 = io_x[33] ? _GEN12627 : _GEN14437;
wire  _GEN14439 = io_x[21] ? _GEN14438 : _GEN12643;
wire  _GEN14440 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14441 = io_x[41] ? _GEN14440 : _GEN6836;
wire  _GEN14442 = io_x[14] ? _GEN14441 : _GEN6843;
wire  _GEN14443 = io_x[0] ? _GEN6845 : _GEN14442;
wire  _GEN14444 = io_x[76] ? _GEN14443 : _GEN6834;
wire  _GEN14445 = io_x[42] ? _GEN14444 : _GEN6874;
wire  _GEN14446 = io_x[38] ? _GEN14445 : _GEN6871;
wire  _GEN14447 = io_x[10] ? _GEN14446 : _GEN7044;
wire  _GEN14448 = io_x[71] ? _GEN14447 : _GEN7203;
wire  _GEN14449 = io_x[70] ? _GEN7020 : _GEN14448;
wire  _GEN14450 = io_x[33] ? _GEN12627 : _GEN14449;
wire  _GEN14451 = io_x[21] ? _GEN14450 : _GEN12933;
wire  _GEN14452 = io_x[18] ? _GEN14451 : _GEN14439;
wire  _GEN14453 = io_x[20] ? _GEN14452 : _GEN14435;
wire  _GEN14454 = io_x[45] ? _GEN14453 : _GEN14429;
wire  _GEN14455 = io_x[28] ? _GEN14454 : _GEN14387;
wire  _GEN14456 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN14457 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14458 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14459 = io_x[6] ? _GEN14458 : _GEN14457;
wire  _GEN14460 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN14461 = io_x[2] ? _GEN6837 : _GEN14460;
wire  _GEN14462 = io_x[6] ? _GEN6850 : _GEN14461;
wire  _GEN14463 = io_x[41] ? _GEN14462 : _GEN14459;
wire  _GEN14464 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14465 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14466 = io_x[6] ? _GEN14465 : _GEN14464;
wire  _GEN14467 = io_x[41] ? _GEN6836 : _GEN14466;
wire  _GEN14468 = io_x[14] ? _GEN14467 : _GEN14463;
wire  _GEN14469 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14470 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14471 = io_x[6] ? _GEN14470 : _GEN14469;
wire  _GEN14472 = io_x[41] ? _GEN6836 : _GEN14471;
wire  _GEN14473 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14474 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14475 = io_x[6] ? _GEN14474 : _GEN14473;
wire  _GEN14476 = io_x[41] ? _GEN6836 : _GEN14475;
wire  _GEN14477 = io_x[14] ? _GEN14476 : _GEN14472;
wire  _GEN14478 = io_x[0] ? _GEN14477 : _GEN14468;
wire  _GEN14479 = io_x[76] ? _GEN14478 : _GEN6834;
wire  _GEN14480 = io_x[42] ? _GEN14479 : _GEN14456;
wire  _GEN14481 = io_x[38] ? _GEN14480 : _GEN6871;
wire  _GEN14482 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14483 = io_x[6] ? _GEN6850 : _GEN14482;
wire  _GEN14484 = io_x[41] ? _GEN6836 : _GEN14483;
wire  _GEN14485 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14486 = io_x[6] ? _GEN6840 : _GEN14485;
wire  _GEN14487 = io_x[41] ? _GEN6836 : _GEN14486;
wire  _GEN14488 = io_x[14] ? _GEN14487 : _GEN14484;
wire  _GEN14489 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14490 = io_x[6] ? _GEN6850 : _GEN14489;
wire  _GEN14491 = io_x[41] ? _GEN6836 : _GEN14490;
wire  _GEN14492 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14493 = io_x[41] ? _GEN6836 : _GEN14492;
wire  _GEN14494 = io_x[14] ? _GEN14493 : _GEN14491;
wire  _GEN14495 = io_x[0] ? _GEN14494 : _GEN14488;
wire  _GEN14496 = io_x[76] ? _GEN14495 : _GEN6834;
wire  _GEN14497 = io_x[42] ? _GEN14496 : _GEN6874;
wire  _GEN14498 = io_x[38] ? _GEN14497 : _GEN6871;
wire  _GEN14499 = io_x[10] ? _GEN14498 : _GEN14481;
wire  _GEN14500 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14501 = io_x[6] ? _GEN6840 : _GEN14500;
wire  _GEN14502 = io_x[41] ? _GEN14501 : _GEN6836;
wire  _GEN14503 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14504 = io_x[6] ? _GEN6850 : _GEN14503;
wire  _GEN14505 = io_x[41] ? _GEN14504 : _GEN6836;
wire  _GEN14506 = io_x[14] ? _GEN14505 : _GEN14502;
wire  _GEN14507 = io_x[0] ? _GEN14506 : _GEN6845;
wire  _GEN14508 = io_x[76] ? _GEN14507 : _GEN6834;
wire  _GEN14509 = io_x[42] ? _GEN6874 : _GEN14508;
wire  _GEN14510 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN14511 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN14512 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14513 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14514 = io_x[6] ? _GEN14513 : _GEN14512;
wire  _GEN14515 = io_x[41] ? _GEN6836 : _GEN14514;
wire  _GEN14516 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14517 = io_x[41] ? _GEN6836 : _GEN14516;
wire  _GEN14518 = io_x[14] ? _GEN14517 : _GEN14515;
wire  _GEN14519 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14520 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14521 = io_x[6] ? _GEN14520 : _GEN14519;
wire  _GEN14522 = io_x[41] ? _GEN6836 : _GEN14521;
wire  _GEN14523 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14524 = io_x[6] ? _GEN6850 : _GEN14523;
wire  _GEN14525 = io_x[41] ? _GEN6836 : _GEN14524;
wire  _GEN14526 = io_x[14] ? _GEN14525 : _GEN14522;
wire  _GEN14527 = io_x[0] ? _GEN14526 : _GEN14518;
wire  _GEN14528 = io_x[76] ? _GEN14527 : _GEN14511;
wire  _GEN14529 = io_x[42] ? _GEN14528 : _GEN14510;
wire  _GEN14530 = io_x[38] ? _GEN14529 : _GEN14509;
wire  _GEN14531 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14532 = io_x[6] ? _GEN6840 : _GEN14531;
wire  _GEN14533 = io_x[41] ? _GEN14532 : _GEN6836;
wire  _GEN14534 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14535 = io_x[6] ? _GEN14534 : _GEN6840;
wire  _GEN14536 = io_x[41] ? _GEN14535 : _GEN6836;
wire  _GEN14537 = io_x[14] ? _GEN14536 : _GEN14533;
wire  _GEN14538 = io_x[0] ? _GEN14537 : _GEN6845;
wire  _GEN14539 = io_x[76] ? _GEN14538 : _GEN6834;
wire  _GEN14540 = io_x[42] ? _GEN6874 : _GEN14539;
wire  _GEN14541 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN14542 = io_x[0] ? _GEN6845 : _GEN14541;
wire  _GEN14543 = io_x[76] ? _GEN14542 : _GEN6833;
wire  _GEN14544 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14545 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14546 = io_x[6] ? _GEN14545 : _GEN14544;
wire  _GEN14547 = io_x[41] ? _GEN6836 : _GEN14546;
wire  _GEN14548 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14549 = io_x[6] ? _GEN6840 : _GEN14548;
wire  _GEN14550 = io_x[41] ? _GEN6836 : _GEN14549;
wire  _GEN14551 = io_x[14] ? _GEN14550 : _GEN14547;
wire  _GEN14552 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14553 = io_x[41] ? _GEN6836 : _GEN14552;
wire  _GEN14554 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14555 = io_x[41] ? _GEN6836 : _GEN14554;
wire  _GEN14556 = io_x[14] ? _GEN14555 : _GEN14553;
wire  _GEN14557 = io_x[0] ? _GEN14556 : _GEN14551;
wire  _GEN14558 = io_x[76] ? _GEN14557 : _GEN6833;
wire  _GEN14559 = io_x[42] ? _GEN14558 : _GEN14543;
wire  _GEN14560 = io_x[38] ? _GEN14559 : _GEN14540;
wire  _GEN14561 = io_x[10] ? _GEN14560 : _GEN14530;
wire  _GEN14562 = io_x[71] ? _GEN14561 : _GEN14499;
wire  _GEN14563 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14564 = io_x[41] ? _GEN14563 : _GEN6836;
wire  _GEN14565 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14566 = io_x[41] ? _GEN14565 : _GEN6836;
wire  _GEN14567 = io_x[14] ? _GEN14566 : _GEN14564;
wire  _GEN14568 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14569 = io_x[41] ? _GEN14568 : _GEN6836;
wire  _GEN14570 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14571 = io_x[41] ? _GEN14570 : _GEN6836;
wire  _GEN14572 = io_x[14] ? _GEN14571 : _GEN14569;
wire  _GEN14573 = io_x[0] ? _GEN14572 : _GEN14567;
wire  _GEN14574 = io_x[76] ? _GEN14573 : _GEN6834;
wire  _GEN14575 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN14576 = io_x[42] ? _GEN14575 : _GEN14574;
wire  _GEN14577 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14578 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14579 = io_x[6] ? _GEN14578 : _GEN14577;
wire  _GEN14580 = io_x[41] ? _GEN14579 : _GEN6836;
wire  _GEN14581 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14582 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14583 = io_x[6] ? _GEN14582 : _GEN14581;
wire  _GEN14584 = io_x[41] ? _GEN14583 : _GEN6836;
wire  _GEN14585 = io_x[14] ? _GEN14584 : _GEN14580;
wire  _GEN14586 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14587 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14588 = io_x[6] ? _GEN14587 : _GEN14586;
wire  _GEN14589 = io_x[41] ? _GEN14588 : _GEN6836;
wire  _GEN14590 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14591 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14592 = io_x[6] ? _GEN14591 : _GEN14590;
wire  _GEN14593 = io_x[41] ? _GEN14592 : _GEN6836;
wire  _GEN14594 = io_x[14] ? _GEN14593 : _GEN14589;
wire  _GEN14595 = io_x[0] ? _GEN14594 : _GEN14585;
wire  _GEN14596 = io_x[76] ? _GEN14595 : _GEN6834;
wire  _GEN14597 = io_x[42] ? _GEN6874 : _GEN14596;
wire  _GEN14598 = io_x[38] ? _GEN14597 : _GEN14576;
wire  _GEN14599 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14600 = io_x[41] ? _GEN14599 : _GEN6836;
wire  _GEN14601 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14602 = io_x[41] ? _GEN14601 : _GEN6836;
wire  _GEN14603 = io_x[14] ? _GEN14602 : _GEN14600;
wire  _GEN14604 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14605 = io_x[41] ? _GEN14604 : _GEN6836;
wire  _GEN14606 = io_x[14] ? _GEN6843 : _GEN14605;
wire  _GEN14607 = io_x[0] ? _GEN14606 : _GEN14603;
wire  _GEN14608 = io_x[76] ? _GEN14607 : _GEN6834;
wire  _GEN14609 = io_x[42] ? _GEN6863 : _GEN14608;
wire  _GEN14610 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14611 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14612 = io_x[6] ? _GEN14611 : _GEN14610;
wire  _GEN14613 = io_x[41] ? _GEN14612 : _GEN6836;
wire  _GEN14614 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14615 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14616 = io_x[6] ? _GEN14615 : _GEN14614;
wire  _GEN14617 = io_x[41] ? _GEN14616 : _GEN6836;
wire  _GEN14618 = io_x[14] ? _GEN14617 : _GEN14613;
wire  _GEN14619 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14620 = io_x[6] ? _GEN6850 : _GEN14619;
wire  _GEN14621 = io_x[41] ? _GEN14620 : _GEN6836;
wire  _GEN14622 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14623 = io_x[6] ? _GEN6850 : _GEN14622;
wire  _GEN14624 = io_x[41] ? _GEN14623 : _GEN6836;
wire  _GEN14625 = io_x[14] ? _GEN14624 : _GEN14621;
wire  _GEN14626 = io_x[0] ? _GEN14625 : _GEN14618;
wire  _GEN14627 = io_x[76] ? _GEN14626 : _GEN6834;
wire  _GEN14628 = io_x[42] ? _GEN6874 : _GEN14627;
wire  _GEN14629 = io_x[38] ? _GEN14628 : _GEN14609;
wire  _GEN14630 = io_x[10] ? _GEN14629 : _GEN14598;
wire  _GEN14631 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14632 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14633 = io_x[6] ? _GEN14632 : _GEN14631;
wire  _GEN14634 = io_x[41] ? _GEN14633 : _GEN6836;
wire  _GEN14635 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14636 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14637 = io_x[6] ? _GEN14636 : _GEN14635;
wire  _GEN14638 = io_x[41] ? _GEN14637 : _GEN6836;
wire  _GEN14639 = io_x[14] ? _GEN14638 : _GEN14634;
wire  _GEN14640 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14641 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14642 = io_x[6] ? _GEN14641 : _GEN14640;
wire  _GEN14643 = io_x[41] ? _GEN14642 : _GEN6836;
wire  _GEN14644 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14645 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14646 = io_x[6] ? _GEN14645 : _GEN14644;
wire  _GEN14647 = io_x[41] ? _GEN14646 : _GEN6836;
wire  _GEN14648 = io_x[14] ? _GEN14647 : _GEN14643;
wire  _GEN14649 = io_x[0] ? _GEN14648 : _GEN14639;
wire  _GEN14650 = io_x[76] ? _GEN14649 : _GEN6833;
wire  _GEN14651 = io_x[42] ? _GEN14650 : _GEN6874;
wire  _GEN14652 = io_x[38] ? _GEN6871 : _GEN14651;
wire  _GEN14653 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14654 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14655 = io_x[6] ? _GEN14654 : _GEN14653;
wire  _GEN14656 = io_x[41] ? _GEN14655 : _GEN6836;
wire  _GEN14657 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14658 = io_x[6] ? _GEN6840 : _GEN14657;
wire  _GEN14659 = io_x[41] ? _GEN14658 : _GEN6836;
wire  _GEN14660 = io_x[14] ? _GEN14659 : _GEN14656;
wire  _GEN14661 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14662 = io_x[6] ? _GEN6850 : _GEN14661;
wire  _GEN14663 = io_x[41] ? _GEN14662 : _GEN6836;
wire  _GEN14664 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14665 = io_x[41] ? _GEN14664 : _GEN6836;
wire  _GEN14666 = io_x[14] ? _GEN14665 : _GEN14663;
wire  _GEN14667 = io_x[0] ? _GEN14666 : _GEN14660;
wire  _GEN14668 = io_x[76] ? _GEN14667 : _GEN6834;
wire  _GEN14669 = io_x[42] ? _GEN14668 : _GEN6874;
wire  _GEN14670 = io_x[38] ? _GEN6871 : _GEN14669;
wire  _GEN14671 = io_x[10] ? _GEN14670 : _GEN14652;
wire  _GEN14672 = io_x[71] ? _GEN14671 : _GEN14630;
wire  _GEN14673 = io_x[70] ? _GEN14672 : _GEN14562;
wire  _GEN14674 = io_x[33] ? _GEN12627 : _GEN14673;
wire  _GEN14675 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14676 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14677 = io_x[6] ? _GEN14676 : _GEN14675;
wire  _GEN14678 = io_x[41] ? _GEN6836 : _GEN14677;
wire  _GEN14679 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14680 = io_x[6] ? _GEN6840 : _GEN14679;
wire  _GEN14681 = io_x[41] ? _GEN6836 : _GEN14680;
wire  _GEN14682 = io_x[14] ? _GEN14681 : _GEN14678;
wire  _GEN14683 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14684 = io_x[6] ? _GEN6840 : _GEN14683;
wire  _GEN14685 = io_x[41] ? _GEN6836 : _GEN14684;
wire  _GEN14686 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14687 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14688 = io_x[6] ? _GEN14687 : _GEN14686;
wire  _GEN14689 = io_x[41] ? _GEN6836 : _GEN14688;
wire  _GEN14690 = io_x[14] ? _GEN14689 : _GEN14685;
wire  _GEN14691 = io_x[0] ? _GEN14690 : _GEN14682;
wire  _GEN14692 = io_x[76] ? _GEN14691 : _GEN6834;
wire  _GEN14693 = io_x[42] ? _GEN14692 : _GEN6874;
wire  _GEN14694 = io_x[38] ? _GEN14693 : _GEN6871;
wire  _GEN14695 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14696 = io_x[6] ? _GEN6840 : _GEN14695;
wire  _GEN14697 = io_x[41] ? _GEN6836 : _GEN14696;
wire  _GEN14698 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14699 = io_x[6] ? _GEN6850 : _GEN14698;
wire  _GEN14700 = io_x[41] ? _GEN6836 : _GEN14699;
wire  _GEN14701 = io_x[14] ? _GEN14700 : _GEN14697;
wire  _GEN14702 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14703 = io_x[6] ? _GEN6850 : _GEN14702;
wire  _GEN14704 = io_x[41] ? _GEN6836 : _GEN14703;
wire  _GEN14705 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14706 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14707 = io_x[6] ? _GEN14706 : _GEN14705;
wire  _GEN14708 = io_x[41] ? _GEN6836 : _GEN14707;
wire  _GEN14709 = io_x[14] ? _GEN14708 : _GEN14704;
wire  _GEN14710 = io_x[0] ? _GEN14709 : _GEN14701;
wire  _GEN14711 = io_x[76] ? _GEN14710 : _GEN6834;
wire  _GEN14712 = io_x[42] ? _GEN14711 : _GEN6863;
wire  _GEN14713 = io_x[38] ? _GEN14712 : _GEN6871;
wire  _GEN14714 = io_x[10] ? _GEN14713 : _GEN14694;
wire  _GEN14715 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN14716 = io_x[0] ? _GEN14715 : _GEN6845;
wire  _GEN14717 = io_x[76] ? _GEN14716 : _GEN6834;
wire  _GEN14718 = io_x[42] ? _GEN6874 : _GEN14717;
wire  _GEN14719 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14720 = io_x[6] ? _GEN6850 : _GEN14719;
wire  _GEN14721 = io_x[41] ? _GEN6836 : _GEN14720;
wire  _GEN14722 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14723 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14724 = io_x[6] ? _GEN14723 : _GEN14722;
wire  _GEN14725 = io_x[41] ? _GEN6836 : _GEN14724;
wire  _GEN14726 = io_x[14] ? _GEN14725 : _GEN14721;
wire  _GEN14727 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14728 = io_x[6] ? _GEN6840 : _GEN14727;
wire  _GEN14729 = io_x[41] ? _GEN6836 : _GEN14728;
wire  _GEN14730 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14731 = io_x[6] ? _GEN6850 : _GEN14730;
wire  _GEN14732 = io_x[41] ? _GEN6836 : _GEN14731;
wire  _GEN14733 = io_x[14] ? _GEN14732 : _GEN14729;
wire  _GEN14734 = io_x[0] ? _GEN14733 : _GEN14726;
wire  _GEN14735 = io_x[76] ? _GEN14734 : _GEN6834;
wire  _GEN14736 = io_x[42] ? _GEN14735 : _GEN6863;
wire  _GEN14737 = io_x[38] ? _GEN14736 : _GEN14718;
wire  _GEN14738 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN14739 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14740 = io_x[6] ? _GEN6840 : _GEN14739;
wire  _GEN14741 = io_x[41] ? _GEN6836 : _GEN14740;
wire  _GEN14742 = io_x[14] ? _GEN14741 : _GEN6843;
wire  _GEN14743 = io_x[0] ? _GEN14742 : _GEN6845;
wire  _GEN14744 = io_x[76] ? _GEN14743 : _GEN6834;
wire  _GEN14745 = io_x[42] ? _GEN14744 : _GEN14738;
wire  _GEN14746 = io_x[38] ? _GEN14745 : _GEN7036;
wire  _GEN14747 = io_x[10] ? _GEN14746 : _GEN14737;
wire  _GEN14748 = io_x[71] ? _GEN14747 : _GEN14714;
wire  _GEN14749 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14750 = io_x[41] ? _GEN14749 : _GEN6836;
wire  _GEN14751 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14752 = io_x[41] ? _GEN14751 : _GEN6836;
wire  _GEN14753 = io_x[14] ? _GEN14752 : _GEN14750;
wire  _GEN14754 = io_x[0] ? _GEN14753 : _GEN6845;
wire  _GEN14755 = io_x[76] ? _GEN14754 : _GEN6834;
wire  _GEN14756 = io_x[42] ? _GEN6874 : _GEN14755;
wire  _GEN14757 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14758 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14759 = io_x[6] ? _GEN14758 : _GEN14757;
wire  _GEN14760 = io_x[41] ? _GEN14759 : _GEN6836;
wire  _GEN14761 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14762 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14763 = io_x[6] ? _GEN14762 : _GEN14761;
wire  _GEN14764 = io_x[41] ? _GEN14763 : _GEN6836;
wire  _GEN14765 = io_x[14] ? _GEN14764 : _GEN14760;
wire  _GEN14766 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14767 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14768 = io_x[6] ? _GEN14767 : _GEN14766;
wire  _GEN14769 = io_x[41] ? _GEN14768 : _GEN6836;
wire  _GEN14770 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14771 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14772 = io_x[6] ? _GEN14771 : _GEN14770;
wire  _GEN14773 = io_x[41] ? _GEN14772 : _GEN6836;
wire  _GEN14774 = io_x[14] ? _GEN14773 : _GEN14769;
wire  _GEN14775 = io_x[0] ? _GEN14774 : _GEN14765;
wire  _GEN14776 = io_x[76] ? _GEN14775 : _GEN6834;
wire  _GEN14777 = io_x[42] ? _GEN6874 : _GEN14776;
wire  _GEN14778 = io_x[38] ? _GEN14777 : _GEN14756;
wire  _GEN14779 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14780 = io_x[41] ? _GEN14779 : _GEN6836;
wire  _GEN14781 = io_x[14] ? _GEN6843 : _GEN14780;
wire  _GEN14782 = io_x[0] ? _GEN14781 : _GEN6845;
wire  _GEN14783 = io_x[76] ? _GEN14782 : _GEN6834;
wire  _GEN14784 = io_x[42] ? _GEN6874 : _GEN14783;
wire  _GEN14785 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14786 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14787 = io_x[6] ? _GEN14786 : _GEN14785;
wire  _GEN14788 = io_x[41] ? _GEN14787 : _GEN6836;
wire  _GEN14789 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14790 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14791 = io_x[6] ? _GEN14790 : _GEN14789;
wire  _GEN14792 = io_x[41] ? _GEN14791 : _GEN6836;
wire  _GEN14793 = io_x[14] ? _GEN14792 : _GEN14788;
wire  _GEN14794 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14795 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14796 = io_x[6] ? _GEN14795 : _GEN14794;
wire  _GEN14797 = io_x[41] ? _GEN14796 : _GEN6836;
wire  _GEN14798 = io_x[14] ? _GEN6856 : _GEN14797;
wire  _GEN14799 = io_x[0] ? _GEN14798 : _GEN14793;
wire  _GEN14800 = io_x[76] ? _GEN14799 : _GEN6834;
wire  _GEN14801 = io_x[42] ? _GEN6874 : _GEN14800;
wire  _GEN14802 = io_x[38] ? _GEN14801 : _GEN14784;
wire  _GEN14803 = io_x[10] ? _GEN14802 : _GEN14778;
wire  _GEN14804 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14805 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14806 = io_x[6] ? _GEN14805 : _GEN14804;
wire  _GEN14807 = io_x[41] ? _GEN14806 : _GEN6836;
wire  _GEN14808 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14809 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14810 = io_x[6] ? _GEN14809 : _GEN14808;
wire  _GEN14811 = io_x[41] ? _GEN14810 : _GEN6836;
wire  _GEN14812 = io_x[14] ? _GEN14811 : _GEN14807;
wire  _GEN14813 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14814 = io_x[6] ? _GEN6840 : _GEN14813;
wire  _GEN14815 = io_x[41] ? _GEN14814 : _GEN6836;
wire  _GEN14816 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14817 = io_x[41] ? _GEN14816 : _GEN6836;
wire  _GEN14818 = io_x[14] ? _GEN14817 : _GEN14815;
wire  _GEN14819 = io_x[0] ? _GEN14818 : _GEN14812;
wire  _GEN14820 = io_x[76] ? _GEN14819 : _GEN6834;
wire  _GEN14821 = io_x[42] ? _GEN14820 : _GEN6874;
wire  _GEN14822 = io_x[38] ? _GEN6871 : _GEN14821;
wire  _GEN14823 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14824 = io_x[6] ? _GEN6850 : _GEN14823;
wire  _GEN14825 = io_x[41] ? _GEN14824 : _GEN6836;
wire  _GEN14826 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14827 = io_x[41] ? _GEN14826 : _GEN6836;
wire  _GEN14828 = io_x[14] ? _GEN14827 : _GEN14825;
wire  _GEN14829 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14830 = io_x[41] ? _GEN14829 : _GEN6836;
wire  _GEN14831 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14832 = io_x[6] ? _GEN6850 : _GEN14831;
wire  _GEN14833 = io_x[41] ? _GEN14832 : _GEN6836;
wire  _GEN14834 = io_x[14] ? _GEN14833 : _GEN14830;
wire  _GEN14835 = io_x[0] ? _GEN14834 : _GEN14828;
wire  _GEN14836 = io_x[76] ? _GEN14835 : _GEN6833;
wire  _GEN14837 = io_x[42] ? _GEN14836 : _GEN6874;
wire  _GEN14838 = io_x[38] ? _GEN6871 : _GEN14837;
wire  _GEN14839 = io_x[10] ? _GEN14838 : _GEN14822;
wire  _GEN14840 = io_x[71] ? _GEN14839 : _GEN14803;
wire  _GEN14841 = io_x[70] ? _GEN14840 : _GEN14748;
wire  _GEN14842 = io_x[33] ? _GEN12641 : _GEN14841;
wire  _GEN14843 = io_x[21] ? _GEN14842 : _GEN14674;
wire  _GEN14844 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14845 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14846 = io_x[6] ? _GEN14845 : _GEN14844;
wire  _GEN14847 = io_x[41] ? _GEN6836 : _GEN14846;
wire  _GEN14848 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14849 = io_x[6] ? _GEN14848 : _GEN6840;
wire  _GEN14850 = io_x[41] ? _GEN6836 : _GEN14849;
wire  _GEN14851 = io_x[14] ? _GEN14850 : _GEN14847;
wire  _GEN14852 = io_x[0] ? _GEN6845 : _GEN14851;
wire  _GEN14853 = io_x[76] ? _GEN14852 : _GEN6833;
wire  _GEN14854 = io_x[42] ? _GEN14853 : _GEN6874;
wire  _GEN14855 = io_x[38] ? _GEN14854 : _GEN6871;
wire  _GEN14856 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14857 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14858 = io_x[6] ? _GEN14857 : _GEN14856;
wire  _GEN14859 = io_x[41] ? _GEN6836 : _GEN14858;
wire  _GEN14860 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14861 = io_x[6] ? _GEN6840 : _GEN14860;
wire  _GEN14862 = io_x[41] ? _GEN6836 : _GEN14861;
wire  _GEN14863 = io_x[14] ? _GEN14862 : _GEN14859;
wire  _GEN14864 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14865 = io_x[41] ? _GEN6836 : _GEN14864;
wire  _GEN14866 = io_x[14] ? _GEN6843 : _GEN14865;
wire  _GEN14867 = io_x[0] ? _GEN14866 : _GEN14863;
wire  _GEN14868 = io_x[76] ? _GEN14867 : _GEN6834;
wire  _GEN14869 = io_x[42] ? _GEN14868 : _GEN6874;
wire  _GEN14870 = io_x[38] ? _GEN14869 : _GEN6871;
wire  _GEN14871 = io_x[10] ? _GEN14870 : _GEN14855;
wire  _GEN14872 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN14873 = io_x[76] ? _GEN6834 : _GEN14872;
wire  _GEN14874 = io_x[42] ? _GEN6874 : _GEN14873;
wire  _GEN14875 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14876 = io_x[6] ? _GEN6850 : _GEN14875;
wire  _GEN14877 = io_x[41] ? _GEN6836 : _GEN14876;
wire  _GEN14878 = io_x[14] ? _GEN6843 : _GEN14877;
wire  _GEN14879 = io_x[0] ? _GEN6845 : _GEN14878;
wire  _GEN14880 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14881 = io_x[6] ? _GEN6850 : _GEN14880;
wire  _GEN14882 = io_x[41] ? _GEN14881 : _GEN6836;
wire  _GEN14883 = io_x[14] ? _GEN6843 : _GEN14882;
wire  _GEN14884 = io_x[0] ? _GEN6845 : _GEN14883;
wire  _GEN14885 = io_x[76] ? _GEN14884 : _GEN14879;
wire  _GEN14886 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14887 = io_x[6] ? _GEN6850 : _GEN14886;
wire  _GEN14888 = io_x[41] ? _GEN14887 : _GEN6836;
wire  _GEN14889 = io_x[14] ? _GEN6843 : _GEN14888;
wire  _GEN14890 = io_x[0] ? _GEN6845 : _GEN14889;
wire  _GEN14891 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14892 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14893 = io_x[6] ? _GEN14892 : _GEN14891;
wire  _GEN14894 = io_x[41] ? _GEN6836 : _GEN14893;
wire  _GEN14895 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14896 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14897 = io_x[6] ? _GEN14896 : _GEN14895;
wire  _GEN14898 = io_x[41] ? _GEN6836 : _GEN14897;
wire  _GEN14899 = io_x[14] ? _GEN14898 : _GEN14894;
wire  _GEN14900 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14901 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14902 = io_x[6] ? _GEN14901 : _GEN14900;
wire  _GEN14903 = io_x[41] ? _GEN6836 : _GEN14902;
wire  _GEN14904 = io_x[14] ? _GEN6856 : _GEN14903;
wire  _GEN14905 = io_x[0] ? _GEN14904 : _GEN14899;
wire  _GEN14906 = io_x[76] ? _GEN14905 : _GEN14890;
wire  _GEN14907 = io_x[42] ? _GEN14906 : _GEN14885;
wire  _GEN14908 = io_x[38] ? _GEN14907 : _GEN14874;
wire  _GEN14909 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14910 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14911 = io_x[6] ? _GEN14910 : _GEN14909;
wire  _GEN14912 = io_x[41] ? _GEN6836 : _GEN14911;
wire  _GEN14913 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14914 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14915 = io_x[6] ? _GEN14914 : _GEN14913;
wire  _GEN14916 = io_x[41] ? _GEN6836 : _GEN14915;
wire  _GEN14917 = io_x[14] ? _GEN14916 : _GEN14912;
wire  _GEN14918 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14919 = io_x[6] ? _GEN14918 : _GEN6850;
wire  _GEN14920 = io_x[41] ? _GEN6836 : _GEN14919;
wire  _GEN14921 = io_x[14] ? _GEN6856 : _GEN14920;
wire  _GEN14922 = io_x[0] ? _GEN14921 : _GEN14917;
wire  _GEN14923 = io_x[76] ? _GEN14922 : _GEN6834;
wire  _GEN14924 = io_x[42] ? _GEN14923 : _GEN6863;
wire  _GEN14925 = io_x[38] ? _GEN14924 : _GEN6871;
wire  _GEN14926 = io_x[10] ? _GEN14925 : _GEN14908;
wire  _GEN14927 = io_x[71] ? _GEN14926 : _GEN14871;
wire  _GEN14928 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14929 = io_x[41] ? _GEN14928 : _GEN6836;
wire  _GEN14930 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14931 = io_x[41] ? _GEN14930 : _GEN6836;
wire  _GEN14932 = io_x[14] ? _GEN14931 : _GEN14929;
wire  _GEN14933 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14934 = io_x[41] ? _GEN14933 : _GEN6836;
wire  _GEN14935 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14936 = io_x[41] ? _GEN14935 : _GEN6836;
wire  _GEN14937 = io_x[14] ? _GEN14936 : _GEN14934;
wire  _GEN14938 = io_x[0] ? _GEN14937 : _GEN14932;
wire  _GEN14939 = io_x[76] ? _GEN14938 : _GEN6833;
wire  _GEN14940 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN14941 = io_x[14] ? _GEN6843 : _GEN14940;
wire  _GEN14942 = io_x[0] ? _GEN6845 : _GEN14941;
wire  _GEN14943 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN14944 = io_x[2] ? _GEN6837 : _GEN14943;
wire  _GEN14945 = io_x[6] ? _GEN6850 : _GEN14944;
wire  _GEN14946 = io_x[41] ? _GEN14945 : _GEN6836;
wire  _GEN14947 = io_x[14] ? _GEN6843 : _GEN14946;
wire  _GEN14948 = io_x[0] ? _GEN6845 : _GEN14947;
wire  _GEN14949 = io_x[76] ? _GEN14948 : _GEN14942;
wire  _GEN14950 = io_x[42] ? _GEN14949 : _GEN14939;
wire  _GEN14951 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14952 = io_x[6] ? _GEN6850 : _GEN14951;
wire  _GEN14953 = io_x[41] ? _GEN14952 : _GEN6836;
wire  _GEN14954 = io_x[14] ? _GEN6843 : _GEN14953;
wire  _GEN14955 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN14956 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14957 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14958 = io_x[6] ? _GEN14957 : _GEN14956;
wire  _GEN14959 = io_x[41] ? _GEN14958 : _GEN14955;
wire  _GEN14960 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14961 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14962 = io_x[6] ? _GEN14961 : _GEN14960;
wire  _GEN14963 = io_x[41] ? _GEN14962 : _GEN6836;
wire  _GEN14964 = io_x[14] ? _GEN14963 : _GEN14959;
wire  _GEN14965 = io_x[0] ? _GEN14964 : _GEN14954;
wire  _GEN14966 = io_x[76] ? _GEN14965 : _GEN6834;
wire  _GEN14967 = io_x[42] ? _GEN6874 : _GEN14966;
wire  _GEN14968 = io_x[38] ? _GEN14967 : _GEN14950;
wire  _GEN14969 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14970 = io_x[41] ? _GEN14969 : _GEN6836;
wire  _GEN14971 = io_x[14] ? _GEN6856 : _GEN14970;
wire  _GEN14972 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN14973 = io_x[41] ? _GEN14972 : _GEN6836;
wire  _GEN14974 = io_x[14] ? _GEN6856 : _GEN14973;
wire  _GEN14975 = io_x[0] ? _GEN14974 : _GEN14971;
wire  _GEN14976 = io_x[76] ? _GEN14975 : _GEN6834;
wire  _GEN14977 = io_x[42] ? _GEN6874 : _GEN14976;
wire  _GEN14978 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14979 = io_x[6] ? _GEN6840 : _GEN14978;
wire  _GEN14980 = io_x[41] ? _GEN14979 : _GEN6836;
wire  _GEN14981 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14982 = io_x[6] ? _GEN6850 : _GEN14981;
wire  _GEN14983 = io_x[41] ? _GEN14982 : _GEN6836;
wire  _GEN14984 = io_x[14] ? _GEN14983 : _GEN14980;
wire  _GEN14985 = io_x[0] ? _GEN14984 : _GEN6858;
wire  _GEN14986 = io_x[76] ? _GEN14985 : _GEN6834;
wire  _GEN14987 = io_x[42] ? _GEN6874 : _GEN14986;
wire  _GEN14988 = io_x[38] ? _GEN14987 : _GEN14977;
wire  _GEN14989 = io_x[10] ? _GEN14988 : _GEN14968;
wire  _GEN14990 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14991 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14992 = io_x[6] ? _GEN14991 : _GEN14990;
wire  _GEN14993 = io_x[41] ? _GEN14992 : _GEN6836;
wire  _GEN14994 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN14995 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN14996 = io_x[6] ? _GEN14995 : _GEN14994;
wire  _GEN14997 = io_x[41] ? _GEN14996 : _GEN6836;
wire  _GEN14998 = io_x[14] ? _GEN14997 : _GEN14993;
wire  _GEN14999 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15000 = io_x[41] ? _GEN14999 : _GEN6836;
wire  _GEN15001 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15002 = io_x[41] ? _GEN15001 : _GEN6836;
wire  _GEN15003 = io_x[14] ? _GEN15002 : _GEN15000;
wire  _GEN15004 = io_x[0] ? _GEN15003 : _GEN14998;
wire  _GEN15005 = io_x[76] ? _GEN15004 : _GEN6834;
wire  _GEN15006 = io_x[42] ? _GEN15005 : _GEN6863;
wire  _GEN15007 = io_x[38] ? _GEN6871 : _GEN15006;
wire  _GEN15008 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15009 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15010 = io_x[6] ? _GEN15009 : _GEN15008;
wire  _GEN15011 = io_x[41] ? _GEN15010 : _GEN6836;
wire  _GEN15012 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15013 = io_x[6] ? _GEN6840 : _GEN15012;
wire  _GEN15014 = io_x[41] ? _GEN15013 : _GEN6836;
wire  _GEN15015 = io_x[14] ? _GEN15014 : _GEN15011;
wire  _GEN15016 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15017 = io_x[0] ? _GEN15016 : _GEN15015;
wire  _GEN15018 = io_x[76] ? _GEN15017 : _GEN6834;
wire  _GEN15019 = io_x[42] ? _GEN15018 : _GEN6874;
wire  _GEN15020 = io_x[38] ? _GEN6871 : _GEN15019;
wire  _GEN15021 = io_x[10] ? _GEN15020 : _GEN15007;
wire  _GEN15022 = io_x[71] ? _GEN15021 : _GEN14989;
wire  _GEN15023 = io_x[70] ? _GEN15022 : _GEN14927;
wire  _GEN15024 = io_x[33] ? _GEN12641 : _GEN15023;
wire  _GEN15025 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN15026 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN15027 = io_x[76] ? _GEN15026 : _GEN6833;
wire  _GEN15028 = io_x[42] ? _GEN15027 : _GEN15025;
wire  _GEN15029 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15030 = io_x[6] ? _GEN6840 : _GEN15029;
wire  _GEN15031 = io_x[41] ? _GEN6924 : _GEN15030;
wire  _GEN15032 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15033 = io_x[6] ? _GEN6850 : _GEN15032;
wire  _GEN15034 = io_x[41] ? _GEN6836 : _GEN15033;
wire  _GEN15035 = io_x[14] ? _GEN15034 : _GEN15031;
wire  _GEN15036 = io_x[0] ? _GEN6858 : _GEN15035;
wire  _GEN15037 = io_x[76] ? _GEN15036 : _GEN6834;
wire  _GEN15038 = io_x[42] ? _GEN15037 : _GEN6874;
wire  _GEN15039 = io_x[38] ? _GEN15038 : _GEN15028;
wire  _GEN15040 = io_x[10] ? _GEN7094 : _GEN15039;
wire  _GEN15041 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15042 = io_x[41] ? _GEN15041 : _GEN6836;
wire  _GEN15043 = io_x[14] ? _GEN15042 : _GEN6843;
wire  _GEN15044 = io_x[0] ? _GEN15043 : _GEN6858;
wire  _GEN15045 = io_x[76] ? _GEN6834 : _GEN15044;
wire  _GEN15046 = io_x[42] ? _GEN6874 : _GEN15045;
wire  _GEN15047 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN15048 = io_x[0] ? _GEN6845 : _GEN15047;
wire  _GEN15049 = io_x[76] ? _GEN6834 : _GEN15048;
wire  _GEN15050 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15051 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15052 = io_x[6] ? _GEN15051 : _GEN15050;
wire  _GEN15053 = io_x[41] ? _GEN6836 : _GEN15052;
wire  _GEN15054 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15055 = io_x[6] ? _GEN6850 : _GEN15054;
wire  _GEN15056 = io_x[41] ? _GEN6836 : _GEN15055;
wire  _GEN15057 = io_x[14] ? _GEN15056 : _GEN15053;
wire  _GEN15058 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15059 = io_x[41] ? _GEN6836 : _GEN15058;
wire  _GEN15060 = io_x[14] ? _GEN15059 : _GEN6856;
wire  _GEN15061 = io_x[0] ? _GEN15060 : _GEN15057;
wire  _GEN15062 = io_x[76] ? _GEN15061 : _GEN6834;
wire  _GEN15063 = io_x[42] ? _GEN15062 : _GEN15049;
wire  _GEN15064 = io_x[38] ? _GEN15063 : _GEN15046;
wire  _GEN15065 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15066 = io_x[6] ? _GEN6840 : _GEN15065;
wire  _GEN15067 = io_x[41] ? _GEN6836 : _GEN15066;
wire  _GEN15068 = io_x[14] ? _GEN6843 : _GEN15067;
wire  _GEN15069 = io_x[0] ? _GEN6845 : _GEN15068;
wire  _GEN15070 = io_x[76] ? _GEN15069 : _GEN6834;
wire  _GEN15071 = io_x[42] ? _GEN15070 : _GEN6874;
wire  _GEN15072 = io_x[38] ? _GEN15071 : _GEN6871;
wire  _GEN15073 = io_x[10] ? _GEN15072 : _GEN15064;
wire  _GEN15074 = io_x[71] ? _GEN15073 : _GEN15040;
wire  _GEN15075 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15076 = io_x[0] ? _GEN15075 : _GEN6845;
wire  _GEN15077 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15078 = io_x[41] ? _GEN15077 : _GEN6836;
wire  _GEN15079 = io_x[14] ? _GEN15078 : _GEN6856;
wire  _GEN15080 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN15081 = io_x[14] ? _GEN6843 : _GEN15080;
wire  _GEN15082 = io_x[0] ? _GEN15081 : _GEN15079;
wire  _GEN15083 = io_x[76] ? _GEN15082 : _GEN15076;
wire  _GEN15084 = io_x[42] ? _GEN6874 : _GEN15083;
wire  _GEN15085 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15086 = io_x[41] ? _GEN15085 : _GEN6836;
wire  _GEN15087 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15088 = io_x[41] ? _GEN15087 : _GEN6836;
wire  _GEN15089 = io_x[14] ? _GEN15088 : _GEN15086;
wire  _GEN15090 = io_x[0] ? _GEN15089 : _GEN6845;
wire  _GEN15091 = io_x[76] ? _GEN15090 : _GEN6834;
wire  _GEN15092 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN15093 = io_x[42] ? _GEN15092 : _GEN15091;
wire  _GEN15094 = io_x[38] ? _GEN15093 : _GEN15084;
wire  _GEN15095 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15096 = io_x[41] ? _GEN15095 : _GEN6836;
wire  _GEN15097 = io_x[14] ? _GEN6843 : _GEN15096;
wire  _GEN15098 = io_x[0] ? _GEN6845 : _GEN15097;
wire  _GEN15099 = io_x[76] ? _GEN15098 : _GEN6834;
wire  _GEN15100 = io_x[42] ? _GEN6874 : _GEN15099;
wire  _GEN15101 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15102 = io_x[41] ? _GEN15101 : _GEN6836;
wire  _GEN15103 = io_x[14] ? _GEN15102 : _GEN6843;
wire  _GEN15104 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15105 = io_x[41] ? _GEN15104 : _GEN6836;
wire  _GEN15106 = io_x[14] ? _GEN6856 : _GEN15105;
wire  _GEN15107 = io_x[0] ? _GEN15106 : _GEN15103;
wire  _GEN15108 = io_x[76] ? _GEN15107 : _GEN6834;
wire  _GEN15109 = io_x[42] ? _GEN6874 : _GEN15108;
wire  _GEN15110 = io_x[38] ? _GEN15109 : _GEN15100;
wire  _GEN15111 = io_x[10] ? _GEN15110 : _GEN15094;
wire  _GEN15112 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15113 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15114 = io_x[6] ? _GEN15113 : _GEN15112;
wire  _GEN15115 = io_x[41] ? _GEN15114 : _GEN6836;
wire  _GEN15116 = io_x[14] ? _GEN6843 : _GEN15115;
wire  _GEN15117 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15118 = io_x[41] ? _GEN15117 : _GEN6836;
wire  _GEN15119 = io_x[14] ? _GEN6843 : _GEN15118;
wire  _GEN15120 = io_x[0] ? _GEN15119 : _GEN15116;
wire  _GEN15121 = io_x[76] ? _GEN15120 : _GEN6834;
wire  _GEN15122 = io_x[42] ? _GEN15121 : _GEN6874;
wire  _GEN15123 = io_x[38] ? _GEN6871 : _GEN15122;
wire  _GEN15124 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN15125 = io_x[42] ? _GEN15124 : _GEN6874;
wire  _GEN15126 = io_x[38] ? _GEN6871 : _GEN15125;
wire  _GEN15127 = io_x[10] ? _GEN15126 : _GEN15123;
wire  _GEN15128 = io_x[71] ? _GEN15127 : _GEN15111;
wire  _GEN15129 = io_x[70] ? _GEN15128 : _GEN15074;
wire  _GEN15130 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15131 = io_x[41] ? _GEN6836 : _GEN15130;
wire  _GEN15132 = io_x[14] ? _GEN15131 : _GEN6843;
wire  _GEN15133 = io_x[0] ? _GEN15132 : _GEN6845;
wire  _GEN15134 = io_x[76] ? _GEN6834 : _GEN15133;
wire  _GEN15135 = io_x[42] ? _GEN15134 : _GEN6874;
wire  _GEN15136 = io_x[38] ? _GEN6871 : _GEN15135;
wire  _GEN15137 = io_x[10] ? _GEN7044 : _GEN15136;
wire  _GEN15138 = io_x[71] ? _GEN7196 : _GEN15137;
wire  _GEN15139 = io_x[70] ? _GEN8474 : _GEN15138;
wire  _GEN15140 = io_x[33] ? _GEN15139 : _GEN15129;
wire  _GEN15141 = io_x[21] ? _GEN15140 : _GEN15024;
wire  _GEN15142 = io_x[18] ? _GEN15141 : _GEN14843;
wire  _GEN15143 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15144 = io_x[41] ? _GEN6836 : _GEN15143;
wire  _GEN15145 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15146 = io_x[41] ? _GEN6836 : _GEN15145;
wire  _GEN15147 = io_x[14] ? _GEN15146 : _GEN15144;
wire  _GEN15148 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15149 = io_x[41] ? _GEN6924 : _GEN15148;
wire  _GEN15150 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15151 = io_x[6] ? _GEN6850 : _GEN15150;
wire  _GEN15152 = io_x[41] ? _GEN6836 : _GEN15151;
wire  _GEN15153 = io_x[14] ? _GEN15152 : _GEN15149;
wire  _GEN15154 = io_x[0] ? _GEN15153 : _GEN15147;
wire  _GEN15155 = io_x[76] ? _GEN15154 : _GEN6834;
wire  _GEN15156 = io_x[42] ? _GEN15155 : _GEN6863;
wire  _GEN15157 = io_x[38] ? _GEN15156 : _GEN6871;
wire  _GEN15158 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15159 = io_x[6] ? _GEN6850 : _GEN15158;
wire  _GEN15160 = io_x[41] ? _GEN15159 : _GEN6836;
wire  _GEN15161 = io_x[14] ? _GEN15160 : _GEN6843;
wire  _GEN15162 = io_x[0] ? _GEN15161 : _GEN6845;
wire  _GEN15163 = io_x[76] ? _GEN6834 : _GEN15162;
wire  _GEN15164 = io_x[42] ? _GEN6863 : _GEN15163;
wire  _GEN15165 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15166 = io_x[41] ? _GEN6836 : _GEN15165;
wire  _GEN15167 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15168 = io_x[41] ? _GEN6836 : _GEN15167;
wire  _GEN15169 = io_x[14] ? _GEN15168 : _GEN15166;
wire  _GEN15170 = io_x[0] ? _GEN6858 : _GEN15169;
wire  _GEN15171 = io_x[76] ? _GEN15170 : _GEN6834;
wire  _GEN15172 = io_x[42] ? _GEN15171 : _GEN6874;
wire  _GEN15173 = io_x[38] ? _GEN15172 : _GEN15164;
wire  _GEN15174 = io_x[10] ? _GEN15173 : _GEN15157;
wire  _GEN15175 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN15176 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15177 = io_x[41] ? _GEN6836 : _GEN15176;
wire  _GEN15178 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15179 = io_x[41] ? _GEN6836 : _GEN15178;
wire  _GEN15180 = io_x[14] ? _GEN15179 : _GEN15177;
wire  _GEN15181 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15182 = io_x[6] ? _GEN6850 : _GEN15181;
wire  _GEN15183 = io_x[41] ? _GEN6836 : _GEN15182;
wire  _GEN15184 = io_x[14] ? _GEN6856 : _GEN15183;
wire  _GEN15185 = io_x[0] ? _GEN15184 : _GEN15180;
wire  _GEN15186 = io_x[76] ? _GEN15185 : _GEN6834;
wire  _GEN15187 = io_x[42] ? _GEN15186 : _GEN15175;
wire  _GEN15188 = io_x[38] ? _GEN15187 : _GEN6871;
wire  _GEN15189 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15190 = io_x[41] ? _GEN6836 : _GEN15189;
wire  _GEN15191 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15192 = io_x[41] ? _GEN6836 : _GEN15191;
wire  _GEN15193 = io_x[14] ? _GEN15192 : _GEN15190;
wire  _GEN15194 = io_x[0] ? _GEN6858 : _GEN15193;
wire  _GEN15195 = io_x[76] ? _GEN15194 : _GEN6834;
wire  _GEN15196 = io_x[42] ? _GEN15195 : _GEN6874;
wire  _GEN15197 = io_x[38] ? _GEN15196 : _GEN6871;
wire  _GEN15198 = io_x[10] ? _GEN15197 : _GEN15188;
wire  _GEN15199 = io_x[71] ? _GEN15198 : _GEN15174;
wire  _GEN15200 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15201 = io_x[41] ? _GEN15200 : _GEN6836;
wire  _GEN15202 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15203 = io_x[41] ? _GEN15202 : _GEN6836;
wire  _GEN15204 = io_x[14] ? _GEN15203 : _GEN15201;
wire  _GEN15205 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15206 = io_x[41] ? _GEN15205 : _GEN6836;
wire  _GEN15207 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15208 = io_x[41] ? _GEN15207 : _GEN6836;
wire  _GEN15209 = io_x[14] ? _GEN15208 : _GEN15206;
wire  _GEN15210 = io_x[0] ? _GEN15209 : _GEN15204;
wire  _GEN15211 = io_x[76] ? _GEN15210 : _GEN6834;
wire  _GEN15212 = io_x[42] ? _GEN6874 : _GEN15211;
wire  _GEN15213 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15214 = io_x[41] ? _GEN15213 : _GEN6836;
wire  _GEN15215 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15216 = io_x[6] ? _GEN6840 : _GEN15215;
wire  _GEN15217 = io_x[41] ? _GEN15216 : _GEN6836;
wire  _GEN15218 = io_x[14] ? _GEN15217 : _GEN15214;
wire  _GEN15219 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15220 = io_x[41] ? _GEN15219 : _GEN6836;
wire  _GEN15221 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15222 = io_x[41] ? _GEN15221 : _GEN6836;
wire  _GEN15223 = io_x[14] ? _GEN15222 : _GEN15220;
wire  _GEN15224 = io_x[0] ? _GEN15223 : _GEN15218;
wire  _GEN15225 = io_x[76] ? _GEN15224 : _GEN6834;
wire  _GEN15226 = io_x[42] ? _GEN6874 : _GEN15225;
wire  _GEN15227 = io_x[38] ? _GEN15226 : _GEN15212;
wire  _GEN15228 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15229 = io_x[41] ? _GEN15228 : _GEN6836;
wire  _GEN15230 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15231 = io_x[41] ? _GEN15230 : _GEN6836;
wire  _GEN15232 = io_x[14] ? _GEN15231 : _GEN15229;
wire  _GEN15233 = io_x[0] ? _GEN6858 : _GEN15232;
wire  _GEN15234 = io_x[76] ? _GEN15233 : _GEN6833;
wire  _GEN15235 = io_x[42] ? _GEN6874 : _GEN15234;
wire  _GEN15236 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15237 = io_x[6] ? _GEN6840 : _GEN15236;
wire  _GEN15238 = io_x[41] ? _GEN15237 : _GEN6836;
wire  _GEN15239 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15240 = io_x[41] ? _GEN15239 : _GEN6836;
wire  _GEN15241 = io_x[14] ? _GEN15240 : _GEN15238;
wire  _GEN15242 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15243 = io_x[41] ? _GEN15242 : _GEN6836;
wire  _GEN15244 = io_x[14] ? _GEN6843 : _GEN15243;
wire  _GEN15245 = io_x[0] ? _GEN15244 : _GEN15241;
wire  _GEN15246 = io_x[76] ? _GEN15245 : _GEN6833;
wire  _GEN15247 = io_x[42] ? _GEN6874 : _GEN15246;
wire  _GEN15248 = io_x[38] ? _GEN15247 : _GEN15235;
wire  _GEN15249 = io_x[10] ? _GEN15248 : _GEN15227;
wire  _GEN15250 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15251 = io_x[41] ? _GEN15250 : _GEN6836;
wire  _GEN15252 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15253 = io_x[41] ? _GEN15252 : _GEN6836;
wire  _GEN15254 = io_x[14] ? _GEN15253 : _GEN15251;
wire  _GEN15255 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15256 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15257 = io_x[6] ? _GEN15256 : _GEN15255;
wire  _GEN15258 = io_x[41] ? _GEN15257 : _GEN6836;
wire  _GEN15259 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15260 = io_x[6] ? _GEN6850 : _GEN15259;
wire  _GEN15261 = io_x[41] ? _GEN15260 : _GEN6836;
wire  _GEN15262 = io_x[14] ? _GEN15261 : _GEN15258;
wire  _GEN15263 = io_x[0] ? _GEN15262 : _GEN15254;
wire  _GEN15264 = io_x[76] ? _GEN15263 : _GEN6834;
wire  _GEN15265 = io_x[42] ? _GEN15264 : _GEN6874;
wire  _GEN15266 = io_x[38] ? _GEN6871 : _GEN15265;
wire  _GEN15267 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15268 = io_x[41] ? _GEN15267 : _GEN6836;
wire  _GEN15269 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15270 = io_x[41] ? _GEN15269 : _GEN6836;
wire  _GEN15271 = io_x[14] ? _GEN15270 : _GEN15268;
wire  _GEN15272 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15273 = io_x[6] ? _GEN15272 : _GEN6840;
wire  _GEN15274 = io_x[41] ? _GEN15273 : _GEN6836;
wire  _GEN15275 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15276 = io_x[6] ? _GEN6840 : _GEN15275;
wire  _GEN15277 = io_x[41] ? _GEN15276 : _GEN6836;
wire  _GEN15278 = io_x[14] ? _GEN15277 : _GEN15274;
wire  _GEN15279 = io_x[0] ? _GEN15278 : _GEN15271;
wire  _GEN15280 = io_x[76] ? _GEN15279 : _GEN6834;
wire  _GEN15281 = io_x[42] ? _GEN15280 : _GEN6863;
wire  _GEN15282 = io_x[38] ? _GEN6871 : _GEN15281;
wire  _GEN15283 = io_x[10] ? _GEN15282 : _GEN15266;
wire  _GEN15284 = io_x[71] ? _GEN15283 : _GEN15249;
wire  _GEN15285 = io_x[70] ? _GEN15284 : _GEN15199;
wire  _GEN15286 = io_x[33] ? _GEN12627 : _GEN15285;
wire  _GEN15287 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15288 = io_x[41] ? _GEN6836 : _GEN15287;
wire  _GEN15289 = io_x[14] ? _GEN15288 : _GEN6843;
wire  _GEN15290 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15291 = io_x[6] ? _GEN6850 : _GEN15290;
wire  _GEN15292 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15293 = io_x[6] ? _GEN6840 : _GEN15292;
wire  _GEN15294 = io_x[41] ? _GEN15293 : _GEN15291;
wire  _GEN15295 = io_x[14] ? _GEN6856 : _GEN15294;
wire  _GEN15296 = io_x[0] ? _GEN15295 : _GEN15289;
wire  _GEN15297 = io_x[76] ? _GEN15296 : _GEN6834;
wire  _GEN15298 = io_x[42] ? _GEN15297 : _GEN6863;
wire  _GEN15299 = io_x[38] ? _GEN15298 : _GEN7036;
wire  _GEN15300 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15301 = io_x[6] ? _GEN6850 : _GEN15300;
wire  _GEN15302 = io_x[41] ? _GEN6836 : _GEN15301;
wire  _GEN15303 = io_x[14] ? _GEN15302 : _GEN6856;
wire  _GEN15304 = io_x[0] ? _GEN6845 : _GEN15303;
wire  _GEN15305 = io_x[76] ? _GEN15304 : _GEN6834;
wire  _GEN15306 = io_x[42] ? _GEN15305 : _GEN6863;
wire  _GEN15307 = io_x[38] ? _GEN15306 : _GEN6871;
wire  _GEN15308 = io_x[10] ? _GEN15307 : _GEN15299;
wire  _GEN15309 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN15310 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN15311 = io_x[76] ? _GEN6834 : _GEN15310;
wire  _GEN15312 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15313 = io_x[6] ? _GEN15312 : _GEN6850;
wire  _GEN15314 = io_x[41] ? _GEN6836 : _GEN15313;
wire  _GEN15315 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15316 = io_x[41] ? _GEN6836 : _GEN15315;
wire  _GEN15317 = io_x[14] ? _GEN15316 : _GEN15314;
wire  _GEN15318 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15319 = io_x[0] ? _GEN15318 : _GEN15317;
wire  _GEN15320 = io_x[76] ? _GEN15319 : _GEN6834;
wire  _GEN15321 = io_x[42] ? _GEN15320 : _GEN15311;
wire  _GEN15322 = io_x[38] ? _GEN15321 : _GEN15309;
wire  _GEN15323 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN15324 = io_x[0] ? _GEN6858 : _GEN15323;
wire  _GEN15325 = io_x[76] ? _GEN15324 : _GEN6834;
wire  _GEN15326 = io_x[42] ? _GEN15325 : _GEN6863;
wire  _GEN15327 = io_x[38] ? _GEN15326 : _GEN6871;
wire  _GEN15328 = io_x[10] ? _GEN15327 : _GEN15322;
wire  _GEN15329 = io_x[71] ? _GEN15328 : _GEN15308;
wire  _GEN15330 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15331 = io_x[41] ? _GEN15330 : _GEN6836;
wire  _GEN15332 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15333 = io_x[41] ? _GEN15332 : _GEN6836;
wire  _GEN15334 = io_x[14] ? _GEN15333 : _GEN15331;
wire  _GEN15335 = io_x[0] ? _GEN6845 : _GEN15334;
wire  _GEN15336 = io_x[76] ? _GEN15335 : _GEN6833;
wire  _GEN15337 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15338 = io_x[41] ? _GEN15337 : _GEN6836;
wire  _GEN15339 = io_x[14] ? _GEN6843 : _GEN15338;
wire  _GEN15340 = io_x[0] ? _GEN6845 : _GEN15339;
wire  _GEN15341 = io_x[76] ? _GEN15340 : _GEN6834;
wire  _GEN15342 = io_x[42] ? _GEN15341 : _GEN15336;
wire  _GEN15343 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15344 = io_x[41] ? _GEN15343 : _GEN6836;
wire  _GEN15345 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15346 = io_x[41] ? _GEN15345 : _GEN6836;
wire  _GEN15347 = io_x[14] ? _GEN15346 : _GEN15344;
wire  _GEN15348 = io_x[0] ? _GEN6845 : _GEN15347;
wire  _GEN15349 = io_x[76] ? _GEN15348 : _GEN6834;
wire  _GEN15350 = io_x[42] ? _GEN6874 : _GEN15349;
wire  _GEN15351 = io_x[38] ? _GEN15350 : _GEN15342;
wire  _GEN15352 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15353 = io_x[41] ? _GEN15352 : _GEN6836;
wire  _GEN15354 = io_x[14] ? _GEN6856 : _GEN15353;
wire  _GEN15355 = io_x[0] ? _GEN6858 : _GEN15354;
wire  _GEN15356 = io_x[76] ? _GEN15355 : _GEN6834;
wire  _GEN15357 = io_x[42] ? _GEN6874 : _GEN15356;
wire  _GEN15358 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15359 = io_x[6] ? _GEN15358 : _GEN6850;
wire  _GEN15360 = io_x[41] ? _GEN15359 : _GEN6836;
wire  _GEN15361 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15362 = io_x[41] ? _GEN15361 : _GEN6836;
wire  _GEN15363 = io_x[14] ? _GEN15362 : _GEN15360;
wire  _GEN15364 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15365 = io_x[0] ? _GEN15364 : _GEN15363;
wire  _GEN15366 = io_x[76] ? _GEN15365 : _GEN6833;
wire  _GEN15367 = io_x[42] ? _GEN6874 : _GEN15366;
wire  _GEN15368 = io_x[38] ? _GEN15367 : _GEN15357;
wire  _GEN15369 = io_x[10] ? _GEN15368 : _GEN15351;
wire  _GEN15370 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN15371 = io_x[2] ? _GEN6837 : _GEN15370;
wire  _GEN15372 = io_x[6] ? _GEN6850 : _GEN15371;
wire  _GEN15373 = io_x[41] ? _GEN6836 : _GEN15372;
wire  _GEN15374 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15375 = io_x[6] ? _GEN6850 : _GEN15374;
wire  _GEN15376 = io_x[41] ? _GEN15375 : _GEN6836;
wire  _GEN15377 = io_x[14] ? _GEN15376 : _GEN15373;
wire  _GEN15378 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15379 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15380 = io_x[6] ? _GEN15379 : _GEN15378;
wire  _GEN15381 = io_x[41] ? _GEN15380 : _GEN6836;
wire  _GEN15382 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15383 = io_x[6] ? _GEN15382 : _GEN6840;
wire  _GEN15384 = io_x[41] ? _GEN15383 : _GEN6836;
wire  _GEN15385 = io_x[14] ? _GEN15384 : _GEN15381;
wire  _GEN15386 = io_x[0] ? _GEN15385 : _GEN15377;
wire  _GEN15387 = io_x[76] ? _GEN15386 : _GEN6834;
wire  _GEN15388 = io_x[42] ? _GEN15387 : _GEN6874;
wire  _GEN15389 = io_x[38] ? _GEN7036 : _GEN15388;
wire  _GEN15390 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15391 = io_x[0] ? _GEN15390 : _GEN6858;
wire  _GEN15392 = io_x[76] ? _GEN15391 : _GEN6834;
wire  _GEN15393 = io_x[42] ? _GEN15392 : _GEN6863;
wire  _GEN15394 = io_x[38] ? _GEN6871 : _GEN15393;
wire  _GEN15395 = io_x[10] ? _GEN15394 : _GEN15389;
wire  _GEN15396 = io_x[71] ? _GEN15395 : _GEN15369;
wire  _GEN15397 = io_x[70] ? _GEN15396 : _GEN15329;
wire  _GEN15398 = io_x[33] ? _GEN12641 : _GEN15397;
wire  _GEN15399 = io_x[21] ? _GEN15398 : _GEN15286;
wire  _GEN15400 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN15401 = io_x[76] ? _GEN15400 : _GEN6833;
wire  _GEN15402 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15403 = io_x[6] ? _GEN6850 : _GEN15402;
wire  _GEN15404 = io_x[41] ? _GEN15403 : _GEN6836;
wire  _GEN15405 = io_x[14] ? _GEN6843 : _GEN15404;
wire  _GEN15406 = io_x[0] ? _GEN15405 : _GEN6858;
wire  _GEN15407 = io_x[76] ? _GEN6834 : _GEN15406;
wire  _GEN15408 = io_x[42] ? _GEN15407 : _GEN15401;
wire  _GEN15409 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15410 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15411 = io_x[6] ? _GEN15410 : _GEN15409;
wire  _GEN15412 = io_x[41] ? _GEN6924 : _GEN15411;
wire  _GEN15413 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15414 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15415 = io_x[6] ? _GEN15414 : _GEN15413;
wire  _GEN15416 = io_x[41] ? _GEN6836 : _GEN15415;
wire  _GEN15417 = io_x[14] ? _GEN15416 : _GEN15412;
wire  _GEN15418 = io_x[0] ? _GEN6845 : _GEN15417;
wire  _GEN15419 = io_x[76] ? _GEN15418 : _GEN6834;
wire  _GEN15420 = io_x[42] ? _GEN15419 : _GEN6863;
wire  _GEN15421 = io_x[38] ? _GEN15420 : _GEN15408;
wire  _GEN15422 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15423 = io_x[41] ? _GEN15422 : _GEN6836;
wire  _GEN15424 = io_x[14] ? _GEN15423 : _GEN6843;
wire  _GEN15425 = io_x[0] ? _GEN15424 : _GEN6845;
wire  _GEN15426 = io_x[76] ? _GEN6834 : _GEN15425;
wire  _GEN15427 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15428 = io_x[41] ? _GEN6836 : _GEN15427;
wire  _GEN15429 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15430 = io_x[6] ? _GEN6850 : _GEN15429;
wire  _GEN15431 = io_x[41] ? _GEN6836 : _GEN15430;
wire  _GEN15432 = io_x[14] ? _GEN15431 : _GEN15428;
wire  _GEN15433 = io_x[0] ? _GEN6845 : _GEN15432;
wire  _GEN15434 = io_x[76] ? _GEN15433 : _GEN6834;
wire  _GEN15435 = io_x[42] ? _GEN15434 : _GEN15426;
wire  _GEN15436 = io_x[38] ? _GEN15435 : _GEN6871;
wire  _GEN15437 = io_x[10] ? _GEN15436 : _GEN15421;
wire  _GEN15438 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15439 = io_x[41] ? _GEN6836 : _GEN15438;
wire  _GEN15440 = io_x[14] ? _GEN6856 : _GEN15439;
wire  _GEN15441 = io_x[0] ? _GEN15440 : _GEN6858;
wire  _GEN15442 = io_x[76] ? _GEN6834 : _GEN15441;
wire  _GEN15443 = io_x[42] ? _GEN6874 : _GEN15442;
wire  _GEN15444 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15445 = io_x[6] ? _GEN6850 : _GEN15444;
wire  _GEN15446 = io_x[41] ? _GEN6924 : _GEN15445;
wire  _GEN15447 = io_x[14] ? _GEN6856 : _GEN15446;
wire  _GEN15448 = io_x[0] ? _GEN6845 : _GEN15447;
wire  _GEN15449 = io_x[76] ? _GEN6834 : _GEN15448;
wire  _GEN15450 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15451 = io_x[6] ? _GEN6840 : _GEN15450;
wire  _GEN15452 = io_x[41] ? _GEN6836 : _GEN15451;
wire  _GEN15453 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15454 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15455 = io_x[6] ? _GEN15454 : _GEN15453;
wire  _GEN15456 = io_x[41] ? _GEN6836 : _GEN15455;
wire  _GEN15457 = io_x[14] ? _GEN15456 : _GEN15452;
wire  _GEN15458 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15459 = io_x[6] ? _GEN15458 : _GEN6850;
wire  _GEN15460 = io_x[41] ? _GEN6836 : _GEN15459;
wire  _GEN15461 = io_x[14] ? _GEN6856 : _GEN15460;
wire  _GEN15462 = io_x[0] ? _GEN15461 : _GEN15457;
wire  _GEN15463 = io_x[76] ? _GEN15462 : _GEN6834;
wire  _GEN15464 = io_x[42] ? _GEN15463 : _GEN15449;
wire  _GEN15465 = io_x[38] ? _GEN15464 : _GEN15443;
wire  _GEN15466 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN15467 = io_x[0] ? _GEN6858 : _GEN15466;
wire  _GEN15468 = io_x[76] ? _GEN6834 : _GEN15467;
wire  _GEN15469 = io_x[42] ? _GEN6863 : _GEN15468;
wire  _GEN15470 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15471 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15472 = io_x[6] ? _GEN15471 : _GEN15470;
wire  _GEN15473 = io_x[41] ? _GEN6836 : _GEN15472;
wire  _GEN15474 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15475 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15476 = io_x[6] ? _GEN15475 : _GEN15474;
wire  _GEN15477 = io_x[41] ? _GEN6836 : _GEN15476;
wire  _GEN15478 = io_x[14] ? _GEN15477 : _GEN15473;
wire  _GEN15479 = io_x[0] ? _GEN6845 : _GEN15478;
wire  _GEN15480 = io_x[76] ? _GEN15479 : _GEN6834;
wire  _GEN15481 = io_x[42] ? _GEN15480 : _GEN6863;
wire  _GEN15482 = io_x[38] ? _GEN15481 : _GEN15469;
wire  _GEN15483 = io_x[10] ? _GEN15482 : _GEN15465;
wire  _GEN15484 = io_x[71] ? _GEN15483 : _GEN15437;
wire  _GEN15485 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15486 = io_x[41] ? _GEN15485 : _GEN6924;
wire  _GEN15487 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15488 = io_x[41] ? _GEN15487 : _GEN6836;
wire  _GEN15489 = io_x[14] ? _GEN15488 : _GEN15486;
wire  _GEN15490 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15491 = io_x[41] ? _GEN15490 : _GEN6836;
wire  _GEN15492 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15493 = io_x[41] ? _GEN15492 : _GEN6836;
wire  _GEN15494 = io_x[14] ? _GEN15493 : _GEN15491;
wire  _GEN15495 = io_x[0] ? _GEN15494 : _GEN15489;
wire  _GEN15496 = io_x[76] ? _GEN15495 : _GEN6834;
wire  _GEN15497 = io_x[42] ? _GEN6874 : _GEN15496;
wire  _GEN15498 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15499 = io_x[6] ? _GEN6840 : _GEN15498;
wire  _GEN15500 = io_x[41] ? _GEN15499 : _GEN6836;
wire  _GEN15501 = io_x[14] ? _GEN6843 : _GEN15500;
wire  _GEN15502 = io_x[0] ? _GEN15501 : _GEN6845;
wire  _GEN15503 = io_x[76] ? _GEN15502 : _GEN6834;
wire  _GEN15504 = io_x[42] ? _GEN6874 : _GEN15503;
wire  _GEN15505 = io_x[38] ? _GEN15504 : _GEN15497;
wire  _GEN15506 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15507 = io_x[41] ? _GEN15506 : _GEN6836;
wire  _GEN15508 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15509 = io_x[41] ? _GEN15508 : _GEN6836;
wire  _GEN15510 = io_x[14] ? _GEN15509 : _GEN15507;
wire  _GEN15511 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15512 = io_x[41] ? _GEN15511 : _GEN6836;
wire  _GEN15513 = io_x[14] ? _GEN6843 : _GEN15512;
wire  _GEN15514 = io_x[0] ? _GEN15513 : _GEN15510;
wire  _GEN15515 = io_x[76] ? _GEN15514 : _GEN6834;
wire  _GEN15516 = io_x[42] ? _GEN6863 : _GEN15515;
wire  _GEN15517 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15518 = io_x[6] ? _GEN6850 : _GEN15517;
wire  _GEN15519 = io_x[41] ? _GEN15518 : _GEN6836;
wire  _GEN15520 = io_x[14] ? _GEN6856 : _GEN15519;
wire  _GEN15521 = io_x[0] ? _GEN15520 : _GEN6858;
wire  _GEN15522 = io_x[76] ? _GEN15521 : _GEN6834;
wire  _GEN15523 = io_x[42] ? _GEN6874 : _GEN15522;
wire  _GEN15524 = io_x[38] ? _GEN15523 : _GEN15516;
wire  _GEN15525 = io_x[10] ? _GEN15524 : _GEN15505;
wire  _GEN15526 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15527 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15528 = io_x[6] ? _GEN15527 : _GEN15526;
wire  _GEN15529 = io_x[41] ? _GEN15528 : _GEN6836;
wire  _GEN15530 = io_x[14] ? _GEN6856 : _GEN15529;
wire  _GEN15531 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15532 = io_x[41] ? _GEN15531 : _GEN6836;
wire  _GEN15533 = io_x[14] ? _GEN15532 : _GEN6856;
wire  _GEN15534 = io_x[0] ? _GEN15533 : _GEN15530;
wire  _GEN15535 = io_x[76] ? _GEN15534 : _GEN6834;
wire  _GEN15536 = io_x[42] ? _GEN15535 : _GEN6874;
wire  _GEN15537 = io_x[38] ? _GEN6871 : _GEN15536;
wire  _GEN15538 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN15539 = io_x[76] ? _GEN15538 : _GEN6834;
wire  _GEN15540 = io_x[42] ? _GEN15539 : _GEN6874;
wire  _GEN15541 = io_x[38] ? _GEN6871 : _GEN15540;
wire  _GEN15542 = io_x[10] ? _GEN15541 : _GEN15537;
wire  _GEN15543 = io_x[71] ? _GEN15542 : _GEN15525;
wire  _GEN15544 = io_x[70] ? _GEN15543 : _GEN15484;
wire  _GEN15545 = io_x[33] ? _GEN12627 : _GEN15544;
wire  _GEN15546 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15547 = io_x[41] ? _GEN6836 : _GEN15546;
wire  _GEN15548 = io_x[14] ? _GEN6856 : _GEN15547;
wire  _GEN15549 = io_x[0] ? _GEN15548 : _GEN6845;
wire  _GEN15550 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15551 = io_x[41] ? _GEN6836 : _GEN15550;
wire  _GEN15552 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN15553 = io_x[14] ? _GEN15552 : _GEN15551;
wire  _GEN15554 = io_x[0] ? _GEN15553 : _GEN6845;
wire  _GEN15555 = io_x[76] ? _GEN15554 : _GEN15549;
wire  _GEN15556 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15557 = io_x[41] ? _GEN15556 : _GEN6836;
wire  _GEN15558 = io_x[14] ? _GEN6843 : _GEN15557;
wire  _GEN15559 = io_x[0] ? _GEN15558 : _GEN6858;
wire  _GEN15560 = io_x[76] ? _GEN6833 : _GEN15559;
wire  _GEN15561 = io_x[42] ? _GEN15560 : _GEN15555;
wire  _GEN15562 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15563 = io_x[41] ? _GEN6836 : _GEN15562;
wire  _GEN15564 = io_x[14] ? _GEN6843 : _GEN15563;
wire  _GEN15565 = io_x[0] ? _GEN6858 : _GEN15564;
wire  _GEN15566 = io_x[76] ? _GEN15565 : _GEN6833;
wire  _GEN15567 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN15568 = io_x[14] ? _GEN6843 : _GEN15567;
wire  _GEN15569 = io_x[0] ? _GEN15568 : _GEN6845;
wire  _GEN15570 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN15571 = io_x[2] ? _GEN6837 : _GEN15570;
wire  _GEN15572 = io_x[6] ? _GEN6850 : _GEN15571;
wire  _GEN15573 = io_x[41] ? _GEN15572 : _GEN6836;
wire  _GEN15574 = io_x[14] ? _GEN6856 : _GEN15573;
wire  _GEN15575 = io_x[0] ? _GEN6845 : _GEN15574;
wire  _GEN15576 = io_x[76] ? _GEN15575 : _GEN15569;
wire  _GEN15577 = io_x[42] ? _GEN15576 : _GEN15566;
wire  _GEN15578 = io_x[38] ? _GEN15577 : _GEN15561;
wire  _GEN15579 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15580 = io_x[6] ? _GEN15579 : _GEN6840;
wire  _GEN15581 = io_x[41] ? _GEN15580 : _GEN6836;
wire  _GEN15582 = io_x[14] ? _GEN15581 : _GEN6843;
wire  _GEN15583 = io_x[0] ? _GEN15582 : _GEN6845;
wire  _GEN15584 = io_x[76] ? _GEN6833 : _GEN15583;
wire  _GEN15585 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN15586 = io_x[14] ? _GEN15585 : _GEN6856;
wire  _GEN15587 = io_x[0] ? _GEN15586 : _GEN6845;
wire  _GEN15588 = io_x[76] ? _GEN6834 : _GEN15587;
wire  _GEN15589 = io_x[42] ? _GEN15588 : _GEN15584;
wire  _GEN15590 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15591 = io_x[0] ? _GEN15590 : _GEN6845;
wire  _GEN15592 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN15593 = io_x[0] ? _GEN6845 : _GEN15592;
wire  _GEN15594 = io_x[76] ? _GEN15593 : _GEN15591;
wire  _GEN15595 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15596 = io_x[6] ? _GEN6850 : _GEN15595;
wire  _GEN15597 = io_x[41] ? _GEN6836 : _GEN15596;
wire  _GEN15598 = io_x[14] ? _GEN15597 : _GEN6856;
wire  _GEN15599 = io_x[0] ? _GEN6845 : _GEN15598;
wire  _GEN15600 = io_x[76] ? _GEN15599 : _GEN6833;
wire  _GEN15601 = io_x[42] ? _GEN15600 : _GEN15594;
wire  _GEN15602 = io_x[38] ? _GEN15601 : _GEN15589;
wire  _GEN15603 = io_x[10] ? _GEN15602 : _GEN15578;
wire  _GEN15604 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15605 = io_x[6] ? _GEN15604 : _GEN6850;
wire  _GEN15606 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15607 = io_x[41] ? _GEN15606 : _GEN15605;
wire  _GEN15608 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15609 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15610 = io_x[41] ? _GEN15609 : _GEN15608;
wire  _GEN15611 = io_x[14] ? _GEN15610 : _GEN15607;
wire  _GEN15612 = io_x[0] ? _GEN15611 : _GEN6858;
wire  _GEN15613 = io_x[76] ? _GEN6834 : _GEN15612;
wire  _GEN15614 = io_x[42] ? _GEN6874 : _GEN15613;
wire  _GEN15615 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15616 = io_x[6] ? _GEN6840 : _GEN15615;
wire  _GEN15617 = io_x[41] ? _GEN6836 : _GEN15616;
wire  _GEN15618 = io_x[14] ? _GEN6843 : _GEN15617;
wire  _GEN15619 = io_x[0] ? _GEN6845 : _GEN15618;
wire  _GEN15620 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15621 = io_x[41] ? _GEN15620 : _GEN6836;
wire  _GEN15622 = io_x[14] ? _GEN6856 : _GEN15621;
wire  _GEN15623 = io_x[0] ? _GEN6845 : _GEN15622;
wire  _GEN15624 = io_x[76] ? _GEN15623 : _GEN15619;
wire  _GEN15625 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15626 = io_x[6] ? _GEN15625 : _GEN6840;
wire  _GEN15627 = io_x[41] ? _GEN15626 : _GEN6836;
wire  _GEN15628 = io_x[14] ? _GEN6843 : _GEN15627;
wire  _GEN15629 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15630 = io_x[41] ? _GEN6836 : _GEN15629;
wire  _GEN15631 = io_x[14] ? _GEN6843 : _GEN15630;
wire  _GEN15632 = io_x[0] ? _GEN15631 : _GEN15628;
wire  _GEN15633 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15634 = io_x[6] ? _GEN6850 : _GEN15633;
wire  _GEN15635 = io_x[41] ? _GEN6836 : _GEN15634;
wire  _GEN15636 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15637 = io_x[41] ? _GEN6836 : _GEN15636;
wire  _GEN15638 = io_x[14] ? _GEN15637 : _GEN15635;
wire  _GEN15639 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15640 = io_x[6] ? _GEN6840 : _GEN15639;
wire  _GEN15641 = io_x[41] ? _GEN6836 : _GEN15640;
wire  _GEN15642 = io_x[14] ? _GEN6843 : _GEN15641;
wire  _GEN15643 = io_x[0] ? _GEN15642 : _GEN15638;
wire  _GEN15644 = io_x[76] ? _GEN15643 : _GEN15632;
wire  _GEN15645 = io_x[42] ? _GEN15644 : _GEN15624;
wire  _GEN15646 = io_x[38] ? _GEN15645 : _GEN15614;
wire  _GEN15647 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15648 = io_x[6] ? _GEN15647 : _GEN6850;
wire  _GEN15649 = io_x[41] ? _GEN6836 : _GEN15648;
wire  _GEN15650 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15651 = io_x[6] ? _GEN6840 : _GEN15650;
wire  _GEN15652 = io_x[41] ? _GEN6836 : _GEN15651;
wire  _GEN15653 = io_x[14] ? _GEN15652 : _GEN15649;
wire  _GEN15654 = io_x[0] ? _GEN15653 : _GEN6845;
wire  _GEN15655 = io_x[76] ? _GEN6834 : _GEN15654;
wire  _GEN15656 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15657 = io_x[0] ? _GEN6845 : _GEN15656;
wire  _GEN15658 = io_x[76] ? _GEN6834 : _GEN15657;
wire  _GEN15659 = io_x[42] ? _GEN15658 : _GEN15655;
wire  _GEN15660 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15661 = io_x[0] ? _GEN6858 : _GEN15660;
wire  _GEN15662 = io_x[76] ? _GEN6833 : _GEN15661;
wire  _GEN15663 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15664 = io_x[6] ? _GEN15663 : _GEN6850;
wire  _GEN15665 = io_x[41] ? _GEN6836 : _GEN15664;
wire  _GEN15666 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15667 = io_x[6] ? _GEN6850 : _GEN15666;
wire  _GEN15668 = io_x[41] ? _GEN6836 : _GEN15667;
wire  _GEN15669 = io_x[14] ? _GEN15668 : _GEN15665;
wire  _GEN15670 = io_x[0] ? _GEN6845 : _GEN15669;
wire  _GEN15671 = io_x[76] ? _GEN15670 : _GEN6834;
wire  _GEN15672 = io_x[42] ? _GEN15671 : _GEN15662;
wire  _GEN15673 = io_x[38] ? _GEN15672 : _GEN15659;
wire  _GEN15674 = io_x[10] ? _GEN15673 : _GEN15646;
wire  _GEN15675 = io_x[71] ? _GEN15674 : _GEN15603;
wire  _GEN15676 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN15677 = io_x[2] ? _GEN6837 : _GEN15676;
wire  _GEN15678 = io_x[6] ? _GEN6850 : _GEN15677;
wire  _GEN15679 = io_x[41] ? _GEN6836 : _GEN15678;
wire  _GEN15680 = io_x[14] ? _GEN6843 : _GEN15679;
wire  _GEN15681 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15682 = io_x[41] ? _GEN6924 : _GEN15681;
wire  _GEN15683 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15684 = io_x[41] ? _GEN15683 : _GEN6836;
wire  _GEN15685 = io_x[14] ? _GEN15684 : _GEN15682;
wire  _GEN15686 = io_x[0] ? _GEN15685 : _GEN15680;
wire  _GEN15687 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15688 = io_x[6] ? _GEN15687 : _GEN6850;
wire  _GEN15689 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15690 = io_x[41] ? _GEN15689 : _GEN15688;
wire  _GEN15691 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15692 = io_x[41] ? _GEN15691 : _GEN6836;
wire  _GEN15693 = io_x[14] ? _GEN15692 : _GEN15690;
wire  _GEN15694 = io_x[0] ? _GEN15693 : _GEN6845;
wire  _GEN15695 = io_x[76] ? _GEN15694 : _GEN15686;
wire  _GEN15696 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15697 = io_x[6] ? _GEN6840 : _GEN15696;
wire  _GEN15698 = io_x[41] ? _GEN6836 : _GEN15697;
wire  _GEN15699 = io_x[14] ? _GEN6843 : _GEN15698;
wire  _GEN15700 = io_x[0] ? _GEN6845 : _GEN15699;
wire  _GEN15701 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN15702 = io_x[2] ? _GEN6837 : _GEN15701;
wire  _GEN15703 = io_x[6] ? _GEN6850 : _GEN15702;
wire  _GEN15704 = io_x[41] ? _GEN15703 : _GEN6836;
wire  _GEN15705 = io_x[14] ? _GEN6843 : _GEN15704;
wire  _GEN15706 = io_x[0] ? _GEN6845 : _GEN15705;
wire  _GEN15707 = io_x[76] ? _GEN15706 : _GEN15700;
wire  _GEN15708 = io_x[42] ? _GEN15707 : _GEN15695;
wire  _GEN15709 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15710 = io_x[6] ? _GEN15709 : _GEN6840;
wire  _GEN15711 = io_x[41] ? _GEN15710 : _GEN6836;
wire  _GEN15712 = io_x[14] ? _GEN15711 : _GEN6843;
wire  _GEN15713 = io_x[0] ? _GEN15712 : _GEN6845;
wire  _GEN15714 = io_x[76] ? _GEN15713 : _GEN6834;
wire  _GEN15715 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15716 = io_x[6] ? _GEN6850 : _GEN15715;
wire  _GEN15717 = io_x[41] ? _GEN15716 : _GEN6836;
wire  _GEN15718 = io_x[14] ? _GEN6843 : _GEN15717;
wire  _GEN15719 = io_x[0] ? _GEN6858 : _GEN15718;
wire  _GEN15720 = io_x[76] ? _GEN6834 : _GEN15719;
wire  _GEN15721 = io_x[42] ? _GEN15720 : _GEN15714;
wire  _GEN15722 = io_x[38] ? _GEN15721 : _GEN15708;
wire  _GEN15723 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15724 = io_x[0] ? _GEN15723 : _GEN6845;
wire  _GEN15725 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15726 = io_x[41] ? _GEN15725 : _GEN6836;
wire  _GEN15727 = io_x[14] ? _GEN6843 : _GEN15726;
wire  _GEN15728 = io_x[0] ? _GEN15727 : _GEN6845;
wire  _GEN15729 = io_x[76] ? _GEN15728 : _GEN15724;
wire  _GEN15730 = io_x[42] ? _GEN6874 : _GEN15729;
wire  _GEN15731 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15732 = io_x[0] ? _GEN6845 : _GEN15731;
wire  _GEN15733 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN15734 = io_x[0] ? _GEN15733 : _GEN6858;
wire  _GEN15735 = io_x[76] ? _GEN15734 : _GEN15732;
wire  _GEN15736 = io_x[42] ? _GEN6874 : _GEN15735;
wire  _GEN15737 = io_x[38] ? _GEN15736 : _GEN15730;
wire  _GEN15738 = io_x[10] ? _GEN15737 : _GEN15722;
wire  _GEN15739 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN15740 = io_x[0] ? _GEN15739 : _GEN6858;
wire  _GEN15741 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15742 = io_x[6] ? _GEN6850 : _GEN15741;
wire  _GEN15743 = io_x[41] ? _GEN15742 : _GEN6836;
wire  _GEN15744 = io_x[14] ? _GEN15743 : _GEN6856;
wire  _GEN15745 = io_x[0] ? _GEN15744 : _GEN6845;
wire  _GEN15746 = io_x[76] ? _GEN15745 : _GEN15740;
wire  _GEN15747 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15748 = io_x[6] ? _GEN6850 : _GEN15747;
wire  _GEN15749 = io_x[41] ? _GEN15748 : _GEN6836;
wire  _GEN15750 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15751 = io_x[6] ? _GEN6840 : _GEN15750;
wire  _GEN15752 = io_x[41] ? _GEN15751 : _GEN6836;
wire  _GEN15753 = io_x[14] ? _GEN15752 : _GEN15749;
wire  _GEN15754 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15755 = io_x[41] ? _GEN15754 : _GEN6836;
wire  _GEN15756 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN15757 = io_x[14] ? _GEN15756 : _GEN15755;
wire  _GEN15758 = io_x[0] ? _GEN15757 : _GEN15753;
wire  _GEN15759 = io_x[76] ? _GEN15758 : _GEN6833;
wire  _GEN15760 = io_x[42] ? _GEN15759 : _GEN15746;
wire  _GEN15761 = io_x[38] ? _GEN7036 : _GEN15760;
wire  _GEN15762 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN15763 = io_x[2] ? _GEN15762 : _GEN6837;
wire  _GEN15764 = io_x[6] ? _GEN15763 : _GEN6850;
wire  _GEN15765 = io_x[41] ? _GEN6836 : _GEN15764;
wire  _GEN15766 = io_x[14] ? _GEN15765 : _GEN6843;
wire  _GEN15767 = io_x[0] ? _GEN15766 : _GEN6845;
wire  _GEN15768 = io_x[76] ? _GEN6833 : _GEN15767;
wire  _GEN15769 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15770 = io_x[0] ? _GEN15769 : _GEN6845;
wire  _GEN15771 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15772 = io_x[6] ? _GEN6850 : _GEN15771;
wire  _GEN15773 = io_x[41] ? _GEN15772 : _GEN6836;
wire  _GEN15774 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15775 = io_x[6] ? _GEN6850 : _GEN15774;
wire  _GEN15776 = io_x[41] ? _GEN15775 : _GEN6836;
wire  _GEN15777 = io_x[14] ? _GEN15776 : _GEN15773;
wire  _GEN15778 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15779 = io_x[41] ? _GEN15778 : _GEN6836;
wire  _GEN15780 = io_x[14] ? _GEN15779 : _GEN6843;
wire  _GEN15781 = io_x[0] ? _GEN15780 : _GEN15777;
wire  _GEN15782 = io_x[76] ? _GEN15781 : _GEN15770;
wire  _GEN15783 = io_x[42] ? _GEN15782 : _GEN15768;
wire  _GEN15784 = io_x[38] ? _GEN7036 : _GEN15783;
wire  _GEN15785 = io_x[10] ? _GEN15784 : _GEN15761;
wire  _GEN15786 = io_x[71] ? _GEN15785 : _GEN15738;
wire  _GEN15787 = io_x[70] ? _GEN15786 : _GEN15675;
wire  _GEN15788 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15789 = io_x[41] ? _GEN6836 : _GEN15788;
wire  _GEN15790 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15791 = io_x[41] ? _GEN6836 : _GEN15790;
wire  _GEN15792 = io_x[14] ? _GEN15791 : _GEN15789;
wire  _GEN15793 = io_x[0] ? _GEN15792 : _GEN6845;
wire  _GEN15794 = io_x[76] ? _GEN6834 : _GEN15793;
wire  _GEN15795 = io_x[42] ? _GEN15794 : _GEN6863;
wire  _GEN15796 = io_x[38] ? _GEN6871 : _GEN15795;
wire  _GEN15797 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15798 = io_x[0] ? _GEN15797 : _GEN6845;
wire  _GEN15799 = io_x[76] ? _GEN6834 : _GEN15798;
wire  _GEN15800 = io_x[42] ? _GEN6874 : _GEN15799;
wire  _GEN15801 = io_x[38] ? _GEN15800 : _GEN6871;
wire  _GEN15802 = io_x[10] ? _GEN15801 : _GEN15796;
wire  _GEN15803 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN15804 = io_x[76] ? _GEN6834 : _GEN15803;
wire  _GEN15805 = io_x[42] ? _GEN6874 : _GEN15804;
wire  _GEN15806 = io_x[38] ? _GEN15805 : _GEN6871;
wire  _GEN15807 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15808 = io_x[0] ? _GEN6845 : _GEN15807;
wire  _GEN15809 = io_x[76] ? _GEN6834 : _GEN15808;
wire  _GEN15810 = io_x[42] ? _GEN6874 : _GEN15809;
wire  _GEN15811 = io_x[38] ? _GEN15810 : _GEN6871;
wire  _GEN15812 = io_x[10] ? _GEN15811 : _GEN15806;
wire  _GEN15813 = io_x[71] ? _GEN15812 : _GEN15802;
wire  _GEN15814 = io_x[70] ? _GEN8474 : _GEN15813;
wire  _GEN15815 = io_x[33] ? _GEN15814 : _GEN15787;
wire  _GEN15816 = io_x[21] ? _GEN15815 : _GEN15545;
wire  _GEN15817 = io_x[18] ? _GEN15816 : _GEN15399;
wire  _GEN15818 = io_x[20] ? _GEN15817 : _GEN15142;
wire  _GEN15819 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN15820 = io_x[2] ? _GEN6837 : _GEN15819;
wire  _GEN15821 = io_x[6] ? _GEN6850 : _GEN15820;
wire  _GEN15822 = io_x[41] ? _GEN6836 : _GEN15821;
wire  _GEN15823 = io_x[14] ? _GEN6843 : _GEN15822;
wire  _GEN15824 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15825 = io_x[6] ? _GEN6850 : _GEN15824;
wire  _GEN15826 = io_x[41] ? _GEN6836 : _GEN15825;
wire  _GEN15827 = io_x[14] ? _GEN6843 : _GEN15826;
wire  _GEN15828 = io_x[0] ? _GEN15827 : _GEN15823;
wire  _GEN15829 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN15830 = io_x[2] ? _GEN6837 : _GEN15829;
wire  _GEN15831 = io_x[6] ? _GEN6850 : _GEN15830;
wire  _GEN15832 = io_x[41] ? _GEN15831 : _GEN6836;
wire  _GEN15833 = io_x[14] ? _GEN6843 : _GEN15832;
wire  _GEN15834 = io_x[0] ? _GEN6845 : _GEN15833;
wire  _GEN15835 = io_x[76] ? _GEN15834 : _GEN15828;
wire  _GEN15836 = io_x[42] ? _GEN6863 : _GEN15835;
wire  _GEN15837 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15838 = io_x[0] ? _GEN6845 : _GEN15837;
wire  _GEN15839 = io_x[76] ? _GEN6834 : _GEN15838;
wire  _GEN15840 = io_x[42] ? _GEN6863 : _GEN15839;
wire  _GEN15841 = io_x[38] ? _GEN15840 : _GEN15836;
wire  _GEN15842 = io_x[10] ? _GEN7044 : _GEN15841;
wire  _GEN15843 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15844 = io_x[41] ? _GEN15843 : _GEN6836;
wire  _GEN15845 = io_x[14] ? _GEN6843 : _GEN15844;
wire  _GEN15846 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15847 = io_x[6] ? _GEN6850 : _GEN15846;
wire  _GEN15848 = io_x[41] ? _GEN6924 : _GEN15847;
wire  _GEN15849 = io_x[14] ? _GEN6843 : _GEN15848;
wire  _GEN15850 = io_x[0] ? _GEN15849 : _GEN15845;
wire  _GEN15851 = io_x[76] ? _GEN6834 : _GEN15850;
wire  _GEN15852 = io_x[42] ? _GEN6863 : _GEN15851;
wire  _GEN15853 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15854 = io_x[41] ? _GEN6836 : _GEN15853;
wire  _GEN15855 = io_x[14] ? _GEN6843 : _GEN15854;
wire  _GEN15856 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN15857 = io_x[14] ? _GEN6843 : _GEN15856;
wire  _GEN15858 = io_x[0] ? _GEN15857 : _GEN15855;
wire  _GEN15859 = io_x[76] ? _GEN6834 : _GEN15858;
wire  _GEN15860 = io_x[42] ? _GEN6874 : _GEN15859;
wire  _GEN15861 = io_x[38] ? _GEN15860 : _GEN15852;
wire  _GEN15862 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15863 = io_x[6] ? _GEN6850 : _GEN15862;
wire  _GEN15864 = io_x[41] ? _GEN15863 : _GEN6836;
wire  _GEN15865 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15866 = io_x[41] ? _GEN15865 : _GEN6836;
wire  _GEN15867 = io_x[14] ? _GEN15866 : _GEN15864;
wire  _GEN15868 = io_x[0] ? _GEN6845 : _GEN15867;
wire  _GEN15869 = io_x[76] ? _GEN6834 : _GEN15868;
wire  _GEN15870 = io_x[42] ? _GEN6874 : _GEN15869;
wire  _GEN15871 = io_x[38] ? _GEN6871 : _GEN15870;
wire  _GEN15872 = io_x[10] ? _GEN15871 : _GEN15861;
wire  _GEN15873 = io_x[71] ? _GEN15872 : _GEN15842;
wire  _GEN15874 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN15875 = io_x[2] ? _GEN6837 : _GEN15874;
wire  _GEN15876 = io_x[6] ? _GEN6850 : _GEN15875;
wire  _GEN15877 = io_x[41] ? _GEN15876 : _GEN6924;
wire  _GEN15878 = io_x[14] ? _GEN6843 : _GEN15877;
wire  _GEN15879 = io_x[0] ? _GEN6845 : _GEN15878;
wire  _GEN15880 = io_x[76] ? _GEN6834 : _GEN15879;
wire  _GEN15881 = io_x[42] ? _GEN6863 : _GEN15880;
wire  _GEN15882 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN15883 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15884 = io_x[6] ? _GEN6850 : _GEN15883;
wire  _GEN15885 = io_x[41] ? _GEN15884 : _GEN6836;
wire  _GEN15886 = io_x[14] ? _GEN6843 : _GEN15885;
wire  _GEN15887 = io_x[0] ? _GEN15886 : _GEN6858;
wire  _GEN15888 = io_x[76] ? _GEN6834 : _GEN15887;
wire  _GEN15889 = io_x[42] ? _GEN15888 : _GEN15882;
wire  _GEN15890 = io_x[38] ? _GEN15889 : _GEN15881;
wire  _GEN15891 = io_x[10] ? _GEN7044 : _GEN15890;
wire  _GEN15892 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN15893 = io_x[14] ? _GEN6843 : _GEN15892;
wire  _GEN15894 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15895 = io_x[6] ? _GEN6850 : _GEN15894;
wire  _GEN15896 = io_x[41] ? _GEN15895 : _GEN6836;
wire  _GEN15897 = io_x[14] ? _GEN6843 : _GEN15896;
wire  _GEN15898 = io_x[0] ? _GEN15897 : _GEN15893;
wire  _GEN15899 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN15900 = io_x[0] ? _GEN6845 : _GEN15899;
wire  _GEN15901 = io_x[76] ? _GEN15900 : _GEN15898;
wire  _GEN15902 = io_x[42] ? _GEN6863 : _GEN15901;
wire  _GEN15903 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN15904 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN15905 = io_x[42] ? _GEN15904 : _GEN15903;
wire  _GEN15906 = io_x[38] ? _GEN15905 : _GEN15902;
wire  _GEN15907 = io_x[10] ? _GEN7094 : _GEN15906;
wire  _GEN15908 = io_x[71] ? _GEN15907 : _GEN15891;
wire  _GEN15909 = io_x[70] ? _GEN15908 : _GEN15873;
wire  _GEN15910 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15911 = io_x[41] ? _GEN6836 : _GEN15910;
wire  _GEN15912 = io_x[14] ? _GEN6843 : _GEN15911;
wire  _GEN15913 = io_x[0] ? _GEN6845 : _GEN15912;
wire  _GEN15914 = io_x[76] ? _GEN6834 : _GEN15913;
wire  _GEN15915 = io_x[42] ? _GEN6874 : _GEN15914;
wire  _GEN15916 = io_x[38] ? _GEN7036 : _GEN15915;
wire  _GEN15917 = io_x[10] ? _GEN7094 : _GEN15916;
wire  _GEN15918 = io_x[71] ? _GEN7203 : _GEN15917;
wire  _GEN15919 = io_x[70] ? _GEN15918 : _GEN8474;
wire  _GEN15920 = io_x[33] ? _GEN15919 : _GEN15909;
wire  _GEN15921 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN15922 = io_x[10] ? _GEN7044 : _GEN15921;
wire  _GEN15923 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN15924 = io_x[42] ? _GEN6874 : _GEN15923;
wire  _GEN15925 = io_x[38] ? _GEN15924 : _GEN7036;
wire  _GEN15926 = io_x[10] ? _GEN7044 : _GEN15925;
wire  _GEN15927 = io_x[71] ? _GEN15926 : _GEN15922;
wire  _GEN15928 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN15929 = io_x[38] ? _GEN15928 : _GEN7036;
wire  _GEN15930 = io_x[10] ? _GEN7044 : _GEN15929;
wire  _GEN15931 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN15932 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN15933 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN15934 = io_x[76] ? _GEN6834 : _GEN15933;
wire  _GEN15935 = io_x[42] ? _GEN15934 : _GEN15932;
wire  _GEN15936 = io_x[38] ? _GEN15935 : _GEN15931;
wire  _GEN15937 = io_x[10] ? _GEN7044 : _GEN15936;
wire  _GEN15938 = io_x[71] ? _GEN15937 : _GEN15930;
wire  _GEN15939 = io_x[70] ? _GEN15938 : _GEN15927;
wire  _GEN15940 = io_x[33] ? _GEN12627 : _GEN15939;
wire  _GEN15941 = io_x[21] ? _GEN15940 : _GEN15920;
wire  _GEN15942 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN15943 = io_x[42] ? _GEN6863 : _GEN15942;
wire  _GEN15944 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN15945 = io_x[76] ? _GEN6834 : _GEN15944;
wire  _GEN15946 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15947 = io_x[6] ? _GEN6850 : _GEN15946;
wire  _GEN15948 = io_x[41] ? _GEN6836 : _GEN15947;
wire  _GEN15949 = io_x[14] ? _GEN6843 : _GEN15948;
wire  _GEN15950 = io_x[0] ? _GEN6845 : _GEN15949;
wire  _GEN15951 = io_x[76] ? _GEN6833 : _GEN15950;
wire  _GEN15952 = io_x[42] ? _GEN15951 : _GEN15945;
wire  _GEN15953 = io_x[38] ? _GEN15952 : _GEN15943;
wire  _GEN15954 = io_x[10] ? _GEN7044 : _GEN15953;
wire  _GEN15955 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN15956 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN15957 = io_x[41] ? _GEN15956 : _GEN6836;
wire  _GEN15958 = io_x[14] ? _GEN6856 : _GEN15957;
wire  _GEN15959 = io_x[0] ? _GEN15958 : _GEN15955;
wire  _GEN15960 = io_x[76] ? _GEN6834 : _GEN15959;
wire  _GEN15961 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15962 = io_x[41] ? _GEN6836 : _GEN15961;
wire  _GEN15963 = io_x[14] ? _GEN6856 : _GEN15962;
wire  _GEN15964 = io_x[0] ? _GEN6845 : _GEN15963;
wire  _GEN15965 = io_x[76] ? _GEN15964 : _GEN6833;
wire  _GEN15966 = io_x[42] ? _GEN15965 : _GEN15960;
wire  _GEN15967 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15968 = io_x[41] ? _GEN15967 : _GEN6836;
wire  _GEN15969 = io_x[14] ? _GEN6843 : _GEN15968;
wire  _GEN15970 = io_x[0] ? _GEN6845 : _GEN15969;
wire  _GEN15971 = io_x[76] ? _GEN6834 : _GEN15970;
wire  _GEN15972 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN15973 = io_x[42] ? _GEN15972 : _GEN15971;
wire  _GEN15974 = io_x[38] ? _GEN15973 : _GEN15966;
wire  _GEN15975 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN15976 = io_x[6] ? _GEN15975 : _GEN6850;
wire  _GEN15977 = io_x[41] ? _GEN6836 : _GEN15976;
wire  _GEN15978 = io_x[14] ? _GEN15977 : _GEN6843;
wire  _GEN15979 = io_x[0] ? _GEN6845 : _GEN15978;
wire  _GEN15980 = io_x[76] ? _GEN15979 : _GEN6834;
wire  _GEN15981 = io_x[42] ? _GEN15980 : _GEN6874;
wire  _GEN15982 = io_x[38] ? _GEN6871 : _GEN15981;
wire  _GEN15983 = io_x[10] ? _GEN15982 : _GEN15974;
wire  _GEN15984 = io_x[71] ? _GEN15983 : _GEN15954;
wire  _GEN15985 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN15986 = io_x[41] ? _GEN15985 : _GEN6836;
wire  _GEN15987 = io_x[14] ? _GEN6856 : _GEN15986;
wire  _GEN15988 = io_x[0] ? _GEN6858 : _GEN15987;
wire  _GEN15989 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN15990 = io_x[76] ? _GEN15989 : _GEN15988;
wire  _GEN15991 = io_x[42] ? _GEN6863 : _GEN15990;
wire  _GEN15992 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN15993 = io_x[6] ? _GEN6850 : _GEN15992;
wire  _GEN15994 = io_x[41] ? _GEN15993 : _GEN6836;
wire  _GEN15995 = io_x[14] ? _GEN6843 : _GEN15994;
wire  _GEN15996 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN15997 = io_x[14] ? _GEN6843 : _GEN15996;
wire  _GEN15998 = io_x[0] ? _GEN15997 : _GEN15995;
wire  _GEN15999 = io_x[76] ? _GEN6834 : _GEN15998;
wire  _GEN16000 = io_x[42] ? _GEN6863 : _GEN15999;
wire  _GEN16001 = io_x[38] ? _GEN16000 : _GEN15991;
wire  _GEN16002 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN16003 = io_x[10] ? _GEN16002 : _GEN16001;
wire  _GEN16004 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN16005 = io_x[42] ? _GEN6863 : _GEN16004;
wire  _GEN16006 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16007 = io_x[6] ? _GEN6850 : _GEN16006;
wire  _GEN16008 = io_x[41] ? _GEN6836 : _GEN16007;
wire  _GEN16009 = io_x[14] ? _GEN6843 : _GEN16008;
wire  _GEN16010 = io_x[0] ? _GEN16009 : _GEN6845;
wire  _GEN16011 = io_x[76] ? _GEN16010 : _GEN6834;
wire  _GEN16012 = io_x[42] ? _GEN6863 : _GEN16011;
wire  _GEN16013 = io_x[38] ? _GEN16012 : _GEN16005;
wire  _GEN16014 = io_x[10] ? _GEN7094 : _GEN16013;
wire  _GEN16015 = io_x[71] ? _GEN16014 : _GEN16003;
wire  _GEN16016 = io_x[70] ? _GEN16015 : _GEN15984;
wire  _GEN16017 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN16018 = io_x[76] ? _GEN6834 : _GEN16017;
wire  _GEN16019 = io_x[42] ? _GEN6874 : _GEN16018;
wire  _GEN16020 = io_x[38] ? _GEN16019 : _GEN6871;
wire  _GEN16021 = io_x[10] ? _GEN7044 : _GEN16020;
wire  _GEN16022 = io_x[71] ? _GEN7203 : _GEN16021;
wire  _GEN16023 = io_x[70] ? _GEN7020 : _GEN16022;
wire  _GEN16024 = io_x[33] ? _GEN16023 : _GEN16016;
wire  _GEN16025 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN16026 = io_x[76] ? _GEN6834 : _GEN16025;
wire  _GEN16027 = io_x[42] ? _GEN6874 : _GEN16026;
wire  _GEN16028 = io_x[38] ? _GEN16027 : _GEN6871;
wire  _GEN16029 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN16030 = io_x[0] ? _GEN16029 : _GEN6845;
wire  _GEN16031 = io_x[76] ? _GEN16030 : _GEN6834;
wire  _GEN16032 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16033 = io_x[0] ? _GEN16032 : _GEN6845;
wire  _GEN16034 = io_x[76] ? _GEN6834 : _GEN16033;
wire  _GEN16035 = io_x[42] ? _GEN16034 : _GEN16031;
wire  _GEN16036 = io_x[38] ? _GEN16035 : _GEN6871;
wire  _GEN16037 = io_x[10] ? _GEN16036 : _GEN16028;
wire  _GEN16038 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN16039 = io_x[2] ? _GEN16038 : _GEN6837;
wire  _GEN16040 = io_x[6] ? _GEN6840 : _GEN16039;
wire  _GEN16041 = io_x[41] ? _GEN16040 : _GEN6836;
wire  _GEN16042 = io_x[14] ? _GEN6843 : _GEN16041;
wire  _GEN16043 = io_x[0] ? _GEN16042 : _GEN6858;
wire  _GEN16044 = io_x[76] ? _GEN6834 : _GEN16043;
wire  _GEN16045 = io_x[42] ? _GEN6874 : _GEN16044;
wire  _GEN16046 = io_x[38] ? _GEN7036 : _GEN16045;
wire  _GEN16047 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16048 = io_x[41] ? _GEN16047 : _GEN6836;
wire  _GEN16049 = io_x[14] ? _GEN16048 : _GEN6843;
wire  _GEN16050 = io_x[0] ? _GEN16049 : _GEN6845;
wire  _GEN16051 = io_x[76] ? _GEN6834 : _GEN16050;
wire  _GEN16052 = io_x[42] ? _GEN6863 : _GEN16051;
wire  _GEN16053 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN16054 = io_x[42] ? _GEN6863 : _GEN16053;
wire  _GEN16055 = io_x[38] ? _GEN16054 : _GEN16052;
wire  _GEN16056 = io_x[10] ? _GEN16055 : _GEN16046;
wire  _GEN16057 = io_x[71] ? _GEN16056 : _GEN16037;
wire  _GEN16058 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN16059 = io_x[76] ? _GEN16058 : _GEN6834;
wire  _GEN16060 = io_x[42] ? _GEN6874 : _GEN16059;
wire  _GEN16061 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN16062 = io_x[14] ? _GEN6843 : _GEN16061;
wire  _GEN16063 = io_x[0] ? _GEN16062 : _GEN6845;
wire  _GEN16064 = io_x[76] ? _GEN6833 : _GEN16063;
wire  _GEN16065 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN16066 = io_x[76] ? _GEN6834 : _GEN16065;
wire  _GEN16067 = io_x[42] ? _GEN16066 : _GEN16064;
wire  _GEN16068 = io_x[38] ? _GEN16067 : _GEN16060;
wire  _GEN16069 = io_x[10] ? _GEN7044 : _GEN16068;
wire  _GEN16070 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN16071 = io_x[76] ? _GEN6834 : _GEN16070;
wire  _GEN16072 = io_x[42] ? _GEN16071 : _GEN6863;
wire  _GEN16073 = io_x[38] ? _GEN6871 : _GEN16072;
wire  _GEN16074 = io_x[10] ? _GEN7094 : _GEN16073;
wire  _GEN16075 = io_x[71] ? _GEN16074 : _GEN16069;
wire  _GEN16076 = io_x[70] ? _GEN16075 : _GEN16057;
wire  _GEN16077 = io_x[33] ? _GEN12627 : _GEN16076;
wire  _GEN16078 = io_x[21] ? _GEN16077 : _GEN16024;
wire  _GEN16079 = io_x[18] ? _GEN16078 : _GEN15941;
wire  _GEN16080 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16081 = io_x[41] ? _GEN6836 : _GEN16080;
wire  _GEN16082 = io_x[14] ? _GEN6843 : _GEN16081;
wire  _GEN16083 = io_x[0] ? _GEN16082 : _GEN6845;
wire  _GEN16084 = io_x[76] ? _GEN6833 : _GEN16083;
wire  _GEN16085 = io_x[42] ? _GEN6874 : _GEN16084;
wire  _GEN16086 = io_x[38] ? _GEN6871 : _GEN16085;
wire  _GEN16087 = io_x[10] ? _GEN7044 : _GEN16086;
wire  _GEN16088 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN16089 = io_x[76] ? _GEN6833 : _GEN16088;
wire  _GEN16090 = io_x[42] ? _GEN6863 : _GEN16089;
wire  _GEN16091 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16092 = io_x[41] ? _GEN6836 : _GEN16091;
wire  _GEN16093 = io_x[14] ? _GEN6843 : _GEN16092;
wire  _GEN16094 = io_x[0] ? _GEN16093 : _GEN6845;
wire  _GEN16095 = io_x[76] ? _GEN6833 : _GEN16094;
wire  _GEN16096 = io_x[42] ? _GEN6874 : _GEN16095;
wire  _GEN16097 = io_x[38] ? _GEN16096 : _GEN16090;
wire  _GEN16098 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16099 = io_x[6] ? _GEN16098 : _GEN6850;
wire  _GEN16100 = io_x[41] ? _GEN16099 : _GEN6836;
wire  _GEN16101 = io_x[14] ? _GEN16100 : _GEN6843;
wire  _GEN16102 = io_x[0] ? _GEN6845 : _GEN16101;
wire  _GEN16103 = io_x[76] ? _GEN6834 : _GEN16102;
wire  _GEN16104 = io_x[42] ? _GEN16103 : _GEN6874;
wire  _GEN16105 = io_x[38] ? _GEN16104 : _GEN6871;
wire  _GEN16106 = io_x[10] ? _GEN16105 : _GEN16097;
wire  _GEN16107 = io_x[71] ? _GEN16106 : _GEN16087;
wire  _GEN16108 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16109 = io_x[41] ? _GEN6836 : _GEN16108;
wire  _GEN16110 = io_x[14] ? _GEN6843 : _GEN16109;
wire  _GEN16111 = io_x[0] ? _GEN16110 : _GEN6845;
wire  _GEN16112 = io_x[76] ? _GEN16111 : _GEN6834;
wire  _GEN16113 = io_x[42] ? _GEN6874 : _GEN16112;
wire  _GEN16114 = io_x[38] ? _GEN16113 : _GEN6871;
wire  _GEN16115 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16116 = io_x[0] ? _GEN6845 : _GEN16115;
wire  _GEN16117 = io_x[76] ? _GEN6834 : _GEN16116;
wire  _GEN16118 = io_x[42] ? _GEN6874 : _GEN16117;
wire  _GEN16119 = io_x[38] ? _GEN6871 : _GEN16118;
wire  _GEN16120 = io_x[10] ? _GEN16119 : _GEN16114;
wire  _GEN16121 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN16122 = io_x[14] ? _GEN6843 : _GEN16121;
wire  _GEN16123 = io_x[0] ? _GEN6845 : _GEN16122;
wire  _GEN16124 = io_x[76] ? _GEN6833 : _GEN16123;
wire  _GEN16125 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16126 = io_x[41] ? _GEN6836 : _GEN16125;
wire  _GEN16127 = io_x[14] ? _GEN16126 : _GEN6843;
wire  _GEN16128 = io_x[0] ? _GEN16127 : _GEN6845;
wire  _GEN16129 = io_x[76] ? _GEN6834 : _GEN16128;
wire  _GEN16130 = io_x[42] ? _GEN16129 : _GEN16124;
wire  _GEN16131 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16132 = io_x[41] ? _GEN6836 : _GEN16131;
wire  _GEN16133 = io_x[14] ? _GEN6843 : _GEN16132;
wire  _GEN16134 = io_x[0] ? _GEN16133 : _GEN6845;
wire  _GEN16135 = io_x[76] ? _GEN6834 : _GEN16134;
wire  _GEN16136 = io_x[42] ? _GEN6863 : _GEN16135;
wire  _GEN16137 = io_x[38] ? _GEN16136 : _GEN16130;
wire  _GEN16138 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16139 = io_x[0] ? _GEN16138 : _GEN6845;
wire  _GEN16140 = io_x[76] ? _GEN6834 : _GEN16139;
wire  _GEN16141 = io_x[42] ? _GEN16140 : _GEN6874;
wire  _GEN16142 = io_x[38] ? _GEN6871 : _GEN16141;
wire  _GEN16143 = io_x[10] ? _GEN16142 : _GEN16137;
wire  _GEN16144 = io_x[71] ? _GEN16143 : _GEN16120;
wire  _GEN16145 = io_x[70] ? _GEN16144 : _GEN16107;
wire  _GEN16146 = io_x[70] ? _GEN7020 : _GEN8474;
wire  _GEN16147 = io_x[33] ? _GEN16146 : _GEN16145;
wire  _GEN16148 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16149 = io_x[41] ? _GEN6836 : _GEN16148;
wire  _GEN16150 = io_x[14] ? _GEN6843 : _GEN16149;
wire  _GEN16151 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16152 = io_x[41] ? _GEN6836 : _GEN16151;
wire  _GEN16153 = io_x[14] ? _GEN6843 : _GEN16152;
wire  _GEN16154 = io_x[0] ? _GEN16153 : _GEN16150;
wire  _GEN16155 = io_x[76] ? _GEN6834 : _GEN16154;
wire  _GEN16156 = io_x[42] ? _GEN6863 : _GEN16155;
wire  _GEN16157 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16158 = io_x[41] ? _GEN16157 : _GEN6836;
wire  _GEN16159 = io_x[14] ? _GEN6843 : _GEN16158;
wire  _GEN16160 = io_x[0] ? _GEN6845 : _GEN16159;
wire  _GEN16161 = io_x[76] ? _GEN6834 : _GEN16160;
wire  _GEN16162 = io_x[42] ? _GEN6874 : _GEN16161;
wire  _GEN16163 = io_x[38] ? _GEN16162 : _GEN16156;
wire  _GEN16164 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16165 = io_x[0] ? _GEN16164 : _GEN6845;
wire  _GEN16166 = io_x[76] ? _GEN6834 : _GEN16165;
wire  _GEN16167 = io_x[42] ? _GEN16166 : _GEN6874;
wire  _GEN16168 = io_x[38] ? _GEN16167 : _GEN6871;
wire  _GEN16169 = io_x[10] ? _GEN16168 : _GEN16163;
wire  _GEN16170 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN16171 = io_x[76] ? _GEN6834 : _GEN16170;
wire  _GEN16172 = io_x[42] ? _GEN6863 : _GEN16171;
wire  _GEN16173 = io_x[38] ? _GEN6871 : _GEN16172;
wire  _GEN16174 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN16175 = io_x[0] ? _GEN16174 : _GEN6845;
wire  _GEN16176 = io_x[76] ? _GEN6834 : _GEN16175;
wire  _GEN16177 = io_x[42] ? _GEN6874 : _GEN16176;
wire  _GEN16178 = io_x[38] ? _GEN16177 : _GEN7036;
wire  _GEN16179 = io_x[10] ? _GEN16178 : _GEN16173;
wire  _GEN16180 = io_x[71] ? _GEN16179 : _GEN16169;
wire  _GEN16181 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN16182 = io_x[42] ? _GEN6874 : _GEN16181;
wire  _GEN16183 = io_x[38] ? _GEN6871 : _GEN16182;
wire  _GEN16184 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16185 = io_x[0] ? _GEN16184 : _GEN6845;
wire  _GEN16186 = io_x[76] ? _GEN6834 : _GEN16185;
wire  _GEN16187 = io_x[42] ? _GEN16186 : _GEN6874;
wire  _GEN16188 = io_x[38] ? _GEN6871 : _GEN16187;
wire  _GEN16189 = io_x[10] ? _GEN16188 : _GEN16183;
wire  _GEN16190 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN16191 = io_x[0] ? _GEN6845 : _GEN16190;
wire  _GEN16192 = io_x[76] ? _GEN6834 : _GEN16191;
wire  _GEN16193 = io_x[42] ? _GEN16192 : _GEN6863;
wire  _GEN16194 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16195 = io_x[41] ? _GEN6836 : _GEN16194;
wire  _GEN16196 = io_x[14] ? _GEN6843 : _GEN16195;
wire  _GEN16197 = io_x[0] ? _GEN16196 : _GEN6858;
wire  _GEN16198 = io_x[76] ? _GEN6834 : _GEN16197;
wire  _GEN16199 = io_x[42] ? _GEN6863 : _GEN16198;
wire  _GEN16200 = io_x[38] ? _GEN16199 : _GEN16193;
wire  _GEN16201 = io_x[10] ? _GEN7044 : _GEN16200;
wire  _GEN16202 = io_x[71] ? _GEN16201 : _GEN16189;
wire  _GEN16203 = io_x[70] ? _GEN16202 : _GEN16180;
wire  _GEN16204 = io_x[33] ? _GEN12627 : _GEN16203;
wire  _GEN16205 = io_x[21] ? _GEN16204 : _GEN16147;
wire  _GEN16206 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16207 = io_x[41] ? _GEN6836 : _GEN16206;
wire  _GEN16208 = io_x[14] ? _GEN6843 : _GEN16207;
wire  _GEN16209 = io_x[0] ? _GEN6845 : _GEN16208;
wire  _GEN16210 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN16211 = io_x[14] ? _GEN6856 : _GEN16210;
wire  _GEN16212 = io_x[0] ? _GEN6845 : _GEN16211;
wire  _GEN16213 = io_x[76] ? _GEN16212 : _GEN16209;
wire  _GEN16214 = io_x[42] ? _GEN6874 : _GEN16213;
wire  _GEN16215 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16216 = io_x[6] ? _GEN6850 : _GEN16215;
wire  _GEN16217 = io_x[41] ? _GEN16216 : _GEN6836;
wire  _GEN16218 = io_x[14] ? _GEN6843 : _GEN16217;
wire  _GEN16219 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16220 = io_x[41] ? _GEN16219 : _GEN6836;
wire  _GEN16221 = io_x[14] ? _GEN6843 : _GEN16220;
wire  _GEN16222 = io_x[0] ? _GEN16221 : _GEN16218;
wire  _GEN16223 = io_x[76] ? _GEN6834 : _GEN16222;
wire  _GEN16224 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16225 = io_x[6] ? _GEN6850 : _GEN16224;
wire  _GEN16226 = io_x[41] ? _GEN16225 : _GEN6836;
wire  _GEN16227 = io_x[14] ? _GEN6843 : _GEN16226;
wire  _GEN16228 = io_x[0] ? _GEN16227 : _GEN6845;
wire  _GEN16229 = io_x[76] ? _GEN16228 : _GEN6834;
wire  _GEN16230 = io_x[42] ? _GEN16229 : _GEN16223;
wire  _GEN16231 = io_x[38] ? _GEN16230 : _GEN16214;
wire  _GEN16232 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN16233 = io_x[42] ? _GEN6874 : _GEN16232;
wire  _GEN16234 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN16235 = io_x[38] ? _GEN16234 : _GEN16233;
wire  _GEN16236 = io_x[10] ? _GEN16235 : _GEN16231;
wire  _GEN16237 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN16238 = io_x[14] ? _GEN6843 : _GEN16237;
wire  _GEN16239 = io_x[0] ? _GEN16238 : _GEN6845;
wire  _GEN16240 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN16241 = io_x[76] ? _GEN16240 : _GEN16239;
wire  _GEN16242 = io_x[42] ? _GEN6874 : _GEN16241;
wire  _GEN16243 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16244 = io_x[41] ? _GEN6836 : _GEN16243;
wire  _GEN16245 = io_x[14] ? _GEN6843 : _GEN16244;
wire  _GEN16246 = io_x[0] ? _GEN16245 : _GEN6858;
wire  _GEN16247 = io_x[76] ? _GEN6833 : _GEN16246;
wire  _GEN16248 = io_x[42] ? _GEN6863 : _GEN16247;
wire  _GEN16249 = io_x[38] ? _GEN16248 : _GEN16242;
wire  _GEN16250 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16251 = io_x[0] ? _GEN16250 : _GEN6845;
wire  _GEN16252 = io_x[76] ? _GEN6834 : _GEN16251;
wire  _GEN16253 = io_x[42] ? _GEN16252 : _GEN6874;
wire  _GEN16254 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16255 = io_x[0] ? _GEN16254 : _GEN6845;
wire  _GEN16256 = io_x[76] ? _GEN6834 : _GEN16255;
wire  _GEN16257 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16258 = io_x[41] ? _GEN16257 : _GEN6836;
wire  _GEN16259 = io_x[14] ? _GEN16258 : _GEN6843;
wire  _GEN16260 = io_x[0] ? _GEN16259 : _GEN6845;
wire  _GEN16261 = io_x[76] ? _GEN6834 : _GEN16260;
wire  _GEN16262 = io_x[42] ? _GEN16261 : _GEN16256;
wire  _GEN16263 = io_x[38] ? _GEN16262 : _GEN16253;
wire  _GEN16264 = io_x[10] ? _GEN16263 : _GEN16249;
wire  _GEN16265 = io_x[71] ? _GEN16264 : _GEN16236;
wire  _GEN16266 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN16267 = io_x[2] ? _GEN6837 : _GEN16266;
wire  _GEN16268 = io_x[6] ? _GEN6850 : _GEN16267;
wire  _GEN16269 = io_x[41] ? _GEN16268 : _GEN6836;
wire  _GEN16270 = io_x[14] ? _GEN6843 : _GEN16269;
wire  _GEN16271 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16272 = io_x[41] ? _GEN6836 : _GEN16271;
wire  _GEN16273 = io_x[14] ? _GEN6856 : _GEN16272;
wire  _GEN16274 = io_x[0] ? _GEN16273 : _GEN16270;
wire  _GEN16275 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN16276 = io_x[76] ? _GEN16275 : _GEN16274;
wire  _GEN16277 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN16278 = io_x[42] ? _GEN16277 : _GEN16276;
wire  _GEN16279 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN16280 = io_x[76] ? _GEN6834 : _GEN16279;
wire  _GEN16281 = io_x[42] ? _GEN16280 : _GEN6863;
wire  _GEN16282 = io_x[38] ? _GEN16281 : _GEN16278;
wire  _GEN16283 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN16284 = io_x[10] ? _GEN16283 : _GEN16282;
wire  _GEN16285 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN16286 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN16287 = io_x[2] ? _GEN16286 : _GEN6837;
wire  _GEN16288 = io_x[6] ? _GEN16287 : _GEN6850;
wire  _GEN16289 = io_x[41] ? _GEN6836 : _GEN16288;
wire  _GEN16290 = io_x[14] ? _GEN6856 : _GEN16289;
wire  _GEN16291 = io_x[0] ? _GEN6845 : _GEN16290;
wire  _GEN16292 = io_x[76] ? _GEN16291 : _GEN16285;
wire  _GEN16293 = io_x[42] ? _GEN6874 : _GEN16292;
wire  _GEN16294 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN16295 = io_x[2] ? _GEN6837 : _GEN16294;
wire  _GEN16296 = io_x[6] ? _GEN6850 : _GEN16295;
wire  _GEN16297 = io_x[41] ? _GEN6836 : _GEN16296;
wire  _GEN16298 = io_x[14] ? _GEN6843 : _GEN16297;
wire  _GEN16299 = io_x[0] ? _GEN6845 : _GEN16298;
wire  _GEN16300 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN16301 = io_x[0] ? _GEN16300 : _GEN6845;
wire  _GEN16302 = io_x[76] ? _GEN16301 : _GEN16299;
wire  _GEN16303 = io_x[42] ? _GEN6874 : _GEN16302;
wire  _GEN16304 = io_x[38] ? _GEN16303 : _GEN16293;
wire  _GEN16305 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN16306 = io_x[0] ? _GEN6845 : _GEN16305;
wire  _GEN16307 = io_x[76] ? _GEN16306 : _GEN6834;
wire  _GEN16308 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN16309 = io_x[0] ? _GEN6845 : _GEN16308;
wire  _GEN16310 = io_x[76] ? _GEN6834 : _GEN16309;
wire  _GEN16311 = io_x[42] ? _GEN16310 : _GEN16307;
wire  _GEN16312 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16313 = io_x[0] ? _GEN6845 : _GEN16312;
wire  _GEN16314 = io_x[76] ? _GEN6834 : _GEN16313;
wire  _GEN16315 = io_x[42] ? _GEN16314 : _GEN6874;
wire  _GEN16316 = io_x[38] ? _GEN16315 : _GEN16311;
wire  _GEN16317 = io_x[10] ? _GEN16316 : _GEN16304;
wire  _GEN16318 = io_x[71] ? _GEN16317 : _GEN16284;
wire  _GEN16319 = io_x[70] ? _GEN16318 : _GEN16265;
wire  _GEN16320 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16321 = io_x[6] ? _GEN6850 : _GEN16320;
wire  _GEN16322 = io_x[41] ? _GEN16321 : _GEN6836;
wire  _GEN16323 = io_x[14] ? _GEN6843 : _GEN16322;
wire  _GEN16324 = io_x[0] ? _GEN16323 : _GEN6845;
wire  _GEN16325 = io_x[76] ? _GEN6834 : _GEN16324;
wire  _GEN16326 = io_x[42] ? _GEN6874 : _GEN16325;
wire  _GEN16327 = io_x[38] ? _GEN16326 : _GEN6871;
wire  _GEN16328 = io_x[10] ? _GEN7094 : _GEN16327;
wire  _GEN16329 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16330 = io_x[41] ? _GEN16329 : _GEN6836;
wire  _GEN16331 = io_x[14] ? _GEN6843 : _GEN16330;
wire  _GEN16332 = io_x[0] ? _GEN16331 : _GEN6845;
wire  _GEN16333 = io_x[76] ? _GEN16332 : _GEN6834;
wire  _GEN16334 = io_x[42] ? _GEN6874 : _GEN16333;
wire  _GEN16335 = io_x[38] ? _GEN16334 : _GEN7036;
wire  _GEN16336 = io_x[10] ? _GEN7044 : _GEN16335;
wire  _GEN16337 = io_x[71] ? _GEN16336 : _GEN16328;
wire  _GEN16338 = io_x[70] ? _GEN16337 : _GEN8474;
wire  _GEN16339 = io_x[33] ? _GEN16338 : _GEN16319;
wire  _GEN16340 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN16341 = io_x[2] ? _GEN16340 : _GEN6837;
wire  _GEN16342 = io_x[6] ? _GEN6850 : _GEN16341;
wire  _GEN16343 = io_x[41] ? _GEN6836 : _GEN16342;
wire  _GEN16344 = io_x[14] ? _GEN6843 : _GEN16343;
wire  _GEN16345 = io_x[0] ? _GEN16344 : _GEN6858;
wire  _GEN16346 = io_x[76] ? _GEN6834 : _GEN16345;
wire  _GEN16347 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16348 = io_x[41] ? _GEN16347 : _GEN6836;
wire  _GEN16349 = io_x[14] ? _GEN6843 : _GEN16348;
wire  _GEN16350 = io_x[0] ? _GEN6845 : _GEN16349;
wire  _GEN16351 = io_x[76] ? _GEN16350 : _GEN6833;
wire  _GEN16352 = io_x[42] ? _GEN16351 : _GEN16346;
wire  _GEN16353 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16354 = io_x[6] ? _GEN6840 : _GEN16353;
wire  _GEN16355 = io_x[41] ? _GEN16354 : _GEN6924;
wire  _GEN16356 = io_x[14] ? _GEN6843 : _GEN16355;
wire  _GEN16357 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16358 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16359 = io_x[6] ? _GEN16358 : _GEN16357;
wire  _GEN16360 = io_x[41] ? _GEN16359 : _GEN6836;
wire  _GEN16361 = io_x[14] ? _GEN6843 : _GEN16360;
wire  _GEN16362 = io_x[0] ? _GEN16361 : _GEN16356;
wire  _GEN16363 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16364 = io_x[41] ? _GEN6836 : _GEN16363;
wire  _GEN16365 = io_x[14] ? _GEN6856 : _GEN16364;
wire  _GEN16366 = io_x[0] ? _GEN16365 : _GEN6845;
wire  _GEN16367 = io_x[76] ? _GEN16366 : _GEN16362;
wire  _GEN16368 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16369 = io_x[6] ? _GEN6840 : _GEN16368;
wire  _GEN16370 = io_x[41] ? _GEN6836 : _GEN16369;
wire  _GEN16371 = io_x[14] ? _GEN6843 : _GEN16370;
wire  _GEN16372 = io_x[0] ? _GEN6845 : _GEN16371;
wire  _GEN16373 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16374 = io_x[6] ? _GEN6840 : _GEN16373;
wire  _GEN16375 = io_x[41] ? _GEN16374 : _GEN6836;
wire  _GEN16376 = io_x[14] ? _GEN6843 : _GEN16375;
wire  _GEN16377 = io_x[0] ? _GEN16376 : _GEN6845;
wire  _GEN16378 = io_x[76] ? _GEN16377 : _GEN16372;
wire  _GEN16379 = io_x[42] ? _GEN16378 : _GEN16367;
wire  _GEN16380 = io_x[38] ? _GEN16379 : _GEN16352;
wire  _GEN16381 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16382 = io_x[41] ? _GEN16381 : _GEN6836;
wire  _GEN16383 = io_x[14] ? _GEN6843 : _GEN16382;
wire  _GEN16384 = io_x[0] ? _GEN16383 : _GEN6845;
wire  _GEN16385 = io_x[76] ? _GEN6834 : _GEN16384;
wire  _GEN16386 = io_x[42] ? _GEN6863 : _GEN16385;
wire  _GEN16387 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16388 = io_x[0] ? _GEN16387 : _GEN6845;
wire  _GEN16389 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16390 = io_x[41] ? _GEN6836 : _GEN16389;
wire  _GEN16391 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16392 = io_x[41] ? _GEN6836 : _GEN16391;
wire  _GEN16393 = io_x[14] ? _GEN16392 : _GEN16390;
wire  _GEN16394 = io_x[0] ? _GEN16393 : _GEN6845;
wire  _GEN16395 = io_x[76] ? _GEN16394 : _GEN16388;
wire  _GEN16396 = io_x[42] ? _GEN6874 : _GEN16395;
wire  _GEN16397 = io_x[38] ? _GEN16396 : _GEN16386;
wire  _GEN16398 = io_x[10] ? _GEN16397 : _GEN16380;
wire  _GEN16399 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16400 = io_x[41] ? _GEN6836 : _GEN16399;
wire  _GEN16401 = io_x[14] ? _GEN6843 : _GEN16400;
wire  _GEN16402 = io_x[0] ? _GEN16401 : _GEN6845;
wire  _GEN16403 = io_x[76] ? _GEN6834 : _GEN16402;
wire  _GEN16404 = io_x[42] ? _GEN6874 : _GEN16403;
wire  _GEN16405 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16406 = io_x[6] ? _GEN6840 : _GEN16405;
wire  _GEN16407 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16408 = io_x[41] ? _GEN16407 : _GEN16406;
wire  _GEN16409 = io_x[14] ? _GEN6843 : _GEN16408;
wire  _GEN16410 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16411 = io_x[41] ? _GEN6836 : _GEN16410;
wire  _GEN16412 = io_x[14] ? _GEN6843 : _GEN16411;
wire  _GEN16413 = io_x[0] ? _GEN16412 : _GEN16409;
wire  _GEN16414 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16415 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN16416 = io_x[14] ? _GEN6856 : _GEN16415;
wire  _GEN16417 = io_x[0] ? _GEN16416 : _GEN16414;
wire  _GEN16418 = io_x[76] ? _GEN16417 : _GEN16413;
wire  _GEN16419 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN16420 = io_x[0] ? _GEN16419 : _GEN6845;
wire  _GEN16421 = io_x[76] ? _GEN6833 : _GEN16420;
wire  _GEN16422 = io_x[42] ? _GEN16421 : _GEN16418;
wire  _GEN16423 = io_x[38] ? _GEN16422 : _GEN16404;
wire  _GEN16424 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16425 = io_x[6] ? _GEN16424 : _GEN6850;
wire  _GEN16426 = io_x[41] ? _GEN16425 : _GEN6836;
wire  _GEN16427 = io_x[14] ? _GEN6843 : _GEN16426;
wire  _GEN16428 = io_x[0] ? _GEN16427 : _GEN6845;
wire  _GEN16429 = io_x[76] ? _GEN6834 : _GEN16428;
wire  _GEN16430 = io_x[42] ? _GEN6863 : _GEN16429;
wire  _GEN16431 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN16432 = io_x[38] ? _GEN16431 : _GEN16430;
wire  _GEN16433 = io_x[10] ? _GEN16432 : _GEN16423;
wire  _GEN16434 = io_x[71] ? _GEN16433 : _GEN16398;
wire  _GEN16435 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN16436 = io_x[14] ? _GEN6843 : _GEN16435;
wire  _GEN16437 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16438 = io_x[6] ? _GEN6840 : _GEN16437;
wire  _GEN16439 = io_x[41] ? _GEN6836 : _GEN16438;
wire  _GEN16440 = io_x[14] ? _GEN6843 : _GEN16439;
wire  _GEN16441 = io_x[0] ? _GEN16440 : _GEN16436;
wire  _GEN16442 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN16443 = io_x[76] ? _GEN16442 : _GEN16441;
wire  _GEN16444 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN16445 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16446 = io_x[41] ? _GEN6836 : _GEN16445;
wire  _GEN16447 = io_x[14] ? _GEN6843 : _GEN16446;
wire  _GEN16448 = io_x[0] ? _GEN16447 : _GEN16444;
wire  _GEN16449 = io_x[76] ? _GEN6834 : _GEN16448;
wire  _GEN16450 = io_x[42] ? _GEN16449 : _GEN16443;
wire  _GEN16451 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN16452 = io_x[14] ? _GEN6843 : _GEN16451;
wire  _GEN16453 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16454 = io_x[41] ? _GEN16453 : _GEN6924;
wire  _GEN16455 = io_x[14] ? _GEN6843 : _GEN16454;
wire  _GEN16456 = io_x[0] ? _GEN16455 : _GEN16452;
wire  _GEN16457 = io_x[76] ? _GEN6834 : _GEN16456;
wire  _GEN16458 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16459 = io_x[41] ? _GEN16458 : _GEN6836;
wire  _GEN16460 = io_x[14] ? _GEN16459 : _GEN6843;
wire  _GEN16461 = io_x[0] ? _GEN16460 : _GEN6858;
wire  _GEN16462 = io_x[76] ? _GEN6834 : _GEN16461;
wire  _GEN16463 = io_x[42] ? _GEN16462 : _GEN16457;
wire  _GEN16464 = io_x[38] ? _GEN16463 : _GEN16450;
wire  _GEN16465 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16466 = io_x[6] ? _GEN6850 : _GEN16465;
wire  _GEN16467 = io_x[41] ? _GEN16466 : _GEN6836;
wire  _GEN16468 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16469 = io_x[6] ? _GEN16468 : _GEN6850;
wire  _GEN16470 = io_x[41] ? _GEN16469 : _GEN6836;
wire  _GEN16471 = io_x[14] ? _GEN16470 : _GEN16467;
wire  _GEN16472 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN16473 = io_x[0] ? _GEN16472 : _GEN16471;
wire  _GEN16474 = io_x[76] ? _GEN6834 : _GEN16473;
wire  _GEN16475 = io_x[42] ? _GEN6863 : _GEN16474;
wire  _GEN16476 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16477 = io_x[0] ? _GEN16476 : _GEN6845;
wire  _GEN16478 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16479 = io_x[0] ? _GEN16478 : _GEN6845;
wire  _GEN16480 = io_x[76] ? _GEN16479 : _GEN16477;
wire  _GEN16481 = io_x[42] ? _GEN16480 : _GEN6863;
wire  _GEN16482 = io_x[38] ? _GEN16481 : _GEN16475;
wire  _GEN16483 = io_x[10] ? _GEN16482 : _GEN16464;
wire  _GEN16484 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16485 = io_x[6] ? _GEN6850 : _GEN16484;
wire  _GEN16486 = io_x[41] ? _GEN6924 : _GEN16485;
wire  _GEN16487 = io_x[14] ? _GEN6843 : _GEN16486;
wire  _GEN16488 = io_x[0] ? _GEN16487 : _GEN6845;
wire  _GEN16489 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16490 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16491 = io_x[6] ? _GEN16490 : _GEN16489;
wire  _GEN16492 = io_x[41] ? _GEN16491 : _GEN6836;
wire  _GEN16493 = io_x[14] ? _GEN6856 : _GEN16492;
wire  _GEN16494 = io_x[0] ? _GEN16493 : _GEN6845;
wire  _GEN16495 = io_x[76] ? _GEN16494 : _GEN16488;
wire  _GEN16496 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN16497 = io_x[76] ? _GEN6834 : _GEN16496;
wire  _GEN16498 = io_x[42] ? _GEN16497 : _GEN16495;
wire  _GEN16499 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN16500 = io_x[2] ? _GEN6837 : _GEN16499;
wire  _GEN16501 = io_x[6] ? _GEN6850 : _GEN16500;
wire  _GEN16502 = io_x[41] ? _GEN6836 : _GEN16501;
wire  _GEN16503 = io_x[14] ? _GEN6843 : _GEN16502;
wire  _GEN16504 = io_x[0] ? _GEN6845 : _GEN16503;
wire  _GEN16505 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN16506 = io_x[14] ? _GEN6843 : _GEN16505;
wire  _GEN16507 = io_x[0] ? _GEN16506 : _GEN6845;
wire  _GEN16508 = io_x[76] ? _GEN16507 : _GEN16504;
wire  _GEN16509 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16510 = io_x[6] ? _GEN16509 : _GEN6850;
wire  _GEN16511 = io_x[41] ? _GEN16510 : _GEN6836;
wire  _GEN16512 = io_x[14] ? _GEN16511 : _GEN6843;
wire  _GEN16513 = io_x[0] ? _GEN16512 : _GEN6858;
wire  _GEN16514 = io_x[76] ? _GEN6834 : _GEN16513;
wire  _GEN16515 = io_x[42] ? _GEN16514 : _GEN16508;
wire  _GEN16516 = io_x[38] ? _GEN16515 : _GEN16498;
wire  _GEN16517 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN16518 = io_x[2] ? _GEN16517 : _GEN6837;
wire  _GEN16519 = io_x[6] ? _GEN16518 : _GEN6840;
wire  _GEN16520 = io_x[41] ? _GEN16519 : _GEN6836;
wire  _GEN16521 = io_x[14] ? _GEN16520 : _GEN6843;
wire  _GEN16522 = io_x[0] ? _GEN16521 : _GEN6858;
wire  _GEN16523 = io_x[76] ? _GEN16522 : _GEN6834;
wire  _GEN16524 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN16525 = io_x[14] ? _GEN16524 : _GEN6843;
wire  _GEN16526 = io_x[0] ? _GEN6845 : _GEN16525;
wire  _GEN16527 = io_x[76] ? _GEN6834 : _GEN16526;
wire  _GEN16528 = io_x[42] ? _GEN16527 : _GEN16523;
wire  _GEN16529 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16530 = io_x[0] ? _GEN16529 : _GEN6845;
wire  _GEN16531 = io_x[76] ? _GEN16530 : _GEN6834;
wire  _GEN16532 = io_x[42] ? _GEN6874 : _GEN16531;
wire  _GEN16533 = io_x[38] ? _GEN16532 : _GEN16528;
wire  _GEN16534 = io_x[10] ? _GEN16533 : _GEN16516;
wire  _GEN16535 = io_x[71] ? _GEN16534 : _GEN16483;
wire  _GEN16536 = io_x[70] ? _GEN16535 : _GEN16434;
wire  _GEN16537 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN16538 = io_x[76] ? _GEN6834 : _GEN16537;
wire  _GEN16539 = io_x[42] ? _GEN6874 : _GEN16538;
wire  _GEN16540 = io_x[38] ? _GEN16539 : _GEN6871;
wire  _GEN16541 = io_x[10] ? _GEN7094 : _GEN16540;
wire  _GEN16542 = io_x[71] ? _GEN7203 : _GEN16541;
wire  _GEN16543 = io_x[70] ? _GEN16542 : _GEN7020;
wire  _GEN16544 = io_x[33] ? _GEN16543 : _GEN16536;
wire  _GEN16545 = io_x[21] ? _GEN16544 : _GEN16339;
wire  _GEN16546 = io_x[18] ? _GEN16545 : _GEN16205;
wire  _GEN16547 = io_x[20] ? _GEN16546 : _GEN16079;
wire  _GEN16548 = io_x[45] ? _GEN16547 : _GEN15818;
wire  _GEN16549 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16550 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16551 = io_x[6] ? _GEN16550 : _GEN16549;
wire  _GEN16552 = io_x[41] ? _GEN6836 : _GEN16551;
wire  _GEN16553 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16554 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16555 = io_x[6] ? _GEN16554 : _GEN16553;
wire  _GEN16556 = io_x[41] ? _GEN6836 : _GEN16555;
wire  _GEN16557 = io_x[14] ? _GEN16556 : _GEN16552;
wire  _GEN16558 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16559 = io_x[6] ? _GEN6840 : _GEN16558;
wire  _GEN16560 = io_x[41] ? _GEN6836 : _GEN16559;
wire  _GEN16561 = io_x[14] ? _GEN6856 : _GEN16560;
wire  _GEN16562 = io_x[0] ? _GEN16561 : _GEN16557;
wire  _GEN16563 = io_x[76] ? _GEN16562 : _GEN6834;
wire  _GEN16564 = io_x[42] ? _GEN16563 : _GEN6874;
wire  _GEN16565 = io_x[38] ? _GEN16564 : _GEN6871;
wire  _GEN16566 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16567 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16568 = io_x[6] ? _GEN16567 : _GEN16566;
wire  _GEN16569 = io_x[41] ? _GEN6836 : _GEN16568;
wire  _GEN16570 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16571 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16572 = io_x[6] ? _GEN16571 : _GEN16570;
wire  _GEN16573 = io_x[41] ? _GEN6836 : _GEN16572;
wire  _GEN16574 = io_x[14] ? _GEN16573 : _GEN16569;
wire  _GEN16575 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16576 = io_x[6] ? _GEN16575 : _GEN6840;
wire  _GEN16577 = io_x[41] ? _GEN6836 : _GEN16576;
wire  _GEN16578 = io_x[14] ? _GEN6843 : _GEN16577;
wire  _GEN16579 = io_x[0] ? _GEN16578 : _GEN16574;
wire  _GEN16580 = io_x[76] ? _GEN16579 : _GEN6834;
wire  _GEN16581 = io_x[42] ? _GEN16580 : _GEN6874;
wire  _GEN16582 = io_x[38] ? _GEN16581 : _GEN6871;
wire  _GEN16583 = io_x[10] ? _GEN16582 : _GEN16565;
wire  _GEN16584 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16585 = io_x[41] ? _GEN16584 : _GEN6836;
wire  _GEN16586 = io_x[14] ? _GEN16585 : _GEN6856;
wire  _GEN16587 = io_x[0] ? _GEN16586 : _GEN6845;
wire  _GEN16588 = io_x[76] ? _GEN16587 : _GEN6834;
wire  _GEN16589 = io_x[42] ? _GEN6874 : _GEN16588;
wire  _GEN16590 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16591 = io_x[0] ? _GEN6845 : _GEN16590;
wire  _GEN16592 = io_x[76] ? _GEN16591 : _GEN6834;
wire  _GEN16593 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16594 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16595 = io_x[6] ? _GEN16594 : _GEN16593;
wire  _GEN16596 = io_x[41] ? _GEN6836 : _GEN16595;
wire  _GEN16597 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16598 = io_x[6] ? _GEN6850 : _GEN16597;
wire  _GEN16599 = io_x[41] ? _GEN6836 : _GEN16598;
wire  _GEN16600 = io_x[14] ? _GEN16599 : _GEN16596;
wire  _GEN16601 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16602 = io_x[6] ? _GEN6840 : _GEN16601;
wire  _GEN16603 = io_x[41] ? _GEN6836 : _GEN16602;
wire  _GEN16604 = io_x[14] ? _GEN6856 : _GEN16603;
wire  _GEN16605 = io_x[0] ? _GEN16604 : _GEN16600;
wire  _GEN16606 = io_x[76] ? _GEN16605 : _GEN6834;
wire  _GEN16607 = io_x[42] ? _GEN16606 : _GEN16592;
wire  _GEN16608 = io_x[38] ? _GEN16607 : _GEN16589;
wire  _GEN16609 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16610 = io_x[41] ? _GEN16609 : _GEN6836;
wire  _GEN16611 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16612 = io_x[6] ? _GEN16611 : _GEN6850;
wire  _GEN16613 = io_x[41] ? _GEN16612 : _GEN6836;
wire  _GEN16614 = io_x[14] ? _GEN16613 : _GEN16610;
wire  _GEN16615 = io_x[0] ? _GEN16614 : _GEN6845;
wire  _GEN16616 = io_x[76] ? _GEN16615 : _GEN6834;
wire  _GEN16617 = io_x[42] ? _GEN6874 : _GEN16616;
wire  _GEN16618 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN16619 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16620 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16621 = io_x[6] ? _GEN16620 : _GEN16619;
wire  _GEN16622 = io_x[41] ? _GEN6836 : _GEN16621;
wire  _GEN16623 = io_x[14] ? _GEN6843 : _GEN16622;
wire  _GEN16624 = io_x[0] ? _GEN6858 : _GEN16623;
wire  _GEN16625 = io_x[76] ? _GEN16624 : _GEN6834;
wire  _GEN16626 = io_x[42] ? _GEN16625 : _GEN16618;
wire  _GEN16627 = io_x[38] ? _GEN16626 : _GEN16617;
wire  _GEN16628 = io_x[10] ? _GEN16627 : _GEN16608;
wire  _GEN16629 = io_x[71] ? _GEN16628 : _GEN16583;
wire  _GEN16630 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16631 = io_x[41] ? _GEN16630 : _GEN6836;
wire  _GEN16632 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16633 = io_x[41] ? _GEN16632 : _GEN6836;
wire  _GEN16634 = io_x[14] ? _GEN16633 : _GEN16631;
wire  _GEN16635 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16636 = io_x[41] ? _GEN16635 : _GEN6836;
wire  _GEN16637 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16638 = io_x[41] ? _GEN16637 : _GEN6836;
wire  _GEN16639 = io_x[14] ? _GEN16638 : _GEN16636;
wire  _GEN16640 = io_x[0] ? _GEN16639 : _GEN16634;
wire  _GEN16641 = io_x[76] ? _GEN16640 : _GEN6834;
wire  _GEN16642 = io_x[42] ? _GEN6874 : _GEN16641;
wire  _GEN16643 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16644 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16645 = io_x[6] ? _GEN16644 : _GEN16643;
wire  _GEN16646 = io_x[41] ? _GEN16645 : _GEN6836;
wire  _GEN16647 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16648 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16649 = io_x[6] ? _GEN16648 : _GEN16647;
wire  _GEN16650 = io_x[41] ? _GEN16649 : _GEN6836;
wire  _GEN16651 = io_x[14] ? _GEN16650 : _GEN16646;
wire  _GEN16652 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16653 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16654 = io_x[6] ? _GEN16653 : _GEN16652;
wire  _GEN16655 = io_x[41] ? _GEN16654 : _GEN6836;
wire  _GEN16656 = io_x[14] ? _GEN6856 : _GEN16655;
wire  _GEN16657 = io_x[0] ? _GEN16656 : _GEN16651;
wire  _GEN16658 = io_x[76] ? _GEN16657 : _GEN6834;
wire  _GEN16659 = io_x[42] ? _GEN6874 : _GEN16658;
wire  _GEN16660 = io_x[38] ? _GEN16659 : _GEN16642;
wire  _GEN16661 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16662 = io_x[41] ? _GEN16661 : _GEN6836;
wire  _GEN16663 = io_x[14] ? _GEN6856 : _GEN16662;
wire  _GEN16664 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16665 = io_x[41] ? _GEN16664 : _GEN6836;
wire  _GEN16666 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16667 = io_x[41] ? _GEN16666 : _GEN6836;
wire  _GEN16668 = io_x[14] ? _GEN16667 : _GEN16665;
wire  _GEN16669 = io_x[0] ? _GEN16668 : _GEN16663;
wire  _GEN16670 = io_x[76] ? _GEN16669 : _GEN6834;
wire  _GEN16671 = io_x[42] ? _GEN6874 : _GEN16670;
wire  _GEN16672 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16673 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16674 = io_x[6] ? _GEN16673 : _GEN16672;
wire  _GEN16675 = io_x[41] ? _GEN16674 : _GEN6836;
wire  _GEN16676 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16677 = io_x[6] ? _GEN16676 : _GEN6840;
wire  _GEN16678 = io_x[41] ? _GEN16677 : _GEN6836;
wire  _GEN16679 = io_x[14] ? _GEN16678 : _GEN16675;
wire  _GEN16680 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16681 = io_x[6] ? _GEN6850 : _GEN16680;
wire  _GEN16682 = io_x[41] ? _GEN16681 : _GEN6836;
wire  _GEN16683 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16684 = io_x[41] ? _GEN16683 : _GEN6836;
wire  _GEN16685 = io_x[14] ? _GEN16684 : _GEN16682;
wire  _GEN16686 = io_x[0] ? _GEN16685 : _GEN16679;
wire  _GEN16687 = io_x[76] ? _GEN16686 : _GEN6834;
wire  _GEN16688 = io_x[42] ? _GEN6863 : _GEN16687;
wire  _GEN16689 = io_x[38] ? _GEN16688 : _GEN16671;
wire  _GEN16690 = io_x[10] ? _GEN16689 : _GEN16660;
wire  _GEN16691 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16692 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16693 = io_x[6] ? _GEN16692 : _GEN16691;
wire  _GEN16694 = io_x[41] ? _GEN16693 : _GEN6836;
wire  _GEN16695 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16696 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16697 = io_x[6] ? _GEN16696 : _GEN16695;
wire  _GEN16698 = io_x[41] ? _GEN16697 : _GEN6836;
wire  _GEN16699 = io_x[14] ? _GEN16698 : _GEN16694;
wire  _GEN16700 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16701 = io_x[6] ? _GEN6840 : _GEN16700;
wire  _GEN16702 = io_x[41] ? _GEN16701 : _GEN6836;
wire  _GEN16703 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16704 = io_x[41] ? _GEN16703 : _GEN6836;
wire  _GEN16705 = io_x[14] ? _GEN16704 : _GEN16702;
wire  _GEN16706 = io_x[0] ? _GEN16705 : _GEN16699;
wire  _GEN16707 = io_x[76] ? _GEN16706 : _GEN6833;
wire  _GEN16708 = io_x[42] ? _GEN16707 : _GEN6874;
wire  _GEN16709 = io_x[38] ? _GEN6871 : _GEN16708;
wire  _GEN16710 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16711 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16712 = io_x[6] ? _GEN16711 : _GEN16710;
wire  _GEN16713 = io_x[41] ? _GEN16712 : _GEN6836;
wire  _GEN16714 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16715 = io_x[6] ? _GEN6840 : _GEN16714;
wire  _GEN16716 = io_x[41] ? _GEN16715 : _GEN6836;
wire  _GEN16717 = io_x[14] ? _GEN16716 : _GEN16713;
wire  _GEN16718 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16719 = io_x[41] ? _GEN16718 : _GEN6836;
wire  _GEN16720 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16721 = io_x[41] ? _GEN16720 : _GEN6836;
wire  _GEN16722 = io_x[14] ? _GEN16721 : _GEN16719;
wire  _GEN16723 = io_x[0] ? _GEN16722 : _GEN16717;
wire  _GEN16724 = io_x[76] ? _GEN16723 : _GEN6834;
wire  _GEN16725 = io_x[42] ? _GEN16724 : _GEN6874;
wire  _GEN16726 = io_x[38] ? _GEN6871 : _GEN16725;
wire  _GEN16727 = io_x[10] ? _GEN16726 : _GEN16709;
wire  _GEN16728 = io_x[71] ? _GEN16727 : _GEN16690;
wire  _GEN16729 = io_x[70] ? _GEN16728 : _GEN16629;
wire  _GEN16730 = io_x[33] ? _GEN12627 : _GEN16729;
wire  _GEN16731 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16732 = io_x[6] ? _GEN16731 : _GEN6840;
wire  _GEN16733 = io_x[41] ? _GEN6836 : _GEN16732;
wire  _GEN16734 = io_x[14] ? _GEN6843 : _GEN16733;
wire  _GEN16735 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16736 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16737 = io_x[6] ? _GEN16736 : _GEN16735;
wire  _GEN16738 = io_x[41] ? _GEN6836 : _GEN16737;
wire  _GEN16739 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16740 = io_x[6] ? _GEN6850 : _GEN16739;
wire  _GEN16741 = io_x[41] ? _GEN6836 : _GEN16740;
wire  _GEN16742 = io_x[14] ? _GEN16741 : _GEN16738;
wire  _GEN16743 = io_x[0] ? _GEN16742 : _GEN16734;
wire  _GEN16744 = io_x[76] ? _GEN16743 : _GEN6834;
wire  _GEN16745 = io_x[42] ? _GEN16744 : _GEN6863;
wire  _GEN16746 = io_x[38] ? _GEN16745 : _GEN7036;
wire  _GEN16747 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16748 = io_x[6] ? _GEN6840 : _GEN16747;
wire  _GEN16749 = io_x[41] ? _GEN6836 : _GEN16748;
wire  _GEN16750 = io_x[14] ? _GEN6843 : _GEN16749;
wire  _GEN16751 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16752 = io_x[6] ? _GEN6850 : _GEN16751;
wire  _GEN16753 = io_x[41] ? _GEN6836 : _GEN16752;
wire  _GEN16754 = io_x[14] ? _GEN6856 : _GEN16753;
wire  _GEN16755 = io_x[0] ? _GEN16754 : _GEN16750;
wire  _GEN16756 = io_x[76] ? _GEN16755 : _GEN6834;
wire  _GEN16757 = io_x[42] ? _GEN16756 : _GEN6874;
wire  _GEN16758 = io_x[38] ? _GEN16757 : _GEN6871;
wire  _GEN16759 = io_x[10] ? _GEN16758 : _GEN16746;
wire  _GEN16760 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16761 = io_x[6] ? _GEN6850 : _GEN16760;
wire  _GEN16762 = io_x[41] ? _GEN6836 : _GEN16761;
wire  _GEN16763 = io_x[14] ? _GEN6856 : _GEN16762;
wire  _GEN16764 = io_x[0] ? _GEN16763 : _GEN6858;
wire  _GEN16765 = io_x[76] ? _GEN16764 : _GEN6834;
wire  _GEN16766 = io_x[42] ? _GEN16765 : _GEN6874;
wire  _GEN16767 = io_x[38] ? _GEN16766 : _GEN6871;
wire  _GEN16768 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16769 = io_x[41] ? _GEN16768 : _GEN6836;
wire  _GEN16770 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16771 = io_x[41] ? _GEN16770 : _GEN6836;
wire  _GEN16772 = io_x[14] ? _GEN16771 : _GEN16769;
wire  _GEN16773 = io_x[0] ? _GEN16772 : _GEN6845;
wire  _GEN16774 = io_x[76] ? _GEN6833 : _GEN16773;
wire  _GEN16775 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN16776 = io_x[76] ? _GEN16775 : _GEN6834;
wire  _GEN16777 = io_x[42] ? _GEN16776 : _GEN16774;
wire  _GEN16778 = io_x[38] ? _GEN16777 : _GEN6871;
wire  _GEN16779 = io_x[10] ? _GEN16778 : _GEN16767;
wire  _GEN16780 = io_x[71] ? _GEN16779 : _GEN16759;
wire  _GEN16781 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16782 = io_x[41] ? _GEN16781 : _GEN6924;
wire  _GEN16783 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16784 = io_x[41] ? _GEN16783 : _GEN6836;
wire  _GEN16785 = io_x[14] ? _GEN16784 : _GEN16782;
wire  _GEN16786 = io_x[0] ? _GEN16785 : _GEN6845;
wire  _GEN16787 = io_x[76] ? _GEN16786 : _GEN6834;
wire  _GEN16788 = io_x[42] ? _GEN6874 : _GEN16787;
wire  _GEN16789 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16790 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16791 = io_x[6] ? _GEN16790 : _GEN16789;
wire  _GEN16792 = io_x[41] ? _GEN16791 : _GEN6836;
wire  _GEN16793 = io_x[14] ? _GEN6856 : _GEN16792;
wire  _GEN16794 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN16795 = io_x[0] ? _GEN16794 : _GEN16793;
wire  _GEN16796 = io_x[76] ? _GEN16795 : _GEN6834;
wire  _GEN16797 = io_x[42] ? _GEN6874 : _GEN16796;
wire  _GEN16798 = io_x[38] ? _GEN16797 : _GEN16788;
wire  _GEN16799 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16800 = io_x[41] ? _GEN16799 : _GEN6836;
wire  _GEN16801 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16802 = io_x[41] ? _GEN16801 : _GEN6836;
wire  _GEN16803 = io_x[14] ? _GEN16802 : _GEN16800;
wire  _GEN16804 = io_x[0] ? _GEN16803 : _GEN6845;
wire  _GEN16805 = io_x[76] ? _GEN16804 : _GEN6834;
wire  _GEN16806 = io_x[42] ? _GEN6874 : _GEN16805;
wire  _GEN16807 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16808 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16809 = io_x[6] ? _GEN16808 : _GEN16807;
wire  _GEN16810 = io_x[41] ? _GEN16809 : _GEN6836;
wire  _GEN16811 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16812 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16813 = io_x[6] ? _GEN16812 : _GEN16811;
wire  _GEN16814 = io_x[41] ? _GEN16813 : _GEN6836;
wire  _GEN16815 = io_x[14] ? _GEN16814 : _GEN16810;
wire  _GEN16816 = io_x[0] ? _GEN6858 : _GEN16815;
wire  _GEN16817 = io_x[76] ? _GEN16816 : _GEN6834;
wire  _GEN16818 = io_x[42] ? _GEN6874 : _GEN16817;
wire  _GEN16819 = io_x[38] ? _GEN16818 : _GEN16806;
wire  _GEN16820 = io_x[10] ? _GEN16819 : _GEN16798;
wire  _GEN16821 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16822 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16823 = io_x[6] ? _GEN16822 : _GEN16821;
wire  _GEN16824 = io_x[41] ? _GEN16823 : _GEN6836;
wire  _GEN16825 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16826 = io_x[6] ? _GEN6850 : _GEN16825;
wire  _GEN16827 = io_x[41] ? _GEN16826 : _GEN6836;
wire  _GEN16828 = io_x[14] ? _GEN16827 : _GEN16824;
wire  _GEN16829 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16830 = io_x[6] ? _GEN6840 : _GEN16829;
wire  _GEN16831 = io_x[41] ? _GEN16830 : _GEN6836;
wire  _GEN16832 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16833 = io_x[6] ? _GEN6850 : _GEN16832;
wire  _GEN16834 = io_x[41] ? _GEN16833 : _GEN6836;
wire  _GEN16835 = io_x[14] ? _GEN16834 : _GEN16831;
wire  _GEN16836 = io_x[0] ? _GEN16835 : _GEN16828;
wire  _GEN16837 = io_x[76] ? _GEN16836 : _GEN6834;
wire  _GEN16838 = io_x[42] ? _GEN16837 : _GEN6874;
wire  _GEN16839 = io_x[38] ? _GEN6871 : _GEN16838;
wire  _GEN16840 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16841 = io_x[6] ? _GEN6840 : _GEN16840;
wire  _GEN16842 = io_x[41] ? _GEN16841 : _GEN6836;
wire  _GEN16843 = io_x[14] ? _GEN6856 : _GEN16842;
wire  _GEN16844 = io_x[0] ? _GEN6858 : _GEN16843;
wire  _GEN16845 = io_x[76] ? _GEN16844 : _GEN6834;
wire  _GEN16846 = io_x[42] ? _GEN16845 : _GEN6874;
wire  _GEN16847 = io_x[38] ? _GEN6871 : _GEN16846;
wire  _GEN16848 = io_x[10] ? _GEN16847 : _GEN16839;
wire  _GEN16849 = io_x[71] ? _GEN16848 : _GEN16820;
wire  _GEN16850 = io_x[70] ? _GEN16849 : _GEN16780;
wire  _GEN16851 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN16852 = io_x[0] ? _GEN16851 : _GEN6845;
wire  _GEN16853 = io_x[76] ? _GEN6834 : _GEN16852;
wire  _GEN16854 = io_x[42] ? _GEN6874 : _GEN16853;
wire  _GEN16855 = io_x[38] ? _GEN16854 : _GEN6871;
wire  _GEN16856 = io_x[10] ? _GEN16855 : _GEN7044;
wire  _GEN16857 = io_x[71] ? _GEN7196 : _GEN16856;
wire  _GEN16858 = io_x[70] ? _GEN8474 : _GEN16857;
wire  _GEN16859 = io_x[33] ? _GEN16858 : _GEN16850;
wire  _GEN16860 = io_x[21] ? _GEN16859 : _GEN16730;
wire  _GEN16861 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN16862 = io_x[0] ? _GEN16861 : _GEN6845;
wire  _GEN16863 = io_x[76] ? _GEN16862 : _GEN6834;
wire  _GEN16864 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16865 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16866 = io_x[6] ? _GEN16865 : _GEN16864;
wire  _GEN16867 = io_x[41] ? _GEN6836 : _GEN16866;
wire  _GEN16868 = io_x[14] ? _GEN6856 : _GEN16867;
wire  _GEN16869 = io_x[0] ? _GEN6858 : _GEN16868;
wire  _GEN16870 = io_x[76] ? _GEN16869 : _GEN6834;
wire  _GEN16871 = io_x[42] ? _GEN16870 : _GEN16863;
wire  _GEN16872 = io_x[38] ? _GEN16871 : _GEN7036;
wire  _GEN16873 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16874 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16875 = io_x[6] ? _GEN16874 : _GEN16873;
wire  _GEN16876 = io_x[41] ? _GEN6836 : _GEN16875;
wire  _GEN16877 = io_x[14] ? _GEN6843 : _GEN16876;
wire  _GEN16878 = io_x[0] ? _GEN6845 : _GEN16877;
wire  _GEN16879 = io_x[76] ? _GEN16878 : _GEN6834;
wire  _GEN16880 = io_x[42] ? _GEN16879 : _GEN6874;
wire  _GEN16881 = io_x[38] ? _GEN16880 : _GEN7036;
wire  _GEN16882 = io_x[10] ? _GEN16881 : _GEN16872;
wire  _GEN16883 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN16884 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16885 = io_x[41] ? _GEN6836 : _GEN16884;
wire  _GEN16886 = io_x[14] ? _GEN16885 : _GEN6856;
wire  _GEN16887 = io_x[0] ? _GEN6845 : _GEN16886;
wire  _GEN16888 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16889 = io_x[6] ? _GEN6850 : _GEN16888;
wire  _GEN16890 = io_x[41] ? _GEN16889 : _GEN6836;
wire  _GEN16891 = io_x[14] ? _GEN6843 : _GEN16890;
wire  _GEN16892 = io_x[0] ? _GEN6845 : _GEN16891;
wire  _GEN16893 = io_x[76] ? _GEN16892 : _GEN16887;
wire  _GEN16894 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16895 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16896 = io_x[6] ? _GEN16895 : _GEN16894;
wire  _GEN16897 = io_x[41] ? _GEN6836 : _GEN16896;
wire  _GEN16898 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16899 = io_x[6] ? _GEN6850 : _GEN16898;
wire  _GEN16900 = io_x[41] ? _GEN6836 : _GEN16899;
wire  _GEN16901 = io_x[14] ? _GEN16900 : _GEN16897;
wire  _GEN16902 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16903 = io_x[6] ? _GEN6850 : _GEN16902;
wire  _GEN16904 = io_x[41] ? _GEN6836 : _GEN16903;
wire  _GEN16905 = io_x[14] ? _GEN6843 : _GEN16904;
wire  _GEN16906 = io_x[0] ? _GEN16905 : _GEN16901;
wire  _GEN16907 = io_x[76] ? _GEN16906 : _GEN6834;
wire  _GEN16908 = io_x[42] ? _GEN16907 : _GEN16893;
wire  _GEN16909 = io_x[38] ? _GEN16908 : _GEN16883;
wire  _GEN16910 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16911 = io_x[41] ? _GEN6836 : _GEN16910;
wire  _GEN16912 = io_x[14] ? _GEN16911 : _GEN6843;
wire  _GEN16913 = io_x[0] ? _GEN6858 : _GEN16912;
wire  _GEN16914 = io_x[76] ? _GEN6833 : _GEN16913;
wire  _GEN16915 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16916 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16917 = io_x[6] ? _GEN16916 : _GEN16915;
wire  _GEN16918 = io_x[41] ? _GEN6836 : _GEN16917;
wire  _GEN16919 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16920 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16921 = io_x[6] ? _GEN16920 : _GEN16919;
wire  _GEN16922 = io_x[41] ? _GEN6836 : _GEN16921;
wire  _GEN16923 = io_x[14] ? _GEN16922 : _GEN16918;
wire  _GEN16924 = io_x[0] ? _GEN6845 : _GEN16923;
wire  _GEN16925 = io_x[76] ? _GEN16924 : _GEN6834;
wire  _GEN16926 = io_x[42] ? _GEN16925 : _GEN16914;
wire  _GEN16927 = io_x[38] ? _GEN16926 : _GEN7036;
wire  _GEN16928 = io_x[10] ? _GEN16927 : _GEN16909;
wire  _GEN16929 = io_x[71] ? _GEN16928 : _GEN16882;
wire  _GEN16930 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16931 = io_x[41] ? _GEN16930 : _GEN6836;
wire  _GEN16932 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16933 = io_x[41] ? _GEN16932 : _GEN6836;
wire  _GEN16934 = io_x[14] ? _GEN16933 : _GEN16931;
wire  _GEN16935 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16936 = io_x[41] ? _GEN16935 : _GEN6836;
wire  _GEN16937 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16938 = io_x[41] ? _GEN16937 : _GEN6836;
wire  _GEN16939 = io_x[14] ? _GEN16938 : _GEN16936;
wire  _GEN16940 = io_x[0] ? _GEN16939 : _GEN16934;
wire  _GEN16941 = io_x[76] ? _GEN16940 : _GEN6834;
wire  _GEN16942 = io_x[42] ? _GEN6874 : _GEN16941;
wire  _GEN16943 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16944 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16945 = io_x[6] ? _GEN16944 : _GEN16943;
wire  _GEN16946 = io_x[41] ? _GEN16945 : _GEN6924;
wire  _GEN16947 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16948 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16949 = io_x[6] ? _GEN16948 : _GEN16947;
wire  _GEN16950 = io_x[41] ? _GEN16949 : _GEN6836;
wire  _GEN16951 = io_x[14] ? _GEN16950 : _GEN16946;
wire  _GEN16952 = io_x[0] ? _GEN16951 : _GEN6845;
wire  _GEN16953 = io_x[76] ? _GEN16952 : _GEN6834;
wire  _GEN16954 = io_x[42] ? _GEN6863 : _GEN16953;
wire  _GEN16955 = io_x[38] ? _GEN16954 : _GEN16942;
wire  _GEN16956 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16957 = io_x[41] ? _GEN16956 : _GEN6836;
wire  _GEN16958 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16959 = io_x[41] ? _GEN16958 : _GEN6836;
wire  _GEN16960 = io_x[14] ? _GEN16959 : _GEN16957;
wire  _GEN16961 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16962 = io_x[41] ? _GEN16961 : _GEN6836;
wire  _GEN16963 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16964 = io_x[41] ? _GEN16963 : _GEN6836;
wire  _GEN16965 = io_x[14] ? _GEN16964 : _GEN16962;
wire  _GEN16966 = io_x[0] ? _GEN16965 : _GEN16960;
wire  _GEN16967 = io_x[76] ? _GEN16966 : _GEN6834;
wire  _GEN16968 = io_x[42] ? _GEN6874 : _GEN16967;
wire  _GEN16969 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN16970 = io_x[41] ? _GEN16969 : _GEN6836;
wire  _GEN16971 = io_x[14] ? _GEN6856 : _GEN16970;
wire  _GEN16972 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16973 = io_x[41] ? _GEN16972 : _GEN6836;
wire  _GEN16974 = io_x[14] ? _GEN16973 : _GEN6856;
wire  _GEN16975 = io_x[0] ? _GEN16974 : _GEN16971;
wire  _GEN16976 = io_x[76] ? _GEN16975 : _GEN6834;
wire  _GEN16977 = io_x[42] ? _GEN6874 : _GEN16976;
wire  _GEN16978 = io_x[38] ? _GEN16977 : _GEN16968;
wire  _GEN16979 = io_x[10] ? _GEN16978 : _GEN16955;
wire  _GEN16980 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN16981 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16982 = io_x[6] ? _GEN16981 : _GEN16980;
wire  _GEN16983 = io_x[41] ? _GEN16982 : _GEN6836;
wire  _GEN16984 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16985 = io_x[6] ? _GEN6850 : _GEN16984;
wire  _GEN16986 = io_x[41] ? _GEN16985 : _GEN6836;
wire  _GEN16987 = io_x[14] ? _GEN16986 : _GEN16983;
wire  _GEN16988 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN16989 = io_x[41] ? _GEN16988 : _GEN6836;
wire  _GEN16990 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16991 = io_x[6] ? _GEN6850 : _GEN16990;
wire  _GEN16992 = io_x[41] ? _GEN16991 : _GEN6836;
wire  _GEN16993 = io_x[14] ? _GEN16992 : _GEN16989;
wire  _GEN16994 = io_x[0] ? _GEN16993 : _GEN16987;
wire  _GEN16995 = io_x[76] ? _GEN16994 : _GEN6834;
wire  _GEN16996 = io_x[42] ? _GEN16995 : _GEN6874;
wire  _GEN16997 = io_x[38] ? _GEN7036 : _GEN16996;
wire  _GEN16998 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN16999 = io_x[6] ? _GEN6840 : _GEN16998;
wire  _GEN17000 = io_x[41] ? _GEN16999 : _GEN6836;
wire  _GEN17001 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17002 = io_x[41] ? _GEN17001 : _GEN6836;
wire  _GEN17003 = io_x[14] ? _GEN17002 : _GEN17000;
wire  _GEN17004 = io_x[0] ? _GEN6845 : _GEN17003;
wire  _GEN17005 = io_x[76] ? _GEN17004 : _GEN6834;
wire  _GEN17006 = io_x[42] ? _GEN17005 : _GEN6863;
wire  _GEN17007 = io_x[38] ? _GEN6871 : _GEN17006;
wire  _GEN17008 = io_x[10] ? _GEN17007 : _GEN16997;
wire  _GEN17009 = io_x[71] ? _GEN17008 : _GEN16979;
wire  _GEN17010 = io_x[70] ? _GEN17009 : _GEN16929;
wire  _GEN17011 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN17012 = io_x[71] ? _GEN17011 : _GEN7196;
wire  _GEN17013 = io_x[70] ? _GEN8474 : _GEN17012;
wire  _GEN17014 = io_x[33] ? _GEN17013 : _GEN17010;
wire  _GEN17015 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17016 = io_x[41] ? _GEN6836 : _GEN17015;
wire  _GEN17017 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17018 = io_x[6] ? _GEN17017 : _GEN6850;
wire  _GEN17019 = io_x[41] ? _GEN6836 : _GEN17018;
wire  _GEN17020 = io_x[14] ? _GEN17019 : _GEN17016;
wire  _GEN17021 = io_x[0] ? _GEN17020 : _GEN6845;
wire  _GEN17022 = io_x[76] ? _GEN17021 : _GEN6834;
wire  _GEN17023 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN17024 = io_x[0] ? _GEN17023 : _GEN6858;
wire  _GEN17025 = io_x[76] ? _GEN17024 : _GEN6834;
wire  _GEN17026 = io_x[42] ? _GEN17025 : _GEN17022;
wire  _GEN17027 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17028 = io_x[41] ? _GEN6924 : _GEN17027;
wire  _GEN17029 = io_x[14] ? _GEN17028 : _GEN6843;
wire  _GEN17030 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17031 = io_x[41] ? _GEN17030 : _GEN6836;
wire  _GEN17032 = io_x[14] ? _GEN17031 : _GEN6856;
wire  _GEN17033 = io_x[0] ? _GEN17032 : _GEN17029;
wire  _GEN17034 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN17035 = io_x[0] ? _GEN6845 : _GEN17034;
wire  _GEN17036 = io_x[76] ? _GEN17035 : _GEN17033;
wire  _GEN17037 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN17038 = io_x[76] ? _GEN6834 : _GEN17037;
wire  _GEN17039 = io_x[42] ? _GEN17038 : _GEN17036;
wire  _GEN17040 = io_x[38] ? _GEN17039 : _GEN17026;
wire  _GEN17041 = io_x[10] ? _GEN17040 : _GEN7094;
wire  _GEN17042 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN17043 = io_x[0] ? _GEN6845 : _GEN17042;
wire  _GEN17044 = io_x[76] ? _GEN6834 : _GEN17043;
wire  _GEN17045 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN17046 = io_x[0] ? _GEN6845 : _GEN17045;
wire  _GEN17047 = io_x[76] ? _GEN6834 : _GEN17046;
wire  _GEN17048 = io_x[42] ? _GEN17047 : _GEN17044;
wire  _GEN17049 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17050 = io_x[41] ? _GEN17049 : _GEN6836;
wire  _GEN17051 = io_x[14] ? _GEN17050 : _GEN6856;
wire  _GEN17052 = io_x[0] ? _GEN6845 : _GEN17051;
wire  _GEN17053 = io_x[76] ? _GEN6834 : _GEN17052;
wire  _GEN17054 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17055 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17056 = io_x[6] ? _GEN17055 : _GEN17054;
wire  _GEN17057 = io_x[41] ? _GEN6836 : _GEN17056;
wire  _GEN17058 = io_x[14] ? _GEN6856 : _GEN17057;
wire  _GEN17059 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17060 = io_x[41] ? _GEN6836 : _GEN17059;
wire  _GEN17061 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17062 = io_x[6] ? _GEN6850 : _GEN17061;
wire  _GEN17063 = io_x[41] ? _GEN6836 : _GEN17062;
wire  _GEN17064 = io_x[14] ? _GEN17063 : _GEN17060;
wire  _GEN17065 = io_x[0] ? _GEN17064 : _GEN17058;
wire  _GEN17066 = io_x[76] ? _GEN17065 : _GEN6834;
wire  _GEN17067 = io_x[42] ? _GEN17066 : _GEN17053;
wire  _GEN17068 = io_x[38] ? _GEN17067 : _GEN17048;
wire  _GEN17069 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17070 = io_x[41] ? _GEN17069 : _GEN6924;
wire  _GEN17071 = io_x[14] ? _GEN17070 : _GEN6856;
wire  _GEN17072 = io_x[0] ? _GEN17071 : _GEN6858;
wire  _GEN17073 = io_x[76] ? _GEN6834 : _GEN17072;
wire  _GEN17074 = io_x[42] ? _GEN6863 : _GEN17073;
wire  _GEN17075 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17076 = io_x[41] ? _GEN6836 : _GEN17075;
wire  _GEN17077 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN17078 = io_x[14] ? _GEN17077 : _GEN17076;
wire  _GEN17079 = io_x[0] ? _GEN6845 : _GEN17078;
wire  _GEN17080 = io_x[76] ? _GEN6834 : _GEN17079;
wire  _GEN17081 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17082 = io_x[6] ? _GEN6850 : _GEN17081;
wire  _GEN17083 = io_x[41] ? _GEN6836 : _GEN17082;
wire  _GEN17084 = io_x[14] ? _GEN6843 : _GEN17083;
wire  _GEN17085 = io_x[0] ? _GEN6845 : _GEN17084;
wire  _GEN17086 = io_x[76] ? _GEN17085 : _GEN6833;
wire  _GEN17087 = io_x[42] ? _GEN17086 : _GEN17080;
wire  _GEN17088 = io_x[38] ? _GEN17087 : _GEN17074;
wire  _GEN17089 = io_x[10] ? _GEN17088 : _GEN17068;
wire  _GEN17090 = io_x[71] ? _GEN17089 : _GEN17041;
wire  _GEN17091 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17092 = io_x[41] ? _GEN17091 : _GEN6836;
wire  _GEN17093 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17094 = io_x[41] ? _GEN17093 : _GEN6836;
wire  _GEN17095 = io_x[14] ? _GEN17094 : _GEN17092;
wire  _GEN17096 = io_x[0] ? _GEN6858 : _GEN17095;
wire  _GEN17097 = io_x[76] ? _GEN17096 : _GEN6833;
wire  _GEN17098 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN17099 = io_x[42] ? _GEN17098 : _GEN17097;
wire  _GEN17100 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN17101 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17102 = io_x[6] ? _GEN6850 : _GEN17101;
wire  _GEN17103 = io_x[41] ? _GEN17102 : _GEN6836;
wire  _GEN17104 = io_x[14] ? _GEN6843 : _GEN17103;
wire  _GEN17105 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17106 = io_x[0] ? _GEN17105 : _GEN17104;
wire  _GEN17107 = io_x[76] ? _GEN17106 : _GEN17100;
wire  _GEN17108 = io_x[42] ? _GEN6874 : _GEN17107;
wire  _GEN17109 = io_x[38] ? _GEN17108 : _GEN17099;
wire  _GEN17110 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17111 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17112 = io_x[6] ? _GEN17111 : _GEN6840;
wire  _GEN17113 = io_x[41] ? _GEN17112 : _GEN17110;
wire  _GEN17114 = io_x[14] ? _GEN17113 : _GEN6856;
wire  _GEN17115 = io_x[0] ? _GEN17114 : _GEN6858;
wire  _GEN17116 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17117 = io_x[41] ? _GEN6924 : _GEN17116;
wire  _GEN17118 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17119 = io_x[41] ? _GEN6836 : _GEN17118;
wire  _GEN17120 = io_x[14] ? _GEN17119 : _GEN17117;
wire  _GEN17121 = io_x[0] ? _GEN17120 : _GEN6845;
wire  _GEN17122 = io_x[76] ? _GEN17121 : _GEN17115;
wire  _GEN17123 = io_x[42] ? _GEN6874 : _GEN17122;
wire  _GEN17124 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17125 = io_x[41] ? _GEN6836 : _GEN17124;
wire  _GEN17126 = io_x[14] ? _GEN17125 : _GEN6843;
wire  _GEN17127 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17128 = io_x[41] ? _GEN17127 : _GEN6836;
wire  _GEN17129 = io_x[14] ? _GEN6843 : _GEN17128;
wire  _GEN17130 = io_x[0] ? _GEN17129 : _GEN17126;
wire  _GEN17131 = io_x[76] ? _GEN17130 : _GEN6834;
wire  _GEN17132 = io_x[42] ? _GEN6874 : _GEN17131;
wire  _GEN17133 = io_x[38] ? _GEN17132 : _GEN17123;
wire  _GEN17134 = io_x[10] ? _GEN17133 : _GEN17109;
wire  _GEN17135 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN17136 = io_x[76] ? _GEN6833 : _GEN17135;
wire  _GEN17137 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17138 = io_x[41] ? _GEN17137 : _GEN6836;
wire  _GEN17139 = io_x[14] ? _GEN6856 : _GEN17138;
wire  _GEN17140 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17141 = io_x[41] ? _GEN17140 : _GEN6836;
wire  _GEN17142 = io_x[14] ? _GEN6843 : _GEN17141;
wire  _GEN17143 = io_x[0] ? _GEN17142 : _GEN17139;
wire  _GEN17144 = io_x[76] ? _GEN17143 : _GEN6833;
wire  _GEN17145 = io_x[42] ? _GEN17144 : _GEN17136;
wire  _GEN17146 = io_x[38] ? _GEN6871 : _GEN17145;
wire  _GEN17147 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17148 = io_x[6] ? _GEN17147 : _GEN6850;
wire  _GEN17149 = io_x[41] ? _GEN6836 : _GEN17148;
wire  _GEN17150 = io_x[14] ? _GEN17149 : _GEN6843;
wire  _GEN17151 = io_x[0] ? _GEN17150 : _GEN6858;
wire  _GEN17152 = io_x[76] ? _GEN6833 : _GEN17151;
wire  _GEN17153 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17154 = io_x[6] ? _GEN17153 : _GEN6850;
wire  _GEN17155 = io_x[41] ? _GEN6836 : _GEN17154;
wire  _GEN17156 = io_x[14] ? _GEN6856 : _GEN17155;
wire  _GEN17157 = io_x[0] ? _GEN17156 : _GEN6845;
wire  _GEN17158 = io_x[76] ? _GEN6834 : _GEN17157;
wire  _GEN17159 = io_x[42] ? _GEN17158 : _GEN17152;
wire  _GEN17160 = io_x[38] ? _GEN7036 : _GEN17159;
wire  _GEN17161 = io_x[10] ? _GEN17160 : _GEN17146;
wire  _GEN17162 = io_x[71] ? _GEN17161 : _GEN17134;
wire  _GEN17163 = io_x[70] ? _GEN17162 : _GEN17090;
wire  _GEN17164 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17165 = io_x[41] ? _GEN6836 : _GEN17164;
wire  _GEN17166 = io_x[14] ? _GEN17165 : _GEN6856;
wire  _GEN17167 = io_x[0] ? _GEN17166 : _GEN6845;
wire  _GEN17168 = io_x[76] ? _GEN6834 : _GEN17167;
wire  _GEN17169 = io_x[42] ? _GEN17168 : _GEN6874;
wire  _GEN17170 = io_x[38] ? _GEN7036 : _GEN17169;
wire  _GEN17171 = io_x[10] ? _GEN17170 : _GEN7044;
wire  _GEN17172 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN17173 = io_x[76] ? _GEN6834 : _GEN17172;
wire  _GEN17174 = io_x[42] ? _GEN6874 : _GEN17173;
wire  _GEN17175 = io_x[38] ? _GEN17174 : _GEN6871;
wire  _GEN17176 = io_x[10] ? _GEN17175 : _GEN7094;
wire  _GEN17177 = io_x[71] ? _GEN17176 : _GEN17171;
wire  _GEN17178 = io_x[70] ? _GEN8474 : _GEN17177;
wire  _GEN17179 = io_x[33] ? _GEN17178 : _GEN17163;
wire  _GEN17180 = io_x[21] ? _GEN17179 : _GEN17014;
wire  _GEN17181 = io_x[18] ? _GEN17180 : _GEN16860;
wire  _GEN17182 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17183 = io_x[41] ? _GEN6836 : _GEN17182;
wire  _GEN17184 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17185 = io_x[41] ? _GEN6836 : _GEN17184;
wire  _GEN17186 = io_x[14] ? _GEN17185 : _GEN17183;
wire  _GEN17187 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN17188 = io_x[0] ? _GEN17187 : _GEN17186;
wire  _GEN17189 = io_x[76] ? _GEN17188 : _GEN6834;
wire  _GEN17190 = io_x[42] ? _GEN17189 : _GEN6874;
wire  _GEN17191 = io_x[38] ? _GEN17190 : _GEN6871;
wire  _GEN17192 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17193 = io_x[41] ? _GEN6836 : _GEN17192;
wire  _GEN17194 = io_x[14] ? _GEN17193 : _GEN6856;
wire  _GEN17195 = io_x[0] ? _GEN6845 : _GEN17194;
wire  _GEN17196 = io_x[76] ? _GEN17195 : _GEN6834;
wire  _GEN17197 = io_x[42] ? _GEN17196 : _GEN6874;
wire  _GEN17198 = io_x[38] ? _GEN17197 : _GEN6871;
wire  _GEN17199 = io_x[10] ? _GEN17198 : _GEN17191;
wire  _GEN17200 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17201 = io_x[6] ? _GEN17200 : _GEN6850;
wire  _GEN17202 = io_x[41] ? _GEN6836 : _GEN17201;
wire  _GEN17203 = io_x[14] ? _GEN6856 : _GEN17202;
wire  _GEN17204 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17205 = io_x[6] ? _GEN6850 : _GEN17204;
wire  _GEN17206 = io_x[41] ? _GEN6836 : _GEN17205;
wire  _GEN17207 = io_x[14] ? _GEN17206 : _GEN6856;
wire  _GEN17208 = io_x[0] ? _GEN17207 : _GEN17203;
wire  _GEN17209 = io_x[76] ? _GEN17208 : _GEN6834;
wire  _GEN17210 = io_x[42] ? _GEN17209 : _GEN6874;
wire  _GEN17211 = io_x[38] ? _GEN17210 : _GEN6871;
wire  _GEN17212 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17213 = io_x[41] ? _GEN17212 : _GEN6836;
wire  _GEN17214 = io_x[14] ? _GEN17213 : _GEN6843;
wire  _GEN17215 = io_x[0] ? _GEN17214 : _GEN6845;
wire  _GEN17216 = io_x[76] ? _GEN6834 : _GEN17215;
wire  _GEN17217 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17218 = io_x[41] ? _GEN6836 : _GEN17217;
wire  _GEN17219 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17220 = io_x[6] ? _GEN6840 : _GEN17219;
wire  _GEN17221 = io_x[41] ? _GEN6836 : _GEN17220;
wire  _GEN17222 = io_x[14] ? _GEN17221 : _GEN17218;
wire  _GEN17223 = io_x[0] ? _GEN6845 : _GEN17222;
wire  _GEN17224 = io_x[76] ? _GEN17223 : _GEN6834;
wire  _GEN17225 = io_x[42] ? _GEN17224 : _GEN17216;
wire  _GEN17226 = io_x[38] ? _GEN17225 : _GEN6871;
wire  _GEN17227 = io_x[10] ? _GEN17226 : _GEN17211;
wire  _GEN17228 = io_x[71] ? _GEN17227 : _GEN17199;
wire  _GEN17229 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17230 = io_x[41] ? _GEN17229 : _GEN6836;
wire  _GEN17231 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17232 = io_x[41] ? _GEN17231 : _GEN6836;
wire  _GEN17233 = io_x[14] ? _GEN17232 : _GEN17230;
wire  _GEN17234 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17235 = io_x[41] ? _GEN17234 : _GEN6836;
wire  _GEN17236 = io_x[14] ? _GEN6856 : _GEN17235;
wire  _GEN17237 = io_x[0] ? _GEN17236 : _GEN17233;
wire  _GEN17238 = io_x[76] ? _GEN17237 : _GEN6834;
wire  _GEN17239 = io_x[42] ? _GEN6874 : _GEN17238;
wire  _GEN17240 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17241 = io_x[6] ? _GEN6850 : _GEN17240;
wire  _GEN17242 = io_x[41] ? _GEN17241 : _GEN6836;
wire  _GEN17243 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17244 = io_x[6] ? _GEN6850 : _GEN17243;
wire  _GEN17245 = io_x[41] ? _GEN17244 : _GEN6836;
wire  _GEN17246 = io_x[14] ? _GEN17245 : _GEN17242;
wire  _GEN17247 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17248 = io_x[0] ? _GEN17247 : _GEN17246;
wire  _GEN17249 = io_x[76] ? _GEN17248 : _GEN6834;
wire  _GEN17250 = io_x[42] ? _GEN6874 : _GEN17249;
wire  _GEN17251 = io_x[38] ? _GEN17250 : _GEN17239;
wire  _GEN17252 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17253 = io_x[41] ? _GEN17252 : _GEN6836;
wire  _GEN17254 = io_x[14] ? _GEN6843 : _GEN17253;
wire  _GEN17255 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17256 = io_x[41] ? _GEN17255 : _GEN6836;
wire  _GEN17257 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN17258 = io_x[14] ? _GEN17257 : _GEN17256;
wire  _GEN17259 = io_x[0] ? _GEN17258 : _GEN17254;
wire  _GEN17260 = io_x[76] ? _GEN17259 : _GEN6833;
wire  _GEN17261 = io_x[42] ? _GEN6874 : _GEN17260;
wire  _GEN17262 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17263 = io_x[41] ? _GEN17262 : _GEN6836;
wire  _GEN17264 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17265 = io_x[41] ? _GEN17264 : _GEN6836;
wire  _GEN17266 = io_x[14] ? _GEN17265 : _GEN17263;
wire  _GEN17267 = io_x[0] ? _GEN17266 : _GEN6845;
wire  _GEN17268 = io_x[76] ? _GEN17267 : _GEN6834;
wire  _GEN17269 = io_x[42] ? _GEN6863 : _GEN17268;
wire  _GEN17270 = io_x[38] ? _GEN17269 : _GEN17261;
wire  _GEN17271 = io_x[10] ? _GEN17270 : _GEN17251;
wire  _GEN17272 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17273 = io_x[41] ? _GEN17272 : _GEN6836;
wire  _GEN17274 = io_x[14] ? _GEN17273 : _GEN6843;
wire  _GEN17275 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17276 = io_x[6] ? _GEN6840 : _GEN17275;
wire  _GEN17277 = io_x[41] ? _GEN17276 : _GEN6836;
wire  _GEN17278 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17279 = io_x[6] ? _GEN6850 : _GEN17278;
wire  _GEN17280 = io_x[41] ? _GEN17279 : _GEN6836;
wire  _GEN17281 = io_x[14] ? _GEN17280 : _GEN17277;
wire  _GEN17282 = io_x[0] ? _GEN17281 : _GEN17274;
wire  _GEN17283 = io_x[76] ? _GEN17282 : _GEN6834;
wire  _GEN17284 = io_x[42] ? _GEN17283 : _GEN6874;
wire  _GEN17285 = io_x[38] ? _GEN6871 : _GEN17284;
wire  _GEN17286 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17287 = io_x[41] ? _GEN17286 : _GEN6836;
wire  _GEN17288 = io_x[14] ? _GEN17287 : _GEN6856;
wire  _GEN17289 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17290 = io_x[6] ? _GEN6850 : _GEN17289;
wire  _GEN17291 = io_x[41] ? _GEN17290 : _GEN6836;
wire  _GEN17292 = io_x[14] ? _GEN6843 : _GEN17291;
wire  _GEN17293 = io_x[0] ? _GEN17292 : _GEN17288;
wire  _GEN17294 = io_x[76] ? _GEN17293 : _GEN6834;
wire  _GEN17295 = io_x[42] ? _GEN17294 : _GEN6874;
wire  _GEN17296 = io_x[38] ? _GEN6871 : _GEN17295;
wire  _GEN17297 = io_x[10] ? _GEN17296 : _GEN17285;
wire  _GEN17298 = io_x[71] ? _GEN17297 : _GEN17271;
wire  _GEN17299 = io_x[70] ? _GEN17298 : _GEN17228;
wire  _GEN17300 = io_x[33] ? _GEN12641 : _GEN17299;
wire  _GEN17301 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17302 = io_x[41] ? _GEN17301 : _GEN6836;
wire  _GEN17303 = io_x[14] ? _GEN17302 : _GEN6843;
wire  _GEN17304 = io_x[0] ? _GEN17303 : _GEN6845;
wire  _GEN17305 = io_x[76] ? _GEN6834 : _GEN17304;
wire  _GEN17306 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN17307 = io_x[76] ? _GEN17306 : _GEN6833;
wire  _GEN17308 = io_x[42] ? _GEN17307 : _GEN17305;
wire  _GEN17309 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17310 = io_x[41] ? _GEN6924 : _GEN17309;
wire  _GEN17311 = io_x[14] ? _GEN6843 : _GEN17310;
wire  _GEN17312 = io_x[0] ? _GEN6858 : _GEN17311;
wire  _GEN17313 = io_x[76] ? _GEN17312 : _GEN6834;
wire  _GEN17314 = io_x[42] ? _GEN17313 : _GEN6863;
wire  _GEN17315 = io_x[38] ? _GEN17314 : _GEN17308;
wire  _GEN17316 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17317 = io_x[0] ? _GEN17316 : _GEN6845;
wire  _GEN17318 = io_x[76] ? _GEN6834 : _GEN17317;
wire  _GEN17319 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN17320 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17321 = io_x[41] ? _GEN17320 : _GEN6836;
wire  _GEN17322 = io_x[14] ? _GEN17321 : _GEN6843;
wire  _GEN17323 = io_x[0] ? _GEN17322 : _GEN6845;
wire  _GEN17324 = io_x[76] ? _GEN17323 : _GEN17319;
wire  _GEN17325 = io_x[42] ? _GEN17324 : _GEN17318;
wire  _GEN17326 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17327 = io_x[0] ? _GEN6845 : _GEN17326;
wire  _GEN17328 = io_x[76] ? _GEN17327 : _GEN6833;
wire  _GEN17329 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17330 = io_x[6] ? _GEN17329 : _GEN6840;
wire  _GEN17331 = io_x[41] ? _GEN6836 : _GEN17330;
wire  _GEN17332 = io_x[14] ? _GEN6843 : _GEN17331;
wire  _GEN17333 = io_x[0] ? _GEN17332 : _GEN6858;
wire  _GEN17334 = io_x[76] ? _GEN17333 : _GEN6833;
wire  _GEN17335 = io_x[42] ? _GEN17334 : _GEN17328;
wire  _GEN17336 = io_x[38] ? _GEN17335 : _GEN17325;
wire  _GEN17337 = io_x[10] ? _GEN17336 : _GEN17315;
wire  _GEN17338 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17339 = io_x[41] ? _GEN6836 : _GEN17338;
wire  _GEN17340 = io_x[14] ? _GEN6856 : _GEN17339;
wire  _GEN17341 = io_x[0] ? _GEN6858 : _GEN17340;
wire  _GEN17342 = io_x[76] ? _GEN17341 : _GEN6834;
wire  _GEN17343 = io_x[42] ? _GEN17342 : _GEN6863;
wire  _GEN17344 = io_x[38] ? _GEN17343 : _GEN6871;
wire  _GEN17345 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17346 = io_x[41] ? _GEN17345 : _GEN6836;
wire  _GEN17347 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17348 = io_x[41] ? _GEN17347 : _GEN6836;
wire  _GEN17349 = io_x[14] ? _GEN17348 : _GEN17346;
wire  _GEN17350 = io_x[0] ? _GEN17349 : _GEN6845;
wire  _GEN17351 = io_x[76] ? _GEN6834 : _GEN17350;
wire  _GEN17352 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17353 = io_x[6] ? _GEN17352 : _GEN6850;
wire  _GEN17354 = io_x[41] ? _GEN6836 : _GEN17353;
wire  _GEN17355 = io_x[14] ? _GEN17354 : _GEN6843;
wire  _GEN17356 = io_x[0] ? _GEN17355 : _GEN6845;
wire  _GEN17357 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17358 = io_x[6] ? _GEN6840 : _GEN17357;
wire  _GEN17359 = io_x[41] ? _GEN6836 : _GEN17358;
wire  _GEN17360 = io_x[14] ? _GEN6843 : _GEN17359;
wire  _GEN17361 = io_x[0] ? _GEN6858 : _GEN17360;
wire  _GEN17362 = io_x[76] ? _GEN17361 : _GEN17356;
wire  _GEN17363 = io_x[42] ? _GEN17362 : _GEN17351;
wire  _GEN17364 = io_x[38] ? _GEN17363 : _GEN6871;
wire  _GEN17365 = io_x[10] ? _GEN17364 : _GEN17344;
wire  _GEN17366 = io_x[71] ? _GEN17365 : _GEN17337;
wire  _GEN17367 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17368 = io_x[41] ? _GEN17367 : _GEN6836;
wire  _GEN17369 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17370 = io_x[41] ? _GEN17369 : _GEN6836;
wire  _GEN17371 = io_x[14] ? _GEN17370 : _GEN17368;
wire  _GEN17372 = io_x[0] ? _GEN6845 : _GEN17371;
wire  _GEN17373 = io_x[76] ? _GEN17372 : _GEN6834;
wire  _GEN17374 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17375 = io_x[6] ? _GEN6850 : _GEN17374;
wire  _GEN17376 = io_x[41] ? _GEN17375 : _GEN6836;
wire  _GEN17377 = io_x[14] ? _GEN6843 : _GEN17376;
wire  _GEN17378 = io_x[0] ? _GEN6845 : _GEN17377;
wire  _GEN17379 = io_x[76] ? _GEN17378 : _GEN6833;
wire  _GEN17380 = io_x[42] ? _GEN17379 : _GEN17373;
wire  _GEN17381 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17382 = io_x[6] ? _GEN6850 : _GEN17381;
wire  _GEN17383 = io_x[41] ? _GEN17382 : _GEN6836;
wire  _GEN17384 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17385 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17386 = io_x[6] ? _GEN17385 : _GEN17384;
wire  _GEN17387 = io_x[41] ? _GEN17386 : _GEN6836;
wire  _GEN17388 = io_x[14] ? _GEN17387 : _GEN17383;
wire  _GEN17389 = io_x[0] ? _GEN6845 : _GEN17388;
wire  _GEN17390 = io_x[76] ? _GEN17389 : _GEN6834;
wire  _GEN17391 = io_x[42] ? _GEN6874 : _GEN17390;
wire  _GEN17392 = io_x[38] ? _GEN17391 : _GEN17380;
wire  _GEN17393 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17394 = io_x[0] ? _GEN6845 : _GEN17393;
wire  _GEN17395 = io_x[76] ? _GEN17394 : _GEN6833;
wire  _GEN17396 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN17397 = io_x[76] ? _GEN6834 : _GEN17396;
wire  _GEN17398 = io_x[42] ? _GEN17397 : _GEN17395;
wire  _GEN17399 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17400 = io_x[6] ? _GEN6850 : _GEN17399;
wire  _GEN17401 = io_x[41] ? _GEN17400 : _GEN6836;
wire  _GEN17402 = io_x[14] ? _GEN6843 : _GEN17401;
wire  _GEN17403 = io_x[0] ? _GEN6845 : _GEN17402;
wire  _GEN17404 = io_x[76] ? _GEN17403 : _GEN6834;
wire  _GEN17405 = io_x[42] ? _GEN6874 : _GEN17404;
wire  _GEN17406 = io_x[38] ? _GEN17405 : _GEN17398;
wire  _GEN17407 = io_x[10] ? _GEN17406 : _GEN17392;
wire  _GEN17408 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN17409 = io_x[0] ? _GEN17408 : _GEN6858;
wire  _GEN17410 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17411 = io_x[6] ? _GEN6850 : _GEN17410;
wire  _GEN17412 = io_x[41] ? _GEN17411 : _GEN6836;
wire  _GEN17413 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17414 = io_x[41] ? _GEN17413 : _GEN6836;
wire  _GEN17415 = io_x[14] ? _GEN17414 : _GEN17412;
wire  _GEN17416 = io_x[0] ? _GEN17415 : _GEN6845;
wire  _GEN17417 = io_x[76] ? _GEN17416 : _GEN17409;
wire  _GEN17418 = io_x[42] ? _GEN17417 : _GEN6874;
wire  _GEN17419 = io_x[38] ? _GEN6871 : _GEN17418;
wire  _GEN17420 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17421 = io_x[6] ? _GEN17420 : _GEN6850;
wire  _GEN17422 = io_x[41] ? _GEN6836 : _GEN17421;
wire  _GEN17423 = io_x[14] ? _GEN17422 : _GEN6843;
wire  _GEN17424 = io_x[0] ? _GEN6858 : _GEN17423;
wire  _GEN17425 = io_x[76] ? _GEN6833 : _GEN17424;
wire  _GEN17426 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17427 = io_x[6] ? _GEN17426 : _GEN6840;
wire  _GEN17428 = io_x[41] ? _GEN17427 : _GEN6836;
wire  _GEN17429 = io_x[14] ? _GEN6856 : _GEN17428;
wire  _GEN17430 = io_x[0] ? _GEN17429 : _GEN6845;
wire  _GEN17431 = io_x[76] ? _GEN17430 : _GEN6833;
wire  _GEN17432 = io_x[42] ? _GEN17431 : _GEN17425;
wire  _GEN17433 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN17434 = io_x[2] ? _GEN17433 : _GEN6837;
wire  _GEN17435 = io_x[6] ? _GEN17434 : _GEN6850;
wire  _GEN17436 = io_x[41] ? _GEN6836 : _GEN17435;
wire  _GEN17437 = io_x[14] ? _GEN17436 : _GEN6843;
wire  _GEN17438 = io_x[0] ? _GEN6845 : _GEN17437;
wire  _GEN17439 = io_x[76] ? _GEN6834 : _GEN17438;
wire  _GEN17440 = io_x[42] ? _GEN6863 : _GEN17439;
wire  _GEN17441 = io_x[38] ? _GEN17440 : _GEN17432;
wire  _GEN17442 = io_x[10] ? _GEN17441 : _GEN17419;
wire  _GEN17443 = io_x[71] ? _GEN17442 : _GEN17407;
wire  _GEN17444 = io_x[70] ? _GEN17443 : _GEN17366;
wire  _GEN17445 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17446 = io_x[41] ? _GEN17445 : _GEN6836;
wire  _GEN17447 = io_x[14] ? _GEN17446 : _GEN6843;
wire  _GEN17448 = io_x[0] ? _GEN17447 : _GEN6845;
wire  _GEN17449 = io_x[76] ? _GEN6834 : _GEN17448;
wire  _GEN17450 = io_x[42] ? _GEN6874 : _GEN17449;
wire  _GEN17451 = io_x[38] ? _GEN17450 : _GEN6871;
wire  _GEN17452 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17453 = io_x[41] ? _GEN17452 : _GEN6836;
wire  _GEN17454 = io_x[14] ? _GEN17453 : _GEN6843;
wire  _GEN17455 = io_x[0] ? _GEN17454 : _GEN6845;
wire  _GEN17456 = io_x[76] ? _GEN6834 : _GEN17455;
wire  _GEN17457 = io_x[42] ? _GEN6874 : _GEN17456;
wire  _GEN17458 = io_x[38] ? _GEN17457 : _GEN6871;
wire  _GEN17459 = io_x[10] ? _GEN17458 : _GEN17451;
wire  _GEN17460 = io_x[71] ? _GEN7196 : _GEN17459;
wire  _GEN17461 = io_x[70] ? _GEN8474 : _GEN17460;
wire  _GEN17462 = io_x[33] ? _GEN17461 : _GEN17444;
wire  _GEN17463 = io_x[21] ? _GEN17462 : _GEN17300;
wire  _GEN17464 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN17465 = io_x[0] ? _GEN6845 : _GEN17464;
wire  _GEN17466 = io_x[76] ? _GEN17465 : _GEN6833;
wire  _GEN17467 = io_x[42] ? _GEN17466 : _GEN6863;
wire  _GEN17468 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17469 = io_x[6] ? _GEN6850 : _GEN17468;
wire  _GEN17470 = io_x[41] ? _GEN6836 : _GEN17469;
wire  _GEN17471 = io_x[14] ? _GEN6856 : _GEN17470;
wire  _GEN17472 = io_x[0] ? _GEN6845 : _GEN17471;
wire  _GEN17473 = io_x[76] ? _GEN17472 : _GEN6834;
wire  _GEN17474 = io_x[42] ? _GEN17473 : _GEN6863;
wire  _GEN17475 = io_x[38] ? _GEN17474 : _GEN17467;
wire  _GEN17476 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17477 = io_x[6] ? _GEN17476 : _GEN6850;
wire  _GEN17478 = io_x[41] ? _GEN17477 : _GEN6836;
wire  _GEN17479 = io_x[14] ? _GEN17478 : _GEN6843;
wire  _GEN17480 = io_x[0] ? _GEN17479 : _GEN6858;
wire  _GEN17481 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17482 = io_x[41] ? _GEN6836 : _GEN17481;
wire  _GEN17483 = io_x[14] ? _GEN17482 : _GEN6856;
wire  _GEN17484 = io_x[0] ? _GEN17483 : _GEN6845;
wire  _GEN17485 = io_x[76] ? _GEN17484 : _GEN17480;
wire  _GEN17486 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN17487 = io_x[42] ? _GEN17486 : _GEN17485;
wire  _GEN17488 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17489 = io_x[0] ? _GEN17488 : _GEN6845;
wire  _GEN17490 = io_x[76] ? _GEN17489 : _GEN6834;
wire  _GEN17491 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17492 = io_x[6] ? _GEN6850 : _GEN17491;
wire  _GEN17493 = io_x[41] ? _GEN6836 : _GEN17492;
wire  _GEN17494 = io_x[14] ? _GEN6856 : _GEN17493;
wire  _GEN17495 = io_x[0] ? _GEN6845 : _GEN17494;
wire  _GEN17496 = io_x[76] ? _GEN17495 : _GEN6833;
wire  _GEN17497 = io_x[42] ? _GEN17496 : _GEN17490;
wire  _GEN17498 = io_x[38] ? _GEN17497 : _GEN17487;
wire  _GEN17499 = io_x[10] ? _GEN17498 : _GEN17475;
wire  _GEN17500 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN17501 = io_x[0] ? _GEN6845 : _GEN17500;
wire  _GEN17502 = io_x[76] ? _GEN6834 : _GEN17501;
wire  _GEN17503 = io_x[42] ? _GEN6874 : _GEN17502;
wire  _GEN17504 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN17505 = io_x[76] ? _GEN6834 : _GEN17504;
wire  _GEN17506 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17507 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17508 = io_x[6] ? _GEN17507 : _GEN17506;
wire  _GEN17509 = io_x[41] ? _GEN6836 : _GEN17508;
wire  _GEN17510 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17511 = io_x[6] ? _GEN6850 : _GEN17510;
wire  _GEN17512 = io_x[41] ? _GEN6836 : _GEN17511;
wire  _GEN17513 = io_x[14] ? _GEN17512 : _GEN17509;
wire  _GEN17514 = io_x[0] ? _GEN6845 : _GEN17513;
wire  _GEN17515 = io_x[76] ? _GEN17514 : _GEN6834;
wire  _GEN17516 = io_x[42] ? _GEN17515 : _GEN17505;
wire  _GEN17517 = io_x[38] ? _GEN17516 : _GEN17503;
wire  _GEN17518 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17519 = io_x[41] ? _GEN6836 : _GEN17518;
wire  _GEN17520 = io_x[14] ? _GEN17519 : _GEN6843;
wire  _GEN17521 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17522 = io_x[41] ? _GEN17521 : _GEN6836;
wire  _GEN17523 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17524 = io_x[41] ? _GEN17523 : _GEN6924;
wire  _GEN17525 = io_x[14] ? _GEN17524 : _GEN17522;
wire  _GEN17526 = io_x[0] ? _GEN17525 : _GEN17520;
wire  _GEN17527 = io_x[76] ? _GEN6834 : _GEN17526;
wire  _GEN17528 = io_x[42] ? _GEN6863 : _GEN17527;
wire  _GEN17529 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17530 = io_x[41] ? _GEN17529 : _GEN6836;
wire  _GEN17531 = io_x[14] ? _GEN6856 : _GEN17530;
wire  _GEN17532 = io_x[0] ? _GEN6845 : _GEN17531;
wire  _GEN17533 = io_x[76] ? _GEN6834 : _GEN17532;
wire  _GEN17534 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17535 = io_x[6] ? _GEN6850 : _GEN17534;
wire  _GEN17536 = io_x[41] ? _GEN6836 : _GEN17535;
wire  _GEN17537 = io_x[14] ? _GEN6856 : _GEN17536;
wire  _GEN17538 = io_x[0] ? _GEN6845 : _GEN17537;
wire  _GEN17539 = io_x[76] ? _GEN17538 : _GEN6834;
wire  _GEN17540 = io_x[42] ? _GEN17539 : _GEN17533;
wire  _GEN17541 = io_x[38] ? _GEN17540 : _GEN17528;
wire  _GEN17542 = io_x[10] ? _GEN17541 : _GEN17517;
wire  _GEN17543 = io_x[71] ? _GEN17542 : _GEN17499;
wire  _GEN17544 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17545 = io_x[41] ? _GEN17544 : _GEN6836;
wire  _GEN17546 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17547 = io_x[41] ? _GEN17546 : _GEN6836;
wire  _GEN17548 = io_x[14] ? _GEN17547 : _GEN17545;
wire  _GEN17549 = io_x[0] ? _GEN6858 : _GEN17548;
wire  _GEN17550 = io_x[76] ? _GEN17549 : _GEN6833;
wire  _GEN17551 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN17552 = io_x[2] ? _GEN6837 : _GEN17551;
wire  _GEN17553 = io_x[6] ? _GEN6850 : _GEN17552;
wire  _GEN17554 = io_x[41] ? _GEN17553 : _GEN6836;
wire  _GEN17555 = io_x[14] ? _GEN6843 : _GEN17554;
wire  _GEN17556 = io_x[0] ? _GEN6845 : _GEN17555;
wire  _GEN17557 = io_x[76] ? _GEN17556 : _GEN6833;
wire  _GEN17558 = io_x[42] ? _GEN17557 : _GEN17550;
wire  _GEN17559 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17560 = io_x[6] ? _GEN6850 : _GEN17559;
wire  _GEN17561 = io_x[41] ? _GEN17560 : _GEN6836;
wire  _GEN17562 = io_x[14] ? _GEN6843 : _GEN17561;
wire  _GEN17563 = io_x[0] ? _GEN17562 : _GEN6845;
wire  _GEN17564 = io_x[76] ? _GEN17563 : _GEN6834;
wire  _GEN17565 = io_x[42] ? _GEN6874 : _GEN17564;
wire  _GEN17566 = io_x[38] ? _GEN17565 : _GEN17558;
wire  _GEN17567 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17568 = io_x[41] ? _GEN17567 : _GEN6924;
wire  _GEN17569 = io_x[14] ? _GEN17568 : _GEN6856;
wire  _GEN17570 = io_x[0] ? _GEN17569 : _GEN6845;
wire  _GEN17571 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17572 = io_x[41] ? _GEN17571 : _GEN6836;
wire  _GEN17573 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17574 = io_x[41] ? _GEN17573 : _GEN6836;
wire  _GEN17575 = io_x[14] ? _GEN17574 : _GEN17572;
wire  _GEN17576 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17577 = io_x[41] ? _GEN17576 : _GEN6836;
wire  _GEN17578 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN17579 = io_x[14] ? _GEN17578 : _GEN17577;
wire  _GEN17580 = io_x[0] ? _GEN17579 : _GEN17575;
wire  _GEN17581 = io_x[76] ? _GEN17580 : _GEN17570;
wire  _GEN17582 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN17583 = io_x[14] ? _GEN17582 : _GEN6843;
wire  _GEN17584 = io_x[0] ? _GEN17583 : _GEN6845;
wire  _GEN17585 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17586 = io_x[0] ? _GEN17585 : _GEN6845;
wire  _GEN17587 = io_x[76] ? _GEN17586 : _GEN17584;
wire  _GEN17588 = io_x[42] ? _GEN17587 : _GEN17581;
wire  _GEN17589 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17590 = io_x[41] ? _GEN17589 : _GEN6924;
wire  _GEN17591 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN17592 = io_x[14] ? _GEN17591 : _GEN17590;
wire  _GEN17593 = io_x[0] ? _GEN6858 : _GEN17592;
wire  _GEN17594 = io_x[76] ? _GEN17593 : _GEN6833;
wire  _GEN17595 = io_x[42] ? _GEN6863 : _GEN17594;
wire  _GEN17596 = io_x[38] ? _GEN17595 : _GEN17588;
wire  _GEN17597 = io_x[10] ? _GEN17596 : _GEN17566;
wire  _GEN17598 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17599 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17600 = io_x[41] ? _GEN17599 : _GEN6836;
wire  _GEN17601 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17602 = io_x[41] ? _GEN17601 : _GEN6836;
wire  _GEN17603 = io_x[14] ? _GEN17602 : _GEN17600;
wire  _GEN17604 = io_x[0] ? _GEN17603 : _GEN17598;
wire  _GEN17605 = io_x[76] ? _GEN17604 : _GEN6833;
wire  _GEN17606 = io_x[42] ? _GEN17605 : _GEN6874;
wire  _GEN17607 = io_x[38] ? _GEN6871 : _GEN17606;
wire  _GEN17608 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17609 = io_x[41] ? _GEN17608 : _GEN6924;
wire  _GEN17610 = io_x[14] ? _GEN17609 : _GEN6856;
wire  _GEN17611 = io_x[0] ? _GEN17610 : _GEN6845;
wire  _GEN17612 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN17613 = io_x[14] ? _GEN17612 : _GEN6843;
wire  _GEN17614 = io_x[0] ? _GEN17613 : _GEN6845;
wire  _GEN17615 = io_x[76] ? _GEN17614 : _GEN17611;
wire  _GEN17616 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17617 = io_x[41] ? _GEN17616 : _GEN6836;
wire  _GEN17618 = io_x[14] ? _GEN6856 : _GEN17617;
wire  _GEN17619 = io_x[0] ? _GEN17618 : _GEN6845;
wire  _GEN17620 = io_x[76] ? _GEN17619 : _GEN6834;
wire  _GEN17621 = io_x[42] ? _GEN17620 : _GEN17615;
wire  _GEN17622 = io_x[38] ? _GEN6871 : _GEN17621;
wire  _GEN17623 = io_x[10] ? _GEN17622 : _GEN17607;
wire  _GEN17624 = io_x[71] ? _GEN17623 : _GEN17597;
wire  _GEN17625 = io_x[70] ? _GEN17624 : _GEN17543;
wire  _GEN17626 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17627 = io_x[41] ? _GEN6836 : _GEN17626;
wire  _GEN17628 = io_x[14] ? _GEN17627 : _GEN6843;
wire  _GEN17629 = io_x[0] ? _GEN17628 : _GEN6845;
wire  _GEN17630 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17631 = io_x[0] ? _GEN17630 : _GEN6845;
wire  _GEN17632 = io_x[76] ? _GEN17631 : _GEN17629;
wire  _GEN17633 = io_x[42] ? _GEN17632 : _GEN6874;
wire  _GEN17634 = io_x[38] ? _GEN7036 : _GEN17633;
wire  _GEN17635 = io_x[10] ? _GEN17634 : _GEN7094;
wire  _GEN17636 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN17637 = io_x[76] ? _GEN6834 : _GEN17636;
wire  _GEN17638 = io_x[42] ? _GEN6874 : _GEN17637;
wire  _GEN17639 = io_x[38] ? _GEN17638 : _GEN6871;
wire  _GEN17640 = io_x[10] ? _GEN17639 : _GEN7044;
wire  _GEN17641 = io_x[71] ? _GEN17640 : _GEN17635;
wire  _GEN17642 = io_x[70] ? _GEN7020 : _GEN17641;
wire  _GEN17643 = io_x[33] ? _GEN17642 : _GEN17625;
wire  _GEN17644 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN17645 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17646 = io_x[6] ? _GEN6850 : _GEN17645;
wire  _GEN17647 = io_x[41] ? _GEN6836 : _GEN17646;
wire  _GEN17648 = io_x[14] ? _GEN6843 : _GEN17647;
wire  _GEN17649 = io_x[0] ? _GEN6845 : _GEN17648;
wire  _GEN17650 = io_x[76] ? _GEN17649 : _GEN17644;
wire  _GEN17651 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN17652 = io_x[14] ? _GEN17651 : _GEN6843;
wire  _GEN17653 = io_x[0] ? _GEN17652 : _GEN6858;
wire  _GEN17654 = io_x[76] ? _GEN6833 : _GEN17653;
wire  _GEN17655 = io_x[42] ? _GEN17654 : _GEN17650;
wire  _GEN17656 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17657 = io_x[41] ? _GEN17656 : _GEN6836;
wire  _GEN17658 = io_x[14] ? _GEN17657 : _GEN6856;
wire  _GEN17659 = io_x[0] ? _GEN17658 : _GEN6858;
wire  _GEN17660 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN17661 = io_x[14] ? _GEN6843 : _GEN17660;
wire  _GEN17662 = io_x[0] ? _GEN6845 : _GEN17661;
wire  _GEN17663 = io_x[76] ? _GEN17662 : _GEN17659;
wire  _GEN17664 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN17665 = io_x[2] ? _GEN6837 : _GEN17664;
wire  _GEN17666 = io_x[6] ? _GEN6850 : _GEN17665;
wire  _GEN17667 = io_x[41] ? _GEN17666 : _GEN6836;
wire  _GEN17668 = io_x[14] ? _GEN6843 : _GEN17667;
wire  _GEN17669 = io_x[0] ? _GEN6845 : _GEN17668;
wire  _GEN17670 = io_x[76] ? _GEN17669 : _GEN6834;
wire  _GEN17671 = io_x[42] ? _GEN17670 : _GEN17663;
wire  _GEN17672 = io_x[38] ? _GEN17671 : _GEN17655;
wire  _GEN17673 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17674 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17675 = io_x[6] ? _GEN17674 : _GEN6850;
wire  _GEN17676 = io_x[41] ? _GEN17675 : _GEN17673;
wire  _GEN17677 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17678 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17679 = io_x[6] ? _GEN17678 : _GEN6850;
wire  _GEN17680 = io_x[41] ? _GEN17679 : _GEN17677;
wire  _GEN17681 = io_x[14] ? _GEN17680 : _GEN17676;
wire  _GEN17682 = io_x[0] ? _GEN17681 : _GEN6858;
wire  _GEN17683 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17684 = io_x[41] ? _GEN6836 : _GEN17683;
wire  _GEN17685 = io_x[14] ? _GEN17684 : _GEN6856;
wire  _GEN17686 = io_x[0] ? _GEN17685 : _GEN6858;
wire  _GEN17687 = io_x[76] ? _GEN17686 : _GEN17682;
wire  _GEN17688 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN17689 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17690 = io_x[6] ? _GEN17689 : _GEN6850;
wire  _GEN17691 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN17692 = io_x[6] ? _GEN17691 : _GEN6840;
wire  _GEN17693 = io_x[41] ? _GEN17692 : _GEN17690;
wire  _GEN17694 = io_x[14] ? _GEN17693 : _GEN17688;
wire  _GEN17695 = io_x[0] ? _GEN17694 : _GEN6858;
wire  _GEN17696 = io_x[76] ? _GEN6834 : _GEN17695;
wire  _GEN17697 = io_x[42] ? _GEN17696 : _GEN17687;
wire  _GEN17698 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17699 = io_x[6] ? _GEN17698 : _GEN6850;
wire  _GEN17700 = io_x[41] ? _GEN17699 : _GEN6924;
wire  _GEN17701 = io_x[14] ? _GEN17700 : _GEN6843;
wire  _GEN17702 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17703 = io_x[6] ? _GEN17702 : _GEN6850;
wire  _GEN17704 = io_x[41] ? _GEN6924 : _GEN17703;
wire  _GEN17705 = io_x[14] ? _GEN17704 : _GEN6843;
wire  _GEN17706 = io_x[0] ? _GEN17705 : _GEN17701;
wire  _GEN17707 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17708 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN17709 = io_x[2] ? _GEN17708 : _GEN6837;
wire  _GEN17710 = io_x[6] ? _GEN17709 : _GEN6850;
wire  _GEN17711 = io_x[41] ? _GEN17710 : _GEN17707;
wire  _GEN17712 = io_x[14] ? _GEN17711 : _GEN6843;
wire  _GEN17713 = io_x[0] ? _GEN6858 : _GEN17712;
wire  _GEN17714 = io_x[76] ? _GEN17713 : _GEN17706;
wire  _GEN17715 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17716 = io_x[41] ? _GEN6924 : _GEN17715;
wire  _GEN17717 = io_x[14] ? _GEN17716 : _GEN6843;
wire  _GEN17718 = io_x[0] ? _GEN17717 : _GEN6845;
wire  _GEN17719 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN17720 = io_x[76] ? _GEN17719 : _GEN17718;
wire  _GEN17721 = io_x[42] ? _GEN17720 : _GEN17714;
wire  _GEN17722 = io_x[38] ? _GEN17721 : _GEN17697;
wire  _GEN17723 = io_x[10] ? _GEN17722 : _GEN17672;
wire  _GEN17724 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17725 = io_x[41] ? _GEN6836 : _GEN17724;
wire  _GEN17726 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17727 = io_x[41] ? _GEN6836 : _GEN17726;
wire  _GEN17728 = io_x[14] ? _GEN17727 : _GEN17725;
wire  _GEN17729 = io_x[0] ? _GEN17728 : _GEN6858;
wire  _GEN17730 = io_x[76] ? _GEN6834 : _GEN17729;
wire  _GEN17731 = io_x[42] ? _GEN6874 : _GEN17730;
wire  _GEN17732 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN17733 = io_x[2] ? _GEN6837 : _GEN17732;
wire  _GEN17734 = io_x[6] ? _GEN6840 : _GEN17733;
wire  _GEN17735 = io_x[41] ? _GEN6836 : _GEN17734;
wire  _GEN17736 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN17737 = io_x[14] ? _GEN17736 : _GEN17735;
wire  _GEN17738 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN17739 = io_x[0] ? _GEN17738 : _GEN17737;
wire  _GEN17740 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN17741 = io_x[2] ? _GEN6837 : _GEN17740;
wire  _GEN17742 = io_x[6] ? _GEN6850 : _GEN17741;
wire  _GEN17743 = io_x[41] ? _GEN17742 : _GEN6836;
wire  _GEN17744 = io_x[14] ? _GEN6856 : _GEN17743;
wire  _GEN17745 = io_x[0] ? _GEN6845 : _GEN17744;
wire  _GEN17746 = io_x[76] ? _GEN17745 : _GEN17739;
wire  _GEN17747 = io_x[42] ? _GEN6874 : _GEN17746;
wire  _GEN17748 = io_x[38] ? _GEN17747 : _GEN17731;
wire  _GEN17749 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17750 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17751 = io_x[41] ? _GEN17750 : _GEN17749;
wire  _GEN17752 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17753 = io_x[6] ? _GEN17752 : _GEN6850;
wire  _GEN17754 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17755 = io_x[41] ? _GEN17754 : _GEN17753;
wire  _GEN17756 = io_x[14] ? _GEN17755 : _GEN17751;
wire  _GEN17757 = io_x[0] ? _GEN17756 : _GEN6858;
wire  _GEN17758 = io_x[76] ? _GEN6833 : _GEN17757;
wire  _GEN17759 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17760 = io_x[41] ? _GEN6836 : _GEN17759;
wire  _GEN17761 = io_x[14] ? _GEN17760 : _GEN6843;
wire  _GEN17762 = io_x[0] ? _GEN6845 : _GEN17761;
wire  _GEN17763 = io_x[76] ? _GEN6834 : _GEN17762;
wire  _GEN17764 = io_x[42] ? _GEN17763 : _GEN17758;
wire  _GEN17765 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17766 = io_x[41] ? _GEN6924 : _GEN17765;
wire  _GEN17767 = io_x[14] ? _GEN17766 : _GEN6843;
wire  _GEN17768 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17769 = io_x[6] ? _GEN17768 : _GEN6850;
wire  _GEN17770 = io_x[41] ? _GEN6924 : _GEN17769;
wire  _GEN17771 = io_x[14] ? _GEN17770 : _GEN6856;
wire  _GEN17772 = io_x[0] ? _GEN17771 : _GEN17767;
wire  _GEN17773 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17774 = io_x[6] ? _GEN17773 : _GEN6850;
wire  _GEN17775 = io_x[41] ? _GEN17774 : _GEN6836;
wire  _GEN17776 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN17777 = io_x[14] ? _GEN17776 : _GEN17775;
wire  _GEN17778 = io_x[0] ? _GEN6858 : _GEN17777;
wire  _GEN17779 = io_x[76] ? _GEN17778 : _GEN17772;
wire  _GEN17780 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17781 = io_x[6] ? _GEN17780 : _GEN6850;
wire  _GEN17782 = io_x[41] ? _GEN6836 : _GEN17781;
wire  _GEN17783 = io_x[14] ? _GEN17782 : _GEN6843;
wire  _GEN17784 = io_x[0] ? _GEN17783 : _GEN6845;
wire  _GEN17785 = io_x[76] ? _GEN6834 : _GEN17784;
wire  _GEN17786 = io_x[42] ? _GEN17785 : _GEN17779;
wire  _GEN17787 = io_x[38] ? _GEN17786 : _GEN17764;
wire  _GEN17788 = io_x[10] ? _GEN17787 : _GEN17748;
wire  _GEN17789 = io_x[71] ? _GEN17788 : _GEN17723;
wire  _GEN17790 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN17791 = io_x[76] ? _GEN17790 : _GEN6834;
wire  _GEN17792 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN17793 = io_x[14] ? _GEN6843 : _GEN17792;
wire  _GEN17794 = io_x[0] ? _GEN6845 : _GEN17793;
wire  _GEN17795 = io_x[76] ? _GEN6833 : _GEN17794;
wire  _GEN17796 = io_x[42] ? _GEN17795 : _GEN17791;
wire  _GEN17797 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17798 = io_x[6] ? _GEN6850 : _GEN17797;
wire  _GEN17799 = io_x[41] ? _GEN6924 : _GEN17798;
wire  _GEN17800 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN17801 = io_x[14] ? _GEN17800 : _GEN17799;
wire  _GEN17802 = io_x[0] ? _GEN6845 : _GEN17801;
wire  _GEN17803 = io_x[76] ? _GEN17802 : _GEN6833;
wire  _GEN17804 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN17805 = io_x[42] ? _GEN17804 : _GEN17803;
wire  _GEN17806 = io_x[38] ? _GEN17805 : _GEN17796;
wire  _GEN17807 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17808 = io_x[41] ? _GEN6836 : _GEN17807;
wire  _GEN17809 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17810 = io_x[6] ? _GEN17809 : _GEN6850;
wire  _GEN17811 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17812 = io_x[41] ? _GEN17811 : _GEN17810;
wire  _GEN17813 = io_x[14] ? _GEN17812 : _GEN17808;
wire  _GEN17814 = io_x[0] ? _GEN17813 : _GEN6858;
wire  _GEN17815 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17816 = io_x[41] ? _GEN6836 : _GEN17815;
wire  _GEN17817 = io_x[14] ? _GEN17816 : _GEN6856;
wire  _GEN17818 = io_x[0] ? _GEN17817 : _GEN6845;
wire  _GEN17819 = io_x[76] ? _GEN17818 : _GEN17814;
wire  _GEN17820 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17821 = io_x[41] ? _GEN6836 : _GEN17820;
wire  _GEN17822 = io_x[14] ? _GEN17821 : _GEN6843;
wire  _GEN17823 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN17824 = io_x[14] ? _GEN17823 : _GEN6843;
wire  _GEN17825 = io_x[0] ? _GEN17824 : _GEN17822;
wire  _GEN17826 = io_x[76] ? _GEN6834 : _GEN17825;
wire  _GEN17827 = io_x[42] ? _GEN17826 : _GEN17819;
wire  _GEN17828 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17829 = io_x[0] ? _GEN17828 : _GEN6858;
wire  _GEN17830 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN17831 = io_x[6] ? _GEN6840 : _GEN17830;
wire  _GEN17832 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN17833 = io_x[2] ? _GEN17832 : _GEN6837;
wire  _GEN17834 = io_x[6] ? _GEN17833 : _GEN6850;
wire  _GEN17835 = io_x[41] ? _GEN17834 : _GEN17831;
wire  _GEN17836 = io_x[14] ? _GEN17835 : _GEN6856;
wire  _GEN17837 = io_x[0] ? _GEN6858 : _GEN17836;
wire  _GEN17838 = io_x[76] ? _GEN17837 : _GEN17829;
wire  _GEN17839 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17840 = io_x[41] ? _GEN17839 : _GEN6836;
wire  _GEN17841 = io_x[14] ? _GEN17840 : _GEN6843;
wire  _GEN17842 = io_x[0] ? _GEN17841 : _GEN6845;
wire  _GEN17843 = io_x[76] ? _GEN17842 : _GEN6834;
wire  _GEN17844 = io_x[42] ? _GEN17843 : _GEN17838;
wire  _GEN17845 = io_x[38] ? _GEN17844 : _GEN17827;
wire  _GEN17846 = io_x[10] ? _GEN17845 : _GEN17806;
wire  _GEN17847 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN17848 = io_x[76] ? _GEN6834 : _GEN17847;
wire  _GEN17849 = io_x[42] ? _GEN17848 : _GEN6863;
wire  _GEN17850 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN17851 = io_x[14] ? _GEN6843 : _GEN17850;
wire  _GEN17852 = io_x[0] ? _GEN6845 : _GEN17851;
wire  _GEN17853 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN17854 = io_x[14] ? _GEN6843 : _GEN17853;
wire  _GEN17855 = io_x[0] ? _GEN6845 : _GEN17854;
wire  _GEN17856 = io_x[76] ? _GEN17855 : _GEN17852;
wire  _GEN17857 = io_x[42] ? _GEN6874 : _GEN17856;
wire  _GEN17858 = io_x[38] ? _GEN17857 : _GEN17849;
wire  _GEN17859 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17860 = io_x[41] ? _GEN6924 : _GEN17859;
wire  _GEN17861 = io_x[14] ? _GEN17860 : _GEN6843;
wire  _GEN17862 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN17863 = io_x[2] ? _GEN17862 : _GEN6837;
wire  _GEN17864 = io_x[6] ? _GEN17863 : _GEN6850;
wire  _GEN17865 = io_x[41] ? _GEN6924 : _GEN17864;
wire  _GEN17866 = io_x[14] ? _GEN17865 : _GEN6843;
wire  _GEN17867 = io_x[0] ? _GEN17866 : _GEN17861;
wire  _GEN17868 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN17869 = io_x[0] ? _GEN17868 : _GEN6845;
wire  _GEN17870 = io_x[76] ? _GEN17869 : _GEN17867;
wire  _GEN17871 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17872 = io_x[41] ? _GEN6924 : _GEN17871;
wire  _GEN17873 = io_x[14] ? _GEN17872 : _GEN6843;
wire  _GEN17874 = io_x[0] ? _GEN17873 : _GEN6858;
wire  _GEN17875 = io_x[76] ? _GEN6833 : _GEN17874;
wire  _GEN17876 = io_x[42] ? _GEN17875 : _GEN17870;
wire  _GEN17877 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17878 = io_x[41] ? _GEN6836 : _GEN17877;
wire  _GEN17879 = io_x[14] ? _GEN17878 : _GEN6843;
wire  _GEN17880 = io_x[0] ? _GEN17879 : _GEN6858;
wire  _GEN17881 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN17882 = io_x[14] ? _GEN17881 : _GEN6843;
wire  _GEN17883 = io_x[0] ? _GEN6845 : _GEN17882;
wire  _GEN17884 = io_x[76] ? _GEN17883 : _GEN17880;
wire  _GEN17885 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17886 = io_x[0] ? _GEN17885 : _GEN6845;
wire  _GEN17887 = io_x[76] ? _GEN6834 : _GEN17886;
wire  _GEN17888 = io_x[42] ? _GEN17887 : _GEN17884;
wire  _GEN17889 = io_x[38] ? _GEN17888 : _GEN17876;
wire  _GEN17890 = io_x[10] ? _GEN17889 : _GEN17858;
wire  _GEN17891 = io_x[71] ? _GEN17890 : _GEN17846;
wire  _GEN17892 = io_x[70] ? _GEN17891 : _GEN17789;
wire  _GEN17893 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN17894 = io_x[38] ? _GEN17893 : _GEN7036;
wire  _GEN17895 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17896 = io_x[41] ? _GEN6836 : _GEN17895;
wire  _GEN17897 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17898 = io_x[41] ? _GEN6836 : _GEN17897;
wire  _GEN17899 = io_x[14] ? _GEN17898 : _GEN17896;
wire  _GEN17900 = io_x[0] ? _GEN17899 : _GEN6845;
wire  _GEN17901 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17902 = io_x[41] ? _GEN17901 : _GEN6836;
wire  _GEN17903 = io_x[14] ? _GEN17902 : _GEN6843;
wire  _GEN17904 = io_x[0] ? _GEN17903 : _GEN6845;
wire  _GEN17905 = io_x[76] ? _GEN17904 : _GEN17900;
wire  _GEN17906 = io_x[42] ? _GEN17905 : _GEN6874;
wire  _GEN17907 = io_x[38] ? _GEN7036 : _GEN17906;
wire  _GEN17908 = io_x[10] ? _GEN17907 : _GEN17894;
wire  _GEN17909 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN17910 = io_x[2] ? _GEN17909 : _GEN6837;
wire  _GEN17911 = io_x[6] ? _GEN17910 : _GEN6850;
wire  _GEN17912 = io_x[41] ? _GEN6836 : _GEN17911;
wire  _GEN17913 = io_x[14] ? _GEN17912 : _GEN6856;
wire  _GEN17914 = io_x[0] ? _GEN6845 : _GEN17913;
wire  _GEN17915 = io_x[76] ? _GEN6834 : _GEN17914;
wire  _GEN17916 = io_x[42] ? _GEN6874 : _GEN17915;
wire  _GEN17917 = io_x[38] ? _GEN17916 : _GEN6871;
wire  _GEN17918 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN17919 = io_x[41] ? _GEN6836 : _GEN17918;
wire  _GEN17920 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17921 = io_x[41] ? _GEN6924 : _GEN17920;
wire  _GEN17922 = io_x[14] ? _GEN17921 : _GEN17919;
wire  _GEN17923 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17924 = io_x[41] ? _GEN6836 : _GEN17923;
wire  _GEN17925 = io_x[14] ? _GEN17924 : _GEN6843;
wire  _GEN17926 = io_x[0] ? _GEN17925 : _GEN17922;
wire  _GEN17927 = io_x[76] ? _GEN6834 : _GEN17926;
wire  _GEN17928 = io_x[42] ? _GEN6874 : _GEN17927;
wire  _GEN17929 = io_x[38] ? _GEN17928 : _GEN6871;
wire  _GEN17930 = io_x[10] ? _GEN17929 : _GEN17917;
wire  _GEN17931 = io_x[71] ? _GEN17930 : _GEN17908;
wire  _GEN17932 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17933 = io_x[41] ? _GEN6836 : _GEN17932;
wire  _GEN17934 = io_x[14] ? _GEN17933 : _GEN6843;
wire  _GEN17935 = io_x[0] ? _GEN17934 : _GEN6845;
wire  _GEN17936 = io_x[76] ? _GEN6834 : _GEN17935;
wire  _GEN17937 = io_x[42] ? _GEN17936 : _GEN6863;
wire  _GEN17938 = io_x[38] ? _GEN6871 : _GEN17937;
wire  _GEN17939 = io_x[10] ? _GEN17938 : _GEN7044;
wire  _GEN17940 = io_x[71] ? _GEN17939 : _GEN7196;
wire  _GEN17941 = io_x[70] ? _GEN17940 : _GEN17931;
wire  _GEN17942 = io_x[33] ? _GEN17941 : _GEN17892;
wire  _GEN17943 = io_x[21] ? _GEN17942 : _GEN17643;
wire  _GEN17944 = io_x[18] ? _GEN17943 : _GEN17463;
wire  _GEN17945 = io_x[20] ? _GEN17944 : _GEN17181;
wire  _GEN17946 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN17947 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN17948 = io_x[2] ? _GEN6837 : _GEN17947;
wire  _GEN17949 = io_x[6] ? _GEN17948 : _GEN6840;
wire  _GEN17950 = io_x[41] ? _GEN6836 : _GEN17949;
wire  _GEN17951 = io_x[14] ? _GEN17950 : _GEN6843;
wire  _GEN17952 = io_x[0] ? _GEN6845 : _GEN17951;
wire  _GEN17953 = io_x[76] ? _GEN6834 : _GEN17952;
wire  _GEN17954 = io_x[42] ? _GEN6874 : _GEN17953;
wire  _GEN17955 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN17956 = io_x[42] ? _GEN6874 : _GEN17955;
wire  _GEN17957 = io_x[38] ? _GEN17956 : _GEN17954;
wire  _GEN17958 = io_x[10] ? _GEN17957 : _GEN17946;
wire  _GEN17959 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17960 = io_x[0] ? _GEN17959 : _GEN6845;
wire  _GEN17961 = io_x[76] ? _GEN6834 : _GEN17960;
wire  _GEN17962 = io_x[42] ? _GEN6863 : _GEN17961;
wire  _GEN17963 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN17964 = io_x[41] ? _GEN6836 : _GEN17963;
wire  _GEN17965 = io_x[14] ? _GEN17964 : _GEN6843;
wire  _GEN17966 = io_x[0] ? _GEN17965 : _GEN6845;
wire  _GEN17967 = io_x[76] ? _GEN6834 : _GEN17966;
wire  _GEN17968 = io_x[42] ? _GEN6874 : _GEN17967;
wire  _GEN17969 = io_x[38] ? _GEN17968 : _GEN17962;
wire  _GEN17970 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17971 = io_x[0] ? _GEN6845 : _GEN17970;
wire  _GEN17972 = io_x[76] ? _GEN6834 : _GEN17971;
wire  _GEN17973 = io_x[42] ? _GEN6874 : _GEN17972;
wire  _GEN17974 = io_x[38] ? _GEN6871 : _GEN17973;
wire  _GEN17975 = io_x[10] ? _GEN17974 : _GEN17969;
wire  _GEN17976 = io_x[71] ? _GEN17975 : _GEN17958;
wire  _GEN17977 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN17978 = io_x[2] ? _GEN6837 : _GEN17977;
wire  _GEN17979 = io_x[6] ? _GEN6850 : _GEN17978;
wire  _GEN17980 = io_x[41] ? _GEN17979 : _GEN6836;
wire  _GEN17981 = io_x[14] ? _GEN6843 : _GEN17980;
wire  _GEN17982 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN17983 = io_x[0] ? _GEN17982 : _GEN17981;
wire  _GEN17984 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN17985 = io_x[2] ? _GEN6837 : _GEN17984;
wire  _GEN17986 = io_x[6] ? _GEN6850 : _GEN17985;
wire  _GEN17987 = io_x[41] ? _GEN6836 : _GEN17986;
wire  _GEN17988 = io_x[14] ? _GEN17987 : _GEN6843;
wire  _GEN17989 = io_x[0] ? _GEN6845 : _GEN17988;
wire  _GEN17990 = io_x[76] ? _GEN17989 : _GEN17983;
wire  _GEN17991 = io_x[42] ? _GEN6874 : _GEN17990;
wire  _GEN17992 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN17993 = io_x[76] ? _GEN6834 : _GEN17992;
wire  _GEN17994 = io_x[42] ? _GEN6874 : _GEN17993;
wire  _GEN17995 = io_x[38] ? _GEN17994 : _GEN17991;
wire  _GEN17996 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN17997 = io_x[2] ? _GEN6837 : _GEN17996;
wire  _GEN17998 = io_x[6] ? _GEN17997 : _GEN6850;
wire  _GEN17999 = io_x[41] ? _GEN6836 : _GEN17998;
wire  _GEN18000 = io_x[14] ? _GEN17999 : _GEN6843;
wire  _GEN18001 = io_x[0] ? _GEN6845 : _GEN18000;
wire  _GEN18002 = io_x[76] ? _GEN18001 : _GEN6834;
wire  _GEN18003 = io_x[42] ? _GEN6874 : _GEN18002;
wire  _GEN18004 = io_x[38] ? _GEN7036 : _GEN18003;
wire  _GEN18005 = io_x[10] ? _GEN18004 : _GEN17995;
wire  _GEN18006 = io_x[71] ? _GEN18005 : _GEN7203;
wire  _GEN18007 = io_x[70] ? _GEN18006 : _GEN17976;
wire  _GEN18008 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN18009 = io_x[10] ? _GEN18008 : _GEN7044;
wire  _GEN18010 = io_x[71] ? _GEN18009 : _GEN7196;
wire  _GEN18011 = io_x[70] ? _GEN8474 : _GEN18010;
wire  _GEN18012 = io_x[33] ? _GEN18011 : _GEN18007;
wire  _GEN18013 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN18014 = io_x[14] ? _GEN6843 : _GEN18013;
wire  _GEN18015 = io_x[0] ? _GEN6845 : _GEN18014;
wire  _GEN18016 = io_x[76] ? _GEN6834 : _GEN18015;
wire  _GEN18017 = io_x[42] ? _GEN6874 : _GEN18016;
wire  _GEN18018 = io_x[38] ? _GEN18017 : _GEN6871;
wire  _GEN18019 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18020 = io_x[41] ? _GEN18019 : _GEN6836;
wire  _GEN18021 = io_x[14] ? _GEN18020 : _GEN6843;
wire  _GEN18022 = io_x[0] ? _GEN18021 : _GEN6845;
wire  _GEN18023 = io_x[76] ? _GEN6834 : _GEN18022;
wire  _GEN18024 = io_x[42] ? _GEN18023 : _GEN6863;
wire  _GEN18025 = io_x[38] ? _GEN18024 : _GEN7036;
wire  _GEN18026 = io_x[10] ? _GEN18025 : _GEN18018;
wire  _GEN18027 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN18028 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN18029 = io_x[42] ? _GEN18028 : _GEN6863;
wire  _GEN18030 = io_x[38] ? _GEN18029 : _GEN18027;
wire  _GEN18031 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN18032 = io_x[76] ? _GEN6834 : _GEN18031;
wire  _GEN18033 = io_x[42] ? _GEN18032 : _GEN6874;
wire  _GEN18034 = io_x[38] ? _GEN18033 : _GEN6871;
wire  _GEN18035 = io_x[10] ? _GEN18034 : _GEN18030;
wire  _GEN18036 = io_x[71] ? _GEN18035 : _GEN18026;
wire  _GEN18037 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18038 = io_x[41] ? _GEN18037 : _GEN6836;
wire  _GEN18039 = io_x[14] ? _GEN18038 : _GEN6843;
wire  _GEN18040 = io_x[0] ? _GEN18039 : _GEN6845;
wire  _GEN18041 = io_x[76] ? _GEN6834 : _GEN18040;
wire  _GEN18042 = io_x[42] ? _GEN18041 : _GEN6874;
wire  _GEN18043 = io_x[38] ? _GEN6871 : _GEN18042;
wire  _GEN18044 = io_x[10] ? _GEN18043 : _GEN7094;
wire  _GEN18045 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN18046 = io_x[76] ? _GEN18045 : _GEN6834;
wire  _GEN18047 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18048 = io_x[0] ? _GEN18047 : _GEN6858;
wire  _GEN18049 = io_x[76] ? _GEN6834 : _GEN18048;
wire  _GEN18050 = io_x[42] ? _GEN18049 : _GEN18046;
wire  _GEN18051 = io_x[38] ? _GEN7036 : _GEN18050;
wire  _GEN18052 = io_x[10] ? _GEN18051 : _GEN7094;
wire  _GEN18053 = io_x[71] ? _GEN18052 : _GEN18044;
wire  _GEN18054 = io_x[70] ? _GEN18053 : _GEN18036;
wire  _GEN18055 = io_x[33] ? _GEN12627 : _GEN18054;
wire  _GEN18056 = io_x[21] ? _GEN18055 : _GEN18012;
wire  _GEN18057 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN18058 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18059 = io_x[6] ? _GEN6840 : _GEN18058;
wire  _GEN18060 = io_x[41] ? _GEN18059 : _GEN6836;
wire  _GEN18061 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18062 = io_x[6] ? _GEN18061 : _GEN6840;
wire  _GEN18063 = io_x[41] ? _GEN18062 : _GEN6836;
wire  _GEN18064 = io_x[14] ? _GEN18063 : _GEN18060;
wire  _GEN18065 = io_x[0] ? _GEN18064 : _GEN6845;
wire  _GEN18066 = io_x[76] ? _GEN6834 : _GEN18065;
wire  _GEN18067 = io_x[42] ? _GEN18066 : _GEN6874;
wire  _GEN18068 = io_x[38] ? _GEN18067 : _GEN6871;
wire  _GEN18069 = io_x[10] ? _GEN18068 : _GEN18057;
wire  _GEN18070 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN18071 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18072 = io_x[6] ? _GEN18071 : _GEN6850;
wire  _GEN18073 = io_x[41] ? _GEN18072 : _GEN6836;
wire  _GEN18074 = io_x[14] ? _GEN18073 : _GEN6843;
wire  _GEN18075 = io_x[0] ? _GEN18074 : _GEN6845;
wire  _GEN18076 = io_x[76] ? _GEN6834 : _GEN18075;
wire  _GEN18077 = io_x[42] ? _GEN6863 : _GEN18076;
wire  _GEN18078 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN18079 = io_x[6] ? _GEN18078 : _GEN6850;
wire  _GEN18080 = io_x[41] ? _GEN18079 : _GEN6836;
wire  _GEN18081 = io_x[14] ? _GEN18080 : _GEN6843;
wire  _GEN18082 = io_x[0] ? _GEN18081 : _GEN6845;
wire  _GEN18083 = io_x[76] ? _GEN18082 : _GEN6833;
wire  _GEN18084 = io_x[42] ? _GEN6874 : _GEN18083;
wire  _GEN18085 = io_x[38] ? _GEN18084 : _GEN18077;
wire  _GEN18086 = io_x[10] ? _GEN18085 : _GEN18070;
wire  _GEN18087 = io_x[71] ? _GEN18086 : _GEN18069;
wire  _GEN18088 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18089 = io_x[0] ? _GEN18088 : _GEN6845;
wire  _GEN18090 = io_x[76] ? _GEN18089 : _GEN6834;
wire  _GEN18091 = io_x[42] ? _GEN18090 : _GEN6874;
wire  _GEN18092 = io_x[38] ? _GEN18091 : _GEN7036;
wire  _GEN18093 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18094 = io_x[0] ? _GEN18093 : _GEN6858;
wire  _GEN18095 = io_x[76] ? _GEN6834 : _GEN18094;
wire  _GEN18096 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18097 = io_x[41] ? _GEN18096 : _GEN6836;
wire  _GEN18098 = io_x[14] ? _GEN18097 : _GEN6843;
wire  _GEN18099 = io_x[0] ? _GEN6845 : _GEN18098;
wire  _GEN18100 = io_x[76] ? _GEN6834 : _GEN18099;
wire  _GEN18101 = io_x[42] ? _GEN18100 : _GEN18095;
wire  _GEN18102 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18103 = io_x[0] ? _GEN18102 : _GEN6845;
wire  _GEN18104 = io_x[76] ? _GEN18103 : _GEN6833;
wire  _GEN18105 = io_x[42] ? _GEN18104 : _GEN6874;
wire  _GEN18106 = io_x[38] ? _GEN18105 : _GEN18101;
wire  _GEN18107 = io_x[10] ? _GEN18106 : _GEN18092;
wire  _GEN18108 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18109 = io_x[6] ? _GEN18108 : _GEN6850;
wire  _GEN18110 = io_x[41] ? _GEN18109 : _GEN6836;
wire  _GEN18111 = io_x[14] ? _GEN18110 : _GEN6843;
wire  _GEN18112 = io_x[0] ? _GEN18111 : _GEN6845;
wire  _GEN18113 = io_x[76] ? _GEN18112 : _GEN6834;
wire  _GEN18114 = io_x[42] ? _GEN6874 : _GEN18113;
wire  _GEN18115 = io_x[38] ? _GEN6871 : _GEN18114;
wire  _GEN18116 = io_x[10] ? _GEN18115 : _GEN7094;
wire  _GEN18117 = io_x[71] ? _GEN18116 : _GEN18107;
wire  _GEN18118 = io_x[70] ? _GEN18117 : _GEN18087;
wire  _GEN18119 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18120 = io_x[0] ? _GEN18119 : _GEN6845;
wire  _GEN18121 = io_x[76] ? _GEN18120 : _GEN6834;
wire  _GEN18122 = io_x[42] ? _GEN18121 : _GEN6874;
wire  _GEN18123 = io_x[38] ? _GEN18122 : _GEN6871;
wire  _GEN18124 = io_x[10] ? _GEN18123 : _GEN7094;
wire  _GEN18125 = io_x[71] ? _GEN7196 : _GEN18124;
wire  _GEN18126 = io_x[70] ? _GEN18125 : _GEN7020;
wire  _GEN18127 = io_x[33] ? _GEN18126 : _GEN18118;
wire  _GEN18128 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN18129 = io_x[38] ? _GEN18128 : _GEN7036;
wire  _GEN18130 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18131 = io_x[0] ? _GEN18130 : _GEN6845;
wire  _GEN18132 = io_x[76] ? _GEN18131 : _GEN6834;
wire  _GEN18133 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18134 = io_x[41] ? _GEN18133 : _GEN6836;
wire  _GEN18135 = io_x[14] ? _GEN18134 : _GEN6843;
wire  _GEN18136 = io_x[0] ? _GEN18135 : _GEN6845;
wire  _GEN18137 = io_x[76] ? _GEN6834 : _GEN18136;
wire  _GEN18138 = io_x[42] ? _GEN18137 : _GEN18132;
wire  _GEN18139 = io_x[38] ? _GEN18138 : _GEN6871;
wire  _GEN18140 = io_x[10] ? _GEN18139 : _GEN18129;
wire  _GEN18141 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN18142 = io_x[38] ? _GEN7036 : _GEN18141;
wire  _GEN18143 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18144 = io_x[41] ? _GEN18143 : _GEN6836;
wire  _GEN18145 = io_x[14] ? _GEN18144 : _GEN6843;
wire  _GEN18146 = io_x[0] ? _GEN18145 : _GEN6845;
wire  _GEN18147 = io_x[76] ? _GEN6834 : _GEN18146;
wire  _GEN18148 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN18149 = io_x[42] ? _GEN18148 : _GEN18147;
wire  _GEN18150 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18151 = io_x[41] ? _GEN18150 : _GEN6836;
wire  _GEN18152 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18153 = io_x[41] ? _GEN18152 : _GEN6836;
wire  _GEN18154 = io_x[14] ? _GEN18153 : _GEN18151;
wire  _GEN18155 = io_x[0] ? _GEN18154 : _GEN6845;
wire  _GEN18156 = io_x[76] ? _GEN18155 : _GEN6833;
wire  _GEN18157 = io_x[42] ? _GEN6863 : _GEN18156;
wire  _GEN18158 = io_x[38] ? _GEN18157 : _GEN18149;
wire  _GEN18159 = io_x[10] ? _GEN18158 : _GEN18142;
wire  _GEN18160 = io_x[71] ? _GEN18159 : _GEN18140;
wire  _GEN18161 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN18162 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN18163 = io_x[14] ? _GEN18162 : _GEN6856;
wire  _GEN18164 = io_x[0] ? _GEN18163 : _GEN6858;
wire  _GEN18165 = io_x[76] ? _GEN6834 : _GEN18164;
wire  _GEN18166 = io_x[42] ? _GEN18165 : _GEN6874;
wire  _GEN18167 = io_x[38] ? _GEN18166 : _GEN18161;
wire  _GEN18168 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18169 = io_x[41] ? _GEN18168 : _GEN6836;
wire  _GEN18170 = io_x[14] ? _GEN18169 : _GEN6843;
wire  _GEN18171 = io_x[0] ? _GEN18170 : _GEN6858;
wire  _GEN18172 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18173 = io_x[0] ? _GEN6845 : _GEN18172;
wire  _GEN18174 = io_x[76] ? _GEN18173 : _GEN18171;
wire  _GEN18175 = io_x[42] ? _GEN18174 : _GEN6874;
wire  _GEN18176 = io_x[38] ? _GEN7036 : _GEN18175;
wire  _GEN18177 = io_x[10] ? _GEN18176 : _GEN18167;
wire  _GEN18178 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18179 = io_x[6] ? _GEN18178 : _GEN6850;
wire  _GEN18180 = io_x[41] ? _GEN18179 : _GEN6836;
wire  _GEN18181 = io_x[14] ? _GEN18180 : _GEN6843;
wire  _GEN18182 = io_x[0] ? _GEN18181 : _GEN6845;
wire  _GEN18183 = io_x[76] ? _GEN18182 : _GEN6834;
wire  _GEN18184 = io_x[42] ? _GEN6874 : _GEN18183;
wire  _GEN18185 = io_x[38] ? _GEN6871 : _GEN18184;
wire  _GEN18186 = io_x[10] ? _GEN18185 : _GEN7044;
wire  _GEN18187 = io_x[71] ? _GEN18186 : _GEN18177;
wire  _GEN18188 = io_x[70] ? _GEN18187 : _GEN18160;
wire  _GEN18189 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN18190 = io_x[71] ? _GEN18189 : _GEN7203;
wire  _GEN18191 = io_x[70] ? _GEN7020 : _GEN18190;
wire  _GEN18192 = io_x[33] ? _GEN18191 : _GEN18188;
wire  _GEN18193 = io_x[21] ? _GEN18192 : _GEN18127;
wire  _GEN18194 = io_x[18] ? _GEN18193 : _GEN18056;
wire  _GEN18195 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN18196 = io_x[14] ? _GEN18195 : _GEN6843;
wire  _GEN18197 = io_x[0] ? _GEN18196 : _GEN6845;
wire  _GEN18198 = io_x[76] ? _GEN6834 : _GEN18197;
wire  _GEN18199 = io_x[42] ? _GEN6874 : _GEN18198;
wire  _GEN18200 = io_x[38] ? _GEN6871 : _GEN18199;
wire  _GEN18201 = io_x[10] ? _GEN18200 : _GEN7044;
wire  _GEN18202 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN18203 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18204 = io_x[0] ? _GEN18203 : _GEN6845;
wire  _GEN18205 = io_x[76] ? _GEN6834 : _GEN18204;
wire  _GEN18206 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18207 = io_x[41] ? _GEN6836 : _GEN18206;
wire  _GEN18208 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18209 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18210 = io_x[6] ? _GEN18209 : _GEN6850;
wire  _GEN18211 = io_x[41] ? _GEN18210 : _GEN18208;
wire  _GEN18212 = io_x[14] ? _GEN18211 : _GEN18207;
wire  _GEN18213 = io_x[0] ? _GEN6845 : _GEN18212;
wire  _GEN18214 = io_x[76] ? _GEN6834 : _GEN18213;
wire  _GEN18215 = io_x[42] ? _GEN18214 : _GEN18205;
wire  _GEN18216 = io_x[38] ? _GEN18215 : _GEN6871;
wire  _GEN18217 = io_x[10] ? _GEN18216 : _GEN18202;
wire  _GEN18218 = io_x[71] ? _GEN18217 : _GEN18201;
wire  _GEN18219 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN18220 = io_x[38] ? _GEN6871 : _GEN18219;
wire  _GEN18221 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18222 = io_x[41] ? _GEN6836 : _GEN18221;
wire  _GEN18223 = io_x[14] ? _GEN18222 : _GEN6843;
wire  _GEN18224 = io_x[0] ? _GEN18223 : _GEN6845;
wire  _GEN18225 = io_x[76] ? _GEN6834 : _GEN18224;
wire  _GEN18226 = io_x[42] ? _GEN18225 : _GEN6863;
wire  _GEN18227 = io_x[38] ? _GEN6871 : _GEN18226;
wire  _GEN18228 = io_x[10] ? _GEN18227 : _GEN18220;
wire  _GEN18229 = io_x[71] ? _GEN18228 : _GEN7196;
wire  _GEN18230 = io_x[70] ? _GEN18229 : _GEN18218;
wire  _GEN18231 = io_x[71] ? _GEN7203 : _GEN7196;
wire  _GEN18232 = io_x[70] ? _GEN8474 : _GEN18231;
wire  _GEN18233 = io_x[33] ? _GEN18232 : _GEN18230;
wire  _GEN18234 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN18235 = io_x[14] ? _GEN6856 : _GEN18234;
wire  _GEN18236 = io_x[0] ? _GEN18235 : _GEN6845;
wire  _GEN18237 = io_x[76] ? _GEN6834 : _GEN18236;
wire  _GEN18238 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN18239 = io_x[42] ? _GEN18238 : _GEN18237;
wire  _GEN18240 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18241 = io_x[41] ? _GEN18240 : _GEN6836;
wire  _GEN18242 = io_x[14] ? _GEN18241 : _GEN6856;
wire  _GEN18243 = io_x[0] ? _GEN18242 : _GEN6845;
wire  _GEN18244 = io_x[76] ? _GEN6834 : _GEN18243;
wire  _GEN18245 = io_x[42] ? _GEN18244 : _GEN6874;
wire  _GEN18246 = io_x[38] ? _GEN18245 : _GEN18239;
wire  _GEN18247 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN18248 = io_x[2] ? _GEN6837 : _GEN18247;
wire  _GEN18249 = io_x[6] ? _GEN18248 : _GEN6850;
wire  _GEN18250 = io_x[41] ? _GEN6836 : _GEN18249;
wire  _GEN18251 = io_x[14] ? _GEN18250 : _GEN6856;
wire  _GEN18252 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18253 = io_x[0] ? _GEN18252 : _GEN18251;
wire  _GEN18254 = io_x[76] ? _GEN6834 : _GEN18253;
wire  _GEN18255 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN18256 = io_x[76] ? _GEN6834 : _GEN18255;
wire  _GEN18257 = io_x[42] ? _GEN18256 : _GEN18254;
wire  _GEN18258 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN18259 = io_x[6] ? _GEN18258 : _GEN6850;
wire  _GEN18260 = io_x[41] ? _GEN6836 : _GEN18259;
wire  _GEN18261 = io_x[14] ? _GEN18260 : _GEN6856;
wire  _GEN18262 = io_x[0] ? _GEN18261 : _GEN6845;
wire  _GEN18263 = io_x[76] ? _GEN6834 : _GEN18262;
wire  _GEN18264 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18265 = io_x[41] ? _GEN18264 : _GEN6836;
wire  _GEN18266 = io_x[14] ? _GEN18265 : _GEN6856;
wire  _GEN18267 = io_x[0] ? _GEN18266 : _GEN6845;
wire  _GEN18268 = io_x[76] ? _GEN6834 : _GEN18267;
wire  _GEN18269 = io_x[42] ? _GEN18268 : _GEN18263;
wire  _GEN18270 = io_x[38] ? _GEN18269 : _GEN18257;
wire  _GEN18271 = io_x[10] ? _GEN18270 : _GEN18246;
wire  _GEN18272 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18273 = io_x[41] ? _GEN6836 : _GEN18272;
wire  _GEN18274 = io_x[14] ? _GEN6843 : _GEN18273;
wire  _GEN18275 = io_x[0] ? _GEN18274 : _GEN6858;
wire  _GEN18276 = io_x[76] ? _GEN6834 : _GEN18275;
wire  _GEN18277 = io_x[42] ? _GEN18276 : _GEN6874;
wire  _GEN18278 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN18279 = io_x[42] ? _GEN6863 : _GEN18278;
wire  _GEN18280 = io_x[38] ? _GEN18279 : _GEN18277;
wire  _GEN18281 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN18282 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18283 = io_x[41] ? _GEN6836 : _GEN18282;
wire  _GEN18284 = io_x[14] ? _GEN18283 : _GEN6856;
wire  _GEN18285 = io_x[0] ? _GEN18284 : _GEN6845;
wire  _GEN18286 = io_x[76] ? _GEN6833 : _GEN18285;
wire  _GEN18287 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN18288 = io_x[6] ? _GEN18287 : _GEN6840;
wire  _GEN18289 = io_x[41] ? _GEN18288 : _GEN6836;
wire  _GEN18290 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18291 = io_x[6] ? _GEN18290 : _GEN6850;
wire  _GEN18292 = io_x[41] ? _GEN18291 : _GEN6924;
wire  _GEN18293 = io_x[14] ? _GEN18292 : _GEN18289;
wire  _GEN18294 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18295 = io_x[0] ? _GEN18294 : _GEN18293;
wire  _GEN18296 = io_x[76] ? _GEN6833 : _GEN18295;
wire  _GEN18297 = io_x[42] ? _GEN18296 : _GEN18286;
wire  _GEN18298 = io_x[38] ? _GEN18297 : _GEN18281;
wire  _GEN18299 = io_x[10] ? _GEN18298 : _GEN18280;
wire  _GEN18300 = io_x[71] ? _GEN18299 : _GEN18271;
wire  _GEN18301 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN18302 = io_x[76] ? _GEN6834 : _GEN18301;
wire  _GEN18303 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN18304 = io_x[14] ? _GEN6843 : _GEN18303;
wire  _GEN18305 = io_x[0] ? _GEN6858 : _GEN18304;
wire  _GEN18306 = io_x[76] ? _GEN6834 : _GEN18305;
wire  _GEN18307 = io_x[42] ? _GEN18306 : _GEN18302;
wire  _GEN18308 = io_x[38] ? _GEN7036 : _GEN18307;
wire  _GEN18309 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18310 = io_x[0] ? _GEN6858 : _GEN18309;
wire  _GEN18311 = io_x[76] ? _GEN6834 : _GEN18310;
wire  _GEN18312 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18313 = io_x[41] ? _GEN18312 : _GEN6836;
wire  _GEN18314 = io_x[14] ? _GEN18313 : _GEN6843;
wire  _GEN18315 = io_x[0] ? _GEN18314 : _GEN6858;
wire  _GEN18316 = io_x[76] ? _GEN6834 : _GEN18315;
wire  _GEN18317 = io_x[42] ? _GEN18316 : _GEN18311;
wire  _GEN18318 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18319 = io_x[41] ? _GEN18318 : _GEN6836;
wire  _GEN18320 = io_x[14] ? _GEN6843 : _GEN18319;
wire  _GEN18321 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18322 = io_x[41] ? _GEN18321 : _GEN6836;
wire  _GEN18323 = io_x[14] ? _GEN18322 : _GEN6843;
wire  _GEN18324 = io_x[0] ? _GEN18323 : _GEN18320;
wire  _GEN18325 = io_x[76] ? _GEN6834 : _GEN18324;
wire  _GEN18326 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18327 = io_x[6] ? _GEN18326 : _GEN6850;
wire  _GEN18328 = io_x[41] ? _GEN18327 : _GEN6924;
wire  _GEN18329 = io_x[14] ? _GEN18328 : _GEN6843;
wire  _GEN18330 = io_x[0] ? _GEN18329 : _GEN6858;
wire  _GEN18331 = io_x[76] ? _GEN6834 : _GEN18330;
wire  _GEN18332 = io_x[42] ? _GEN18331 : _GEN18325;
wire  _GEN18333 = io_x[38] ? _GEN18332 : _GEN18317;
wire  _GEN18334 = io_x[10] ? _GEN18333 : _GEN18308;
wire  _GEN18335 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN18336 = io_x[76] ? _GEN6834 : _GEN18335;
wire  _GEN18337 = io_x[42] ? _GEN18336 : _GEN6863;
wire  _GEN18338 = io_x[38] ? _GEN7036 : _GEN18337;
wire  _GEN18339 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18340 = io_x[41] ? _GEN6836 : _GEN18339;
wire  _GEN18341 = io_x[14] ? _GEN6856 : _GEN18340;
wire  _GEN18342 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18343 = io_x[0] ? _GEN18342 : _GEN18341;
wire  _GEN18344 = io_x[76] ? _GEN6834 : _GEN18343;
wire  _GEN18345 = io_x[42] ? _GEN18344 : _GEN6863;
wire  _GEN18346 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18347 = io_x[0] ? _GEN18346 : _GEN6858;
wire  _GEN18348 = io_x[76] ? _GEN6834 : _GEN18347;
wire  _GEN18349 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18350 = io_x[41] ? _GEN18349 : _GEN6836;
wire  _GEN18351 = io_x[14] ? _GEN18350 : _GEN6843;
wire  _GEN18352 = io_x[0] ? _GEN18351 : _GEN6858;
wire  _GEN18353 = io_x[76] ? _GEN6833 : _GEN18352;
wire  _GEN18354 = io_x[42] ? _GEN18353 : _GEN18348;
wire  _GEN18355 = io_x[38] ? _GEN18354 : _GEN18345;
wire  _GEN18356 = io_x[10] ? _GEN18355 : _GEN18338;
wire  _GEN18357 = io_x[71] ? _GEN18356 : _GEN18334;
wire  _GEN18358 = io_x[70] ? _GEN18357 : _GEN18300;
wire  _GEN18359 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18360 = io_x[0] ? _GEN6845 : _GEN18359;
wire  _GEN18361 = io_x[76] ? _GEN6834 : _GEN18360;
wire  _GEN18362 = io_x[42] ? _GEN6874 : _GEN18361;
wire  _GEN18363 = io_x[38] ? _GEN18362 : _GEN6871;
wire  _GEN18364 = io_x[10] ? _GEN18363 : _GEN7044;
wire  _GEN18365 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN18366 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN18367 = io_x[38] ? _GEN18366 : _GEN18365;
wire  _GEN18368 = io_x[10] ? _GEN18367 : _GEN7044;
wire  _GEN18369 = io_x[71] ? _GEN18368 : _GEN18364;
wire  _GEN18370 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN18371 = io_x[38] ? _GEN18370 : _GEN6871;
wire  _GEN18372 = io_x[10] ? _GEN18371 : _GEN7044;
wire  _GEN18373 = io_x[71] ? _GEN7196 : _GEN18372;
wire  _GEN18374 = io_x[70] ? _GEN18373 : _GEN18369;
wire  _GEN18375 = io_x[33] ? _GEN18374 : _GEN18358;
wire  _GEN18376 = io_x[21] ? _GEN18375 : _GEN18233;
wire  _GEN18377 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN18378 = io_x[14] ? _GEN18377 : _GEN6843;
wire  _GEN18379 = io_x[0] ? _GEN18378 : _GEN6845;
wire  _GEN18380 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18381 = io_x[41] ? _GEN6836 : _GEN18380;
wire  _GEN18382 = io_x[14] ? _GEN18381 : _GEN6843;
wire  _GEN18383 = io_x[0] ? _GEN6845 : _GEN18382;
wire  _GEN18384 = io_x[76] ? _GEN18383 : _GEN18379;
wire  _GEN18385 = io_x[42] ? _GEN6863 : _GEN18384;
wire  _GEN18386 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18387 = io_x[6] ? _GEN6840 : _GEN18386;
wire  _GEN18388 = io_x[41] ? _GEN6924 : _GEN18387;
wire  _GEN18389 = io_x[14] ? _GEN18388 : _GEN6856;
wire  _GEN18390 = io_x[0] ? _GEN6845 : _GEN18389;
wire  _GEN18391 = io_x[76] ? _GEN6834 : _GEN18390;
wire  _GEN18392 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN18393 = io_x[76] ? _GEN6834 : _GEN18392;
wire  _GEN18394 = io_x[42] ? _GEN18393 : _GEN18391;
wire  _GEN18395 = io_x[38] ? _GEN18394 : _GEN18385;
wire  _GEN18396 = io_x[10] ? _GEN18395 : _GEN7094;
wire  _GEN18397 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN18398 = io_x[42] ? _GEN6874 : _GEN18397;
wire  _GEN18399 = io_x[38] ? _GEN18398 : _GEN6871;
wire  _GEN18400 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18401 = io_x[0] ? _GEN18400 : _GEN6845;
wire  _GEN18402 = io_x[76] ? _GEN6834 : _GEN18401;
wire  _GEN18403 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18404 = io_x[0] ? _GEN18403 : _GEN6845;
wire  _GEN18405 = io_x[76] ? _GEN6833 : _GEN18404;
wire  _GEN18406 = io_x[42] ? _GEN18405 : _GEN18402;
wire  _GEN18407 = io_x[38] ? _GEN18406 : _GEN7036;
wire  _GEN18408 = io_x[10] ? _GEN18407 : _GEN18399;
wire  _GEN18409 = io_x[71] ? _GEN18408 : _GEN18396;
wire  _GEN18410 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN18411 = io_x[42] ? _GEN6863 : _GEN18410;
wire  _GEN18412 = io_x[38] ? _GEN7036 : _GEN18411;
wire  _GEN18413 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN18414 = io_x[76] ? _GEN6834 : _GEN18413;
wire  _GEN18415 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18416 = io_x[0] ? _GEN6845 : _GEN18415;
wire  _GEN18417 = io_x[76] ? _GEN6834 : _GEN18416;
wire  _GEN18418 = io_x[42] ? _GEN18417 : _GEN18414;
wire  _GEN18419 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN18420 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18421 = io_x[0] ? _GEN18420 : _GEN6845;
wire  _GEN18422 = io_x[76] ? _GEN6834 : _GEN18421;
wire  _GEN18423 = io_x[42] ? _GEN18422 : _GEN18419;
wire  _GEN18424 = io_x[38] ? _GEN18423 : _GEN18418;
wire  _GEN18425 = io_x[10] ? _GEN18424 : _GEN18412;
wire  _GEN18426 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18427 = io_x[0] ? _GEN18426 : _GEN6858;
wire  _GEN18428 = io_x[76] ? _GEN6834 : _GEN18427;
wire  _GEN18429 = io_x[42] ? _GEN18428 : _GEN6863;
wire  _GEN18430 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN18431 = io_x[14] ? _GEN18430 : _GEN6856;
wire  _GEN18432 = io_x[0] ? _GEN18431 : _GEN6845;
wire  _GEN18433 = io_x[76] ? _GEN6834 : _GEN18432;
wire  _GEN18434 = io_x[42] ? _GEN18433 : _GEN6874;
wire  _GEN18435 = io_x[38] ? _GEN18434 : _GEN18429;
wire  _GEN18436 = io_x[10] ? _GEN18435 : _GEN7094;
wire  _GEN18437 = io_x[71] ? _GEN18436 : _GEN18425;
wire  _GEN18438 = io_x[70] ? _GEN18437 : _GEN18409;
wire  _GEN18439 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN18440 = io_x[71] ? _GEN7196 : _GEN18439;
wire  _GEN18441 = io_x[70] ? _GEN18440 : _GEN8474;
wire  _GEN18442 = io_x[33] ? _GEN18441 : _GEN18438;
wire  _GEN18443 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18444 = io_x[41] ? _GEN18443 : _GEN6836;
wire  _GEN18445 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18446 = io_x[41] ? _GEN6924 : _GEN18445;
wire  _GEN18447 = io_x[14] ? _GEN18446 : _GEN18444;
wire  _GEN18448 = io_x[0] ? _GEN18447 : _GEN6845;
wire  _GEN18449 = io_x[76] ? _GEN6834 : _GEN18448;
wire  _GEN18450 = io_x[42] ? _GEN6863 : _GEN18449;
wire  _GEN18451 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18452 = io_x[41] ? _GEN6836 : _GEN18451;
wire  _GEN18453 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18454 = io_x[41] ? _GEN6836 : _GEN18453;
wire  _GEN18455 = io_x[14] ? _GEN18454 : _GEN18452;
wire  _GEN18456 = io_x[0] ? _GEN18455 : _GEN6845;
wire  _GEN18457 = io_x[76] ? _GEN18456 : _GEN6833;
wire  _GEN18458 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18459 = io_x[41] ? _GEN6924 : _GEN18458;
wire  _GEN18460 = io_x[14] ? _GEN18459 : _GEN6856;
wire  _GEN18461 = io_x[0] ? _GEN6845 : _GEN18460;
wire  _GEN18462 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN18463 = io_x[6] ? _GEN6850 : _GEN18462;
wire  _GEN18464 = io_x[41] ? _GEN18463 : _GEN6836;
wire  _GEN18465 = io_x[14] ? _GEN6843 : _GEN18464;
wire  _GEN18466 = io_x[0] ? _GEN18465 : _GEN6845;
wire  _GEN18467 = io_x[76] ? _GEN18466 : _GEN18461;
wire  _GEN18468 = io_x[42] ? _GEN18467 : _GEN18457;
wire  _GEN18469 = io_x[38] ? _GEN18468 : _GEN18450;
wire  _GEN18470 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18471 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18472 = io_x[6] ? _GEN18471 : _GEN6850;
wire  _GEN18473 = io_x[41] ? _GEN18472 : _GEN6924;
wire  _GEN18474 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18475 = io_x[41] ? _GEN18474 : _GEN6836;
wire  _GEN18476 = io_x[14] ? _GEN18475 : _GEN18473;
wire  _GEN18477 = io_x[0] ? _GEN18476 : _GEN18470;
wire  _GEN18478 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18479 = io_x[0] ? _GEN18478 : _GEN6845;
wire  _GEN18480 = io_x[76] ? _GEN18479 : _GEN18477;
wire  _GEN18481 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN18482 = io_x[2] ? _GEN18481 : _GEN6837;
wire  _GEN18483 = io_x[6] ? _GEN18482 : _GEN6840;
wire  _GEN18484 = io_x[41] ? _GEN18483 : _GEN6836;
wire  _GEN18485 = io_x[14] ? _GEN18484 : _GEN6843;
wire  _GEN18486 = io_x[0] ? _GEN6845 : _GEN18485;
wire  _GEN18487 = io_x[76] ? _GEN18486 : _GEN6833;
wire  _GEN18488 = io_x[42] ? _GEN18487 : _GEN18480;
wire  _GEN18489 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18490 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18491 = io_x[6] ? _GEN18490 : _GEN6850;
wire  _GEN18492 = io_x[41] ? _GEN18491 : _GEN6836;
wire  _GEN18493 = io_x[14] ? _GEN18492 : _GEN6843;
wire  _GEN18494 = io_x[0] ? _GEN18493 : _GEN18489;
wire  _GEN18495 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18496 = io_x[41] ? _GEN6836 : _GEN18495;
wire  _GEN18497 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18498 = io_x[41] ? _GEN6836 : _GEN18497;
wire  _GEN18499 = io_x[14] ? _GEN18498 : _GEN18496;
wire  _GEN18500 = io_x[0] ? _GEN18499 : _GEN6845;
wire  _GEN18501 = io_x[76] ? _GEN18500 : _GEN18494;
wire  _GEN18502 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18503 = io_x[41] ? _GEN6924 : _GEN18502;
wire  _GEN18504 = io_x[14] ? _GEN18503 : _GEN6843;
wire  _GEN18505 = io_x[0] ? _GEN6858 : _GEN18504;
wire  _GEN18506 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18507 = io_x[41] ? _GEN18506 : _GEN6836;
wire  _GEN18508 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18509 = io_x[41] ? _GEN18508 : _GEN6836;
wire  _GEN18510 = io_x[14] ? _GEN18509 : _GEN18507;
wire  _GEN18511 = io_x[0] ? _GEN18510 : _GEN6845;
wire  _GEN18512 = io_x[76] ? _GEN18511 : _GEN18505;
wire  _GEN18513 = io_x[42] ? _GEN18512 : _GEN18501;
wire  _GEN18514 = io_x[38] ? _GEN18513 : _GEN18488;
wire  _GEN18515 = io_x[10] ? _GEN18514 : _GEN18469;
wire  _GEN18516 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18517 = io_x[6] ? _GEN18516 : _GEN6850;
wire  _GEN18518 = io_x[41] ? _GEN18517 : _GEN6924;
wire  _GEN18519 = io_x[14] ? _GEN6843 : _GEN18518;
wire  _GEN18520 = io_x[0] ? _GEN18519 : _GEN6845;
wire  _GEN18521 = io_x[76] ? _GEN6834 : _GEN18520;
wire  _GEN18522 = io_x[42] ? _GEN6863 : _GEN18521;
wire  _GEN18523 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18524 = io_x[41] ? _GEN6836 : _GEN18523;
wire  _GEN18525 = io_x[14] ? _GEN6843 : _GEN18524;
wire  _GEN18526 = io_x[0] ? _GEN18525 : _GEN6845;
wire  _GEN18527 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18528 = io_x[41] ? _GEN18527 : _GEN6836;
wire  _GEN18529 = io_x[14] ? _GEN6843 : _GEN18528;
wire  _GEN18530 = io_x[0] ? _GEN18529 : _GEN6845;
wire  _GEN18531 = io_x[76] ? _GEN18530 : _GEN18526;
wire  _GEN18532 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN18533 = io_x[42] ? _GEN18532 : _GEN18531;
wire  _GEN18534 = io_x[38] ? _GEN18533 : _GEN18522;
wire  _GEN18535 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18536 = io_x[6] ? _GEN18535 : _GEN6850;
wire  _GEN18537 = io_x[41] ? _GEN18536 : _GEN6836;
wire  _GEN18538 = io_x[14] ? _GEN18537 : _GEN6843;
wire  _GEN18539 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN18540 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN18541 = io_x[2] ? _GEN18540 : _GEN6837;
wire  _GEN18542 = io_x[6] ? _GEN18541 : _GEN6850;
wire  _GEN18543 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN18544 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18545 = io_x[6] ? _GEN18544 : _GEN18543;
wire  _GEN18546 = io_x[41] ? _GEN18545 : _GEN18542;
wire  _GEN18547 = io_x[14] ? _GEN18546 : _GEN18539;
wire  _GEN18548 = io_x[0] ? _GEN18547 : _GEN18538;
wire  _GEN18549 = io_x[76] ? _GEN6834 : _GEN18548;
wire  _GEN18550 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18551 = io_x[41] ? _GEN6836 : _GEN18550;
wire  _GEN18552 = io_x[14] ? _GEN18551 : _GEN6843;
wire  _GEN18553 = io_x[0] ? _GEN6845 : _GEN18552;
wire  _GEN18554 = io_x[76] ? _GEN18553 : _GEN6833;
wire  _GEN18555 = io_x[42] ? _GEN18554 : _GEN18549;
wire  _GEN18556 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18557 = io_x[41] ? _GEN6836 : _GEN18556;
wire  _GEN18558 = io_x[14] ? _GEN18557 : _GEN6843;
wire  _GEN18559 = io_x[0] ? _GEN18558 : _GEN6845;
wire  _GEN18560 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18561 = io_x[41] ? _GEN18560 : _GEN6836;
wire  _GEN18562 = io_x[14] ? _GEN18561 : _GEN6856;
wire  _GEN18563 = io_x[0] ? _GEN18562 : _GEN6858;
wire  _GEN18564 = io_x[76] ? _GEN18563 : _GEN18559;
wire  _GEN18565 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18566 = io_x[41] ? _GEN6836 : _GEN18565;
wire  _GEN18567 = io_x[14] ? _GEN18566 : _GEN6843;
wire  _GEN18568 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18569 = io_x[41] ? _GEN18568 : _GEN6836;
wire  _GEN18570 = io_x[14] ? _GEN18569 : _GEN6843;
wire  _GEN18571 = io_x[0] ? _GEN18570 : _GEN18567;
wire  _GEN18572 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18573 = io_x[0] ? _GEN18572 : _GEN6845;
wire  _GEN18574 = io_x[76] ? _GEN18573 : _GEN18571;
wire  _GEN18575 = io_x[42] ? _GEN18574 : _GEN18564;
wire  _GEN18576 = io_x[38] ? _GEN18575 : _GEN18555;
wire  _GEN18577 = io_x[10] ? _GEN18576 : _GEN18534;
wire  _GEN18578 = io_x[71] ? _GEN18577 : _GEN18515;
wire  _GEN18579 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN18580 = io_x[2] ? _GEN6837 : _GEN18579;
wire  _GEN18581 = io_x[6] ? _GEN6840 : _GEN18580;
wire  _GEN18582 = io_x[41] ? _GEN18581 : _GEN6836;
wire  _GEN18583 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18584 = io_x[6] ? _GEN6850 : _GEN18583;
wire  _GEN18585 = io_x[41] ? _GEN18584 : _GEN6836;
wire  _GEN18586 = io_x[14] ? _GEN18585 : _GEN18582;
wire  _GEN18587 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18588 = io_x[41] ? _GEN18587 : _GEN6924;
wire  _GEN18589 = io_x[14] ? _GEN6843 : _GEN18588;
wire  _GEN18590 = io_x[0] ? _GEN18589 : _GEN18586;
wire  _GEN18591 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18592 = io_x[0] ? _GEN18591 : _GEN6845;
wire  _GEN18593 = io_x[76] ? _GEN18592 : _GEN18590;
wire  _GEN18594 = io_x[42] ? _GEN6863 : _GEN18593;
wire  _GEN18595 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN18596 = io_x[14] ? _GEN6843 : _GEN18595;
wire  _GEN18597 = io_x[0] ? _GEN6858 : _GEN18596;
wire  _GEN18598 = io_x[76] ? _GEN6834 : _GEN18597;
wire  _GEN18599 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18600 = io_x[0] ? _GEN18599 : _GEN6858;
wire  _GEN18601 = io_x[76] ? _GEN6834 : _GEN18600;
wire  _GEN18602 = io_x[42] ? _GEN18601 : _GEN18598;
wire  _GEN18603 = io_x[38] ? _GEN18602 : _GEN18594;
wire  _GEN18604 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18605 = io_x[44] ? _GEN6913 : _GEN6914;
wire  _GEN18606 = io_x[2] ? _GEN18605 : _GEN6837;
wire  _GEN18607 = io_x[6] ? _GEN18606 : _GEN6850;
wire  _GEN18608 = io_x[41] ? _GEN18607 : _GEN6836;
wire  _GEN18609 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18610 = io_x[6] ? _GEN18609 : _GEN6850;
wire  _GEN18611 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN18612 = io_x[2] ? _GEN18611 : _GEN6837;
wire  _GEN18613 = io_x[6] ? _GEN18612 : _GEN6850;
wire  _GEN18614 = io_x[41] ? _GEN18613 : _GEN18610;
wire  _GEN18615 = io_x[14] ? _GEN18614 : _GEN18608;
wire  _GEN18616 = io_x[0] ? _GEN18615 : _GEN18604;
wire  _GEN18617 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN18618 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN18619 = io_x[6] ? _GEN18618 : _GEN6850;
wire  _GEN18620 = io_x[41] ? _GEN18619 : _GEN6836;
wire  _GEN18621 = io_x[14] ? _GEN18620 : _GEN18617;
wire  _GEN18622 = io_x[0] ? _GEN18621 : _GEN6845;
wire  _GEN18623 = io_x[76] ? _GEN18622 : _GEN18616;
wire  _GEN18624 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN18625 = io_x[14] ? _GEN18624 : _GEN6856;
wire  _GEN18626 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18627 = io_x[0] ? _GEN18626 : _GEN18625;
wire  _GEN18628 = io_x[76] ? _GEN6833 : _GEN18627;
wire  _GEN18629 = io_x[42] ? _GEN18628 : _GEN18623;
wire  _GEN18630 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18631 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18632 = io_x[0] ? _GEN18631 : _GEN18630;
wire  _GEN18633 = io_x[76] ? _GEN6834 : _GEN18632;
wire  _GEN18634 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN18635 = io_x[2] ? _GEN18634 : _GEN6837;
wire  _GEN18636 = io_x[6] ? _GEN18635 : _GEN6850;
wire  _GEN18637 = io_x[41] ? _GEN18636 : _GEN6924;
wire  _GEN18638 = io_x[14] ? _GEN18637 : _GEN6843;
wire  _GEN18639 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN18640 = io_x[6] ? _GEN18639 : _GEN6840;
wire  _GEN18641 = io_x[41] ? _GEN18640 : _GEN6836;
wire  _GEN18642 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18643 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18644 = io_x[6] ? _GEN18643 : _GEN6850;
wire  _GEN18645 = io_x[41] ? _GEN18644 : _GEN18642;
wire  _GEN18646 = io_x[14] ? _GEN18645 : _GEN18641;
wire  _GEN18647 = io_x[0] ? _GEN18646 : _GEN18638;
wire  _GEN18648 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18649 = io_x[41] ? _GEN6924 : _GEN18648;
wire  _GEN18650 = io_x[14] ? _GEN18649 : _GEN6843;
wire  _GEN18651 = io_x[0] ? _GEN18650 : _GEN6845;
wire  _GEN18652 = io_x[76] ? _GEN18651 : _GEN18647;
wire  _GEN18653 = io_x[42] ? _GEN18652 : _GEN18633;
wire  _GEN18654 = io_x[38] ? _GEN18653 : _GEN18629;
wire  _GEN18655 = io_x[10] ? _GEN18654 : _GEN18603;
wire  _GEN18656 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18657 = io_x[6] ? _GEN6850 : _GEN18656;
wire  _GEN18658 = io_x[41] ? _GEN6836 : _GEN18657;
wire  _GEN18659 = io_x[14] ? _GEN6843 : _GEN18658;
wire  _GEN18660 = io_x[0] ? _GEN18659 : _GEN6845;
wire  _GEN18661 = io_x[76] ? _GEN6834 : _GEN18660;
wire  _GEN18662 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN18663 = io_x[76] ? _GEN6834 : _GEN18662;
wire  _GEN18664 = io_x[42] ? _GEN18663 : _GEN18661;
wire  _GEN18665 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN18666 = io_x[2] ? _GEN6837 : _GEN18665;
wire  _GEN18667 = io_x[6] ? _GEN6850 : _GEN18666;
wire  _GEN18668 = io_x[41] ? _GEN6836 : _GEN18667;
wire  _GEN18669 = io_x[14] ? _GEN6843 : _GEN18668;
wire  _GEN18670 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18671 = io_x[41] ? _GEN6836 : _GEN18670;
wire  _GEN18672 = io_x[14] ? _GEN18671 : _GEN6843;
wire  _GEN18673 = io_x[0] ? _GEN18672 : _GEN18669;
wire  _GEN18674 = io_x[76] ? _GEN6834 : _GEN18673;
wire  _GEN18675 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN18676 = io_x[76] ? _GEN6834 : _GEN18675;
wire  _GEN18677 = io_x[42] ? _GEN18676 : _GEN18674;
wire  _GEN18678 = io_x[38] ? _GEN18677 : _GEN18664;
wire  _GEN18679 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18680 = io_x[41] ? _GEN6836 : _GEN18679;
wire  _GEN18681 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18682 = io_x[41] ? _GEN6924 : _GEN18681;
wire  _GEN18683 = io_x[14] ? _GEN18682 : _GEN18680;
wire  _GEN18684 = io_x[0] ? _GEN18683 : _GEN6845;
wire  _GEN18685 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18686 = io_x[41] ? _GEN6836 : _GEN18685;
wire  _GEN18687 = io_x[14] ? _GEN18686 : _GEN6856;
wire  _GEN18688 = io_x[44] ? _GEN6914 : _GEN6913;
wire  _GEN18689 = io_x[2] ? _GEN18688 : _GEN6837;
wire  _GEN18690 = io_x[6] ? _GEN18689 : _GEN6840;
wire  _GEN18691 = io_x[41] ? _GEN18690 : _GEN6836;
wire  _GEN18692 = io_x[14] ? _GEN18691 : _GEN6856;
wire  _GEN18693 = io_x[0] ? _GEN18692 : _GEN18687;
wire  _GEN18694 = io_x[76] ? _GEN18693 : _GEN18684;
wire  _GEN18695 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN18696 = io_x[14] ? _GEN6856 : _GEN18695;
wire  _GEN18697 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18698 = io_x[41] ? _GEN6924 : _GEN18697;
wire  _GEN18699 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18700 = io_x[41] ? _GEN6924 : _GEN18699;
wire  _GEN18701 = io_x[14] ? _GEN18700 : _GEN18698;
wire  _GEN18702 = io_x[0] ? _GEN18701 : _GEN18696;
wire  _GEN18703 = io_x[76] ? _GEN6834 : _GEN18702;
wire  _GEN18704 = io_x[42] ? _GEN18703 : _GEN18694;
wire  _GEN18705 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18706 = io_x[0] ? _GEN18705 : _GEN6845;
wire  _GEN18707 = io_x[76] ? _GEN6834 : _GEN18706;
wire  _GEN18708 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18709 = io_x[6] ? _GEN18708 : _GEN6850;
wire  _GEN18710 = io_x[41] ? _GEN18709 : _GEN6924;
wire  _GEN18711 = io_x[14] ? _GEN18710 : _GEN6843;
wire  _GEN18712 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18713 = io_x[41] ? _GEN18712 : _GEN6836;
wire  _GEN18714 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18715 = io_x[41] ? _GEN18714 : _GEN6924;
wire  _GEN18716 = io_x[14] ? _GEN18715 : _GEN18713;
wire  _GEN18717 = io_x[0] ? _GEN18716 : _GEN18711;
wire  _GEN18718 = io_x[76] ? _GEN6833 : _GEN18717;
wire  _GEN18719 = io_x[42] ? _GEN18718 : _GEN18707;
wire  _GEN18720 = io_x[38] ? _GEN18719 : _GEN18704;
wire  _GEN18721 = io_x[10] ? _GEN18720 : _GEN18678;
wire  _GEN18722 = io_x[71] ? _GEN18721 : _GEN18655;
wire  _GEN18723 = io_x[70] ? _GEN18722 : _GEN18578;
wire  _GEN18724 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18725 = io_x[41] ? _GEN6836 : _GEN18724;
wire  _GEN18726 = io_x[14] ? _GEN18725 : _GEN6843;
wire  _GEN18727 = io_x[0] ? _GEN18726 : _GEN6845;
wire  _GEN18728 = io_x[76] ? _GEN18727 : _GEN6834;
wire  _GEN18729 = io_x[42] ? _GEN6863 : _GEN18728;
wire  _GEN18730 = io_x[38] ? _GEN18729 : _GEN6871;
wire  _GEN18731 = io_x[10] ? _GEN18730 : _GEN7044;
wire  _GEN18732 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN18733 = io_x[10] ? _GEN7094 : _GEN18732;
wire  _GEN18734 = io_x[71] ? _GEN18733 : _GEN18731;
wire  _GEN18735 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18736 = io_x[0] ? _GEN18735 : _GEN6845;
wire  _GEN18737 = io_x[76] ? _GEN18736 : _GEN6834;
wire  _GEN18738 = io_x[42] ? _GEN18737 : _GEN6863;
wire  _GEN18739 = io_x[38] ? _GEN18738 : _GEN6871;
wire  _GEN18740 = io_x[10] ? _GEN18739 : _GEN7094;
wire  _GEN18741 = io_x[71] ? _GEN7196 : _GEN18740;
wire  _GEN18742 = io_x[70] ? _GEN18741 : _GEN18734;
wire  _GEN18743 = io_x[33] ? _GEN18742 : _GEN18723;
wire  _GEN18744 = io_x[21] ? _GEN18743 : _GEN18442;
wire  _GEN18745 = io_x[18] ? _GEN18744 : _GEN18376;
wire  _GEN18746 = io_x[20] ? _GEN18745 : _GEN18194;
wire  _GEN18747 = io_x[45] ? _GEN18746 : _GEN17945;
wire  _GEN18748 = io_x[28] ? _GEN18747 : _GEN16548;
wire  _GEN18749 = io_x[79] ? _GEN18748 : _GEN14455;
wire  _GEN18750 = io_x[70] ? _GEN7020 : _GEN8474;
wire  _GEN18751 = io_x[33] ? _GEN12627 : _GEN18750;
wire  _GEN18752 = io_x[21] ? _GEN18751 : _GEN12643;
wire  _GEN18753 = io_x[21] ? _GEN12933 : _GEN12643;
wire  _GEN18754 = io_x[18] ? _GEN18753 : _GEN18752;
wire  _GEN18755 = io_x[20] ? _GEN18754 : _GEN14273;
wire  _GEN18756 = 1'b0;
wire  _GEN18757 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN18758 = io_x[76] ? _GEN6834 : _GEN18757;
wire  _GEN18759 = io_x[42] ? _GEN18758 : _GEN6874;
wire  _GEN18760 = io_x[38] ? _GEN6871 : _GEN18759;
wire  _GEN18761 = io_x[10] ? _GEN7094 : _GEN18760;
wire  _GEN18762 = io_x[71] ? _GEN18761 : _GEN7203;
wire  _GEN18763 = io_x[70] ? _GEN18762 : _GEN7020;
wire  _GEN18764 = io_x[33] ? _GEN12627 : _GEN18763;
wire  _GEN18765 = io_x[21] ? _GEN18764 : _GEN12643;
wire  _GEN18766 = io_x[18] ? _GEN14264 : _GEN18765;
wire  _GEN18767 = io_x[20] ? _GEN18766 : _GEN18756;
wire  _GEN18768 = io_x[45] ? _GEN18767 : _GEN18755;
wire  _GEN18769 = io_x[70] ? _GEN7020 : _GEN8474;
wire  _GEN18770 = io_x[33] ? _GEN12627 : _GEN18769;
wire  _GEN18771 = io_x[21] ? _GEN12643 : _GEN18770;
wire  _GEN18772 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18773 = io_x[0] ? _GEN6845 : _GEN18772;
wire  _GEN18774 = io_x[76] ? _GEN18773 : _GEN6834;
wire  _GEN18775 = io_x[42] ? _GEN18774 : _GEN6874;
wire  _GEN18776 = io_x[38] ? _GEN18775 : _GEN6871;
wire  _GEN18777 = io_x[10] ? _GEN18776 : _GEN7044;
wire  _GEN18778 = io_x[71] ? _GEN18777 : _GEN7196;
wire  _GEN18779 = io_x[70] ? _GEN18778 : _GEN8474;
wire  _GEN18780 = io_x[33] ? _GEN12627 : _GEN18779;
wire  _GEN18781 = io_x[21] ? _GEN12643 : _GEN18780;
wire  _GEN18782 = io_x[18] ? _GEN18781 : _GEN18771;
wire  _GEN18783 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN18784 = io_x[38] ? _GEN18783 : _GEN6871;
wire  _GEN18785 = io_x[10] ? _GEN7044 : _GEN18784;
wire  _GEN18786 = io_x[71] ? _GEN18785 : _GEN7196;
wire  _GEN18787 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN18788 = io_x[71] ? _GEN18787 : _GEN7196;
wire  _GEN18789 = io_x[70] ? _GEN18788 : _GEN18786;
wire  _GEN18790 = io_x[33] ? _GEN12627 : _GEN18789;
wire  _GEN18791 = io_x[21] ? _GEN18790 : _GEN12643;
wire  _GEN18792 = io_x[71] ? _GEN7196 : _GEN7203;
wire  _GEN18793 = io_x[70] ? _GEN18792 : _GEN8474;
wire  _GEN18794 = io_x[33] ? _GEN12627 : _GEN18793;
wire  _GEN18795 = io_x[21] ? _GEN18794 : _GEN12643;
wire  _GEN18796 = io_x[18] ? _GEN18795 : _GEN18791;
wire  _GEN18797 = io_x[20] ? _GEN18796 : _GEN18782;
wire  _GEN18798 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN18799 = io_x[10] ? _GEN7044 : _GEN18798;
wire  _GEN18800 = io_x[71] ? _GEN7203 : _GEN18799;
wire  _GEN18801 = io_x[70] ? _GEN18800 : _GEN8474;
wire  _GEN18802 = io_x[33] ? _GEN12627 : _GEN18801;
wire  _GEN18803 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN18804 = io_x[10] ? _GEN7044 : _GEN18803;
wire  _GEN18805 = io_x[71] ? _GEN18804 : _GEN7203;
wire  _GEN18806 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN18807 = io_x[38] ? _GEN6871 : _GEN18806;
wire  _GEN18808 = io_x[10] ? _GEN7094 : _GEN18807;
wire  _GEN18809 = io_x[71] ? _GEN18808 : _GEN7203;
wire  _GEN18810 = io_x[70] ? _GEN18809 : _GEN18805;
wire  _GEN18811 = io_x[33] ? _GEN12627 : _GEN18810;
wire  _GEN18812 = io_x[21] ? _GEN18811 : _GEN18802;
wire  _GEN18813 = io_x[18] ? _GEN12920 : _GEN18812;
wire  _GEN18814 = io_x[71] ? _GEN7196 : _GEN7203;
wire  _GEN18815 = io_x[70] ? _GEN18814 : _GEN8474;
wire  _GEN18816 = io_x[33] ? _GEN12627 : _GEN18815;
wire  _GEN18817 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN18818 = io_x[71] ? _GEN7203 : _GEN18817;
wire  _GEN18819 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN18820 = io_x[71] ? _GEN7203 : _GEN18819;
wire  _GEN18821 = io_x[70] ? _GEN18820 : _GEN18818;
wire  _GEN18822 = io_x[33] ? _GEN12627 : _GEN18821;
wire  _GEN18823 = io_x[21] ? _GEN18822 : _GEN18816;
wire  _GEN18824 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN18825 = io_x[10] ? _GEN18824 : _GEN7044;
wire  _GEN18826 = io_x[71] ? _GEN7196 : _GEN18825;
wire  _GEN18827 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN18828 = io_x[10] ? _GEN18827 : _GEN7044;
wire  _GEN18829 = io_x[71] ? _GEN18828 : _GEN7196;
wire  _GEN18830 = io_x[70] ? _GEN18829 : _GEN18826;
wire  _GEN18831 = io_x[33] ? _GEN12627 : _GEN18830;
wire  _GEN18832 = io_x[21] ? _GEN18831 : _GEN12643;
wire  _GEN18833 = io_x[18] ? _GEN18832 : _GEN18823;
wire  _GEN18834 = io_x[20] ? _GEN18833 : _GEN18813;
wire  _GEN18835 = io_x[45] ? _GEN18834 : _GEN18797;
wire  _GEN18836 = io_x[28] ? _GEN18835 : _GEN18768;
wire  _GEN18837 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN18838 = io_x[42] ? _GEN18837 : _GEN6874;
wire  _GEN18839 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18840 = io_x[41] ? _GEN6836 : _GEN18839;
wire  _GEN18841 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18842 = io_x[41] ? _GEN6836 : _GEN18841;
wire  _GEN18843 = io_x[14] ? _GEN18842 : _GEN18840;
wire  _GEN18844 = io_x[0] ? _GEN6845 : _GEN18843;
wire  _GEN18845 = io_x[76] ? _GEN18844 : _GEN6834;
wire  _GEN18846 = io_x[42] ? _GEN18845 : _GEN6863;
wire  _GEN18847 = io_x[38] ? _GEN18846 : _GEN18838;
wire  _GEN18848 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18849 = io_x[41] ? _GEN6836 : _GEN18848;
wire  _GEN18850 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18851 = io_x[41] ? _GEN6836 : _GEN18850;
wire  _GEN18852 = io_x[14] ? _GEN18851 : _GEN18849;
wire  _GEN18853 = io_x[0] ? _GEN6845 : _GEN18852;
wire  _GEN18854 = io_x[76] ? _GEN18853 : _GEN6834;
wire  _GEN18855 = io_x[42] ? _GEN18854 : _GEN6874;
wire  _GEN18856 = io_x[38] ? _GEN18855 : _GEN6871;
wire  _GEN18857 = io_x[10] ? _GEN18856 : _GEN18847;
wire  _GEN18858 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18859 = io_x[41] ? _GEN18858 : _GEN6836;
wire  _GEN18860 = io_x[14] ? _GEN6856 : _GEN18859;
wire  _GEN18861 = io_x[0] ? _GEN6845 : _GEN18860;
wire  _GEN18862 = io_x[76] ? _GEN18861 : _GEN6834;
wire  _GEN18863 = io_x[42] ? _GEN18862 : _GEN6874;
wire  _GEN18864 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN18865 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18866 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18867 = io_x[41] ? _GEN6836 : _GEN18866;
wire  _GEN18868 = io_x[14] ? _GEN6856 : _GEN18867;
wire  _GEN18869 = io_x[0] ? _GEN18868 : _GEN18865;
wire  _GEN18870 = io_x[76] ? _GEN18869 : _GEN6834;
wire  _GEN18871 = io_x[42] ? _GEN18870 : _GEN18864;
wire  _GEN18872 = io_x[38] ? _GEN18871 : _GEN18863;
wire  _GEN18873 = io_x[10] ? _GEN7094 : _GEN18872;
wire  _GEN18874 = io_x[71] ? _GEN18873 : _GEN18857;
wire  _GEN18875 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18876 = io_x[41] ? _GEN18875 : _GEN6836;
wire  _GEN18877 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN18878 = io_x[14] ? _GEN18877 : _GEN18876;
wire  _GEN18879 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN18880 = io_x[14] ? _GEN18879 : _GEN6856;
wire  _GEN18881 = io_x[0] ? _GEN18880 : _GEN18878;
wire  _GEN18882 = io_x[76] ? _GEN18881 : _GEN6833;
wire  _GEN18883 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN18884 = io_x[42] ? _GEN18883 : _GEN18882;
wire  _GEN18885 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18886 = io_x[41] ? _GEN18885 : _GEN6836;
wire  _GEN18887 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18888 = io_x[41] ? _GEN18887 : _GEN6836;
wire  _GEN18889 = io_x[14] ? _GEN18888 : _GEN18886;
wire  _GEN18890 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18891 = io_x[41] ? _GEN18890 : _GEN6836;
wire  _GEN18892 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18893 = io_x[41] ? _GEN18892 : _GEN6836;
wire  _GEN18894 = io_x[14] ? _GEN18893 : _GEN18891;
wire  _GEN18895 = io_x[0] ? _GEN18894 : _GEN18889;
wire  _GEN18896 = io_x[76] ? _GEN18895 : _GEN6834;
wire  _GEN18897 = io_x[42] ? _GEN6874 : _GEN18896;
wire  _GEN18898 = io_x[38] ? _GEN18897 : _GEN18884;
wire  _GEN18899 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN18900 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18901 = io_x[0] ? _GEN18900 : _GEN18899;
wire  _GEN18902 = io_x[76] ? _GEN18901 : _GEN6834;
wire  _GEN18903 = io_x[42] ? _GEN6874 : _GEN18902;
wire  _GEN18904 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18905 = io_x[41] ? _GEN18904 : _GEN6836;
wire  _GEN18906 = io_x[14] ? _GEN6843 : _GEN18905;
wire  _GEN18907 = io_x[0] ? _GEN6845 : _GEN18906;
wire  _GEN18908 = io_x[76] ? _GEN18907 : _GEN6834;
wire  _GEN18909 = io_x[42] ? _GEN6874 : _GEN18908;
wire  _GEN18910 = io_x[38] ? _GEN18909 : _GEN18903;
wire  _GEN18911 = io_x[10] ? _GEN18910 : _GEN18898;
wire  _GEN18912 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18913 = io_x[0] ? _GEN6845 : _GEN18912;
wire  _GEN18914 = io_x[76] ? _GEN18913 : _GEN6834;
wire  _GEN18915 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN18916 = io_x[42] ? _GEN18915 : _GEN18914;
wire  _GEN18917 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN18918 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18919 = io_x[41] ? _GEN18918 : _GEN6836;
wire  _GEN18920 = io_x[14] ? _GEN6843 : _GEN18919;
wire  _GEN18921 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18922 = io_x[41] ? _GEN6836 : _GEN18921;
wire  _GEN18923 = io_x[14] ? _GEN6843 : _GEN18922;
wire  _GEN18924 = io_x[0] ? _GEN18923 : _GEN18920;
wire  _GEN18925 = io_x[76] ? _GEN18924 : _GEN6833;
wire  _GEN18926 = io_x[42] ? _GEN18925 : _GEN18917;
wire  _GEN18927 = io_x[38] ? _GEN18926 : _GEN18916;
wire  _GEN18928 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18929 = io_x[41] ? _GEN6836 : _GEN18928;
wire  _GEN18930 = io_x[14] ? _GEN6843 : _GEN18929;
wire  _GEN18931 = io_x[0] ? _GEN6845 : _GEN18930;
wire  _GEN18932 = io_x[76] ? _GEN18931 : _GEN6834;
wire  _GEN18933 = io_x[42] ? _GEN6863 : _GEN18932;
wire  _GEN18934 = io_x[38] ? _GEN6871 : _GEN18933;
wire  _GEN18935 = io_x[10] ? _GEN18934 : _GEN18927;
wire  _GEN18936 = io_x[71] ? _GEN18935 : _GEN18911;
wire  _GEN18937 = io_x[70] ? _GEN18936 : _GEN18874;
wire  _GEN18938 = io_x[33] ? _GEN12627 : _GEN18937;
wire  _GEN18939 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18940 = io_x[41] ? _GEN6836 : _GEN18939;
wire  _GEN18941 = io_x[14] ? _GEN6843 : _GEN18940;
wire  _GEN18942 = io_x[0] ? _GEN6845 : _GEN18941;
wire  _GEN18943 = io_x[76] ? _GEN18942 : _GEN6833;
wire  _GEN18944 = io_x[42] ? _GEN18943 : _GEN6874;
wire  _GEN18945 = io_x[38] ? _GEN18944 : _GEN6871;
wire  _GEN18946 = io_x[10] ? _GEN7044 : _GEN18945;
wire  _GEN18947 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18948 = io_x[6] ? _GEN6850 : _GEN18947;
wire  _GEN18949 = io_x[41] ? _GEN18948 : _GEN6836;
wire  _GEN18950 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18951 = io_x[6] ? _GEN18950 : _GEN6840;
wire  _GEN18952 = io_x[41] ? _GEN18951 : _GEN6836;
wire  _GEN18953 = io_x[14] ? _GEN18952 : _GEN18949;
wire  _GEN18954 = io_x[0] ? _GEN6845 : _GEN18953;
wire  _GEN18955 = io_x[76] ? _GEN18954 : _GEN6834;
wire  _GEN18956 = io_x[42] ? _GEN18955 : _GEN6874;
wire  _GEN18957 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN18958 = io_x[41] ? _GEN6836 : _GEN18957;
wire  _GEN18959 = io_x[14] ? _GEN6843 : _GEN18958;
wire  _GEN18960 = io_x[0] ? _GEN18959 : _GEN6845;
wire  _GEN18961 = io_x[76] ? _GEN18960 : _GEN6834;
wire  _GEN18962 = io_x[42] ? _GEN18961 : _GEN6874;
wire  _GEN18963 = io_x[38] ? _GEN18962 : _GEN18956;
wire  _GEN18964 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN18965 = io_x[6] ? _GEN18964 : _GEN6840;
wire  _GEN18966 = io_x[41] ? _GEN18965 : _GEN6836;
wire  _GEN18967 = io_x[14] ? _GEN6843 : _GEN18966;
wire  _GEN18968 = io_x[0] ? _GEN6845 : _GEN18967;
wire  _GEN18969 = io_x[76] ? _GEN18968 : _GEN6834;
wire  _GEN18970 = io_x[42] ? _GEN18969 : _GEN6874;
wire  _GEN18971 = io_x[38] ? _GEN6871 : _GEN18970;
wire  _GEN18972 = io_x[10] ? _GEN18971 : _GEN18963;
wire  _GEN18973 = io_x[71] ? _GEN18972 : _GEN18946;
wire  _GEN18974 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN18975 = io_x[41] ? _GEN18974 : _GEN6836;
wire  _GEN18976 = io_x[14] ? _GEN18975 : _GEN6843;
wire  _GEN18977 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN18978 = io_x[14] ? _GEN6843 : _GEN18977;
wire  _GEN18979 = io_x[0] ? _GEN18978 : _GEN18976;
wire  _GEN18980 = io_x[76] ? _GEN18979 : _GEN6834;
wire  _GEN18981 = io_x[42] ? _GEN6874 : _GEN18980;
wire  _GEN18982 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN18983 = io_x[42] ? _GEN6874 : _GEN18982;
wire  _GEN18984 = io_x[38] ? _GEN18983 : _GEN18981;
wire  _GEN18985 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN18986 = io_x[0] ? _GEN6845 : _GEN18985;
wire  _GEN18987 = io_x[76] ? _GEN18986 : _GEN6834;
wire  _GEN18988 = io_x[42] ? _GEN6874 : _GEN18987;
wire  _GEN18989 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN18990 = io_x[38] ? _GEN18989 : _GEN18988;
wire  _GEN18991 = io_x[10] ? _GEN18990 : _GEN18984;
wire  _GEN18992 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN18993 = io_x[6] ? _GEN6850 : _GEN18992;
wire  _GEN18994 = io_x[41] ? _GEN6836 : _GEN18993;
wire  _GEN18995 = io_x[14] ? _GEN18994 : _GEN6856;
wire  _GEN18996 = io_x[0] ? _GEN6845 : _GEN18995;
wire  _GEN18997 = io_x[76] ? _GEN18996 : _GEN6834;
wire  _GEN18998 = io_x[42] ? _GEN6874 : _GEN18997;
wire  _GEN18999 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19000 = io_x[41] ? _GEN18999 : _GEN6836;
wire  _GEN19001 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19002 = io_x[41] ? _GEN19001 : _GEN6836;
wire  _GEN19003 = io_x[14] ? _GEN19002 : _GEN19000;
wire  _GEN19004 = io_x[0] ? _GEN6845 : _GEN19003;
wire  _GEN19005 = io_x[76] ? _GEN19004 : _GEN6834;
wire  _GEN19006 = io_x[42] ? _GEN19005 : _GEN6874;
wire  _GEN19007 = io_x[38] ? _GEN19006 : _GEN18998;
wire  _GEN19008 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19009 = io_x[0] ? _GEN6845 : _GEN19008;
wire  _GEN19010 = io_x[76] ? _GEN19009 : _GEN6834;
wire  _GEN19011 = io_x[42] ? _GEN6874 : _GEN19010;
wire  _GEN19012 = io_x[38] ? _GEN6871 : _GEN19011;
wire  _GEN19013 = io_x[10] ? _GEN19012 : _GEN19007;
wire  _GEN19014 = io_x[71] ? _GEN19013 : _GEN18991;
wire  _GEN19015 = io_x[70] ? _GEN19014 : _GEN18973;
wire  _GEN19016 = io_x[33] ? _GEN12627 : _GEN19015;
wire  _GEN19017 = io_x[21] ? _GEN19016 : _GEN18938;
wire  _GEN19018 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19019 = io_x[38] ? _GEN19018 : _GEN6871;
wire  _GEN19020 = io_x[10] ? _GEN7094 : _GEN19019;
wire  _GEN19021 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19022 = io_x[0] ? _GEN6845 : _GEN19021;
wire  _GEN19023 = io_x[76] ? _GEN19022 : _GEN6833;
wire  _GEN19024 = io_x[42] ? _GEN19023 : _GEN6874;
wire  _GEN19025 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19026 = io_x[41] ? _GEN19025 : _GEN6836;
wire  _GEN19027 = io_x[14] ? _GEN6856 : _GEN19026;
wire  _GEN19028 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19029 = io_x[41] ? _GEN19028 : _GEN6836;
wire  _GEN19030 = io_x[14] ? _GEN6843 : _GEN19029;
wire  _GEN19031 = io_x[0] ? _GEN19030 : _GEN19027;
wire  _GEN19032 = io_x[76] ? _GEN19031 : _GEN6833;
wire  _GEN19033 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN19034 = io_x[6] ? _GEN6850 : _GEN19033;
wire  _GEN19035 = io_x[41] ? _GEN19034 : _GEN6836;
wire  _GEN19036 = io_x[14] ? _GEN6843 : _GEN19035;
wire  _GEN19037 = io_x[0] ? _GEN6845 : _GEN19036;
wire  _GEN19038 = io_x[76] ? _GEN19037 : _GEN6834;
wire  _GEN19039 = io_x[42] ? _GEN19038 : _GEN19032;
wire  _GEN19040 = io_x[38] ? _GEN19039 : _GEN19024;
wire  _GEN19041 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19042 = io_x[0] ? _GEN6845 : _GEN19041;
wire  _GEN19043 = io_x[76] ? _GEN19042 : _GEN6834;
wire  _GEN19044 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19045 = io_x[0] ? _GEN19044 : _GEN6845;
wire  _GEN19046 = io_x[76] ? _GEN19045 : _GEN6833;
wire  _GEN19047 = io_x[42] ? _GEN19046 : _GEN19043;
wire  _GEN19048 = io_x[38] ? _GEN19047 : _GEN7036;
wire  _GEN19049 = io_x[10] ? _GEN19048 : _GEN19040;
wire  _GEN19050 = io_x[71] ? _GEN19049 : _GEN19020;
wire  _GEN19051 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN19052 = io_x[6] ? _GEN6850 : _GEN19051;
wire  _GEN19053 = io_x[41] ? _GEN19052 : _GEN6836;
wire  _GEN19054 = io_x[14] ? _GEN6843 : _GEN19053;
wire  _GEN19055 = io_x[0] ? _GEN19054 : _GEN6845;
wire  _GEN19056 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19057 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19058 = io_x[41] ? _GEN19057 : _GEN19056;
wire  _GEN19059 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19060 = io_x[41] ? _GEN6836 : _GEN19059;
wire  _GEN19061 = io_x[14] ? _GEN19060 : _GEN19058;
wire  _GEN19062 = io_x[0] ? _GEN19061 : _GEN6845;
wire  _GEN19063 = io_x[76] ? _GEN19062 : _GEN19055;
wire  _GEN19064 = io_x[42] ? _GEN6874 : _GEN19063;
wire  _GEN19065 = io_x[38] ? _GEN7036 : _GEN19064;
wire  _GEN19066 = io_x[10] ? _GEN7044 : _GEN19065;
wire  _GEN19067 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19068 = io_x[41] ? _GEN19067 : _GEN6836;
wire  _GEN19069 = io_x[14] ? _GEN6843 : _GEN19068;
wire  _GEN19070 = io_x[0] ? _GEN19069 : _GEN6845;
wire  _GEN19071 = io_x[76] ? _GEN19070 : _GEN6834;
wire  _GEN19072 = io_x[42] ? _GEN6874 : _GEN19071;
wire  _GEN19073 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN19074 = io_x[6] ? _GEN6850 : _GEN19073;
wire  _GEN19075 = io_x[41] ? _GEN19074 : _GEN6836;
wire  _GEN19076 = io_x[14] ? _GEN6856 : _GEN19075;
wire  _GEN19077 = io_x[0] ? _GEN19076 : _GEN6845;
wire  _GEN19078 = io_x[76] ? _GEN6834 : _GEN19077;
wire  _GEN19079 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19080 = io_x[41] ? _GEN19079 : _GEN6836;
wire  _GEN19081 = io_x[14] ? _GEN6856 : _GEN19080;
wire  _GEN19082 = io_x[0] ? _GEN19081 : _GEN6845;
wire  _GEN19083 = io_x[76] ? _GEN19082 : _GEN6833;
wire  _GEN19084 = io_x[42] ? _GEN19083 : _GEN19078;
wire  _GEN19085 = io_x[38] ? _GEN19084 : _GEN19072;
wire  _GEN19086 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19087 = io_x[41] ? _GEN6836 : _GEN19086;
wire  _GEN19088 = io_x[14] ? _GEN6843 : _GEN19087;
wire  _GEN19089 = io_x[0] ? _GEN6845 : _GEN19088;
wire  _GEN19090 = io_x[76] ? _GEN19089 : _GEN6834;
wire  _GEN19091 = io_x[42] ? _GEN6874 : _GEN19090;
wire  _GEN19092 = io_x[38] ? _GEN6871 : _GEN19091;
wire  _GEN19093 = io_x[10] ? _GEN19092 : _GEN19085;
wire  _GEN19094 = io_x[71] ? _GEN19093 : _GEN19066;
wire  _GEN19095 = io_x[70] ? _GEN19094 : _GEN19050;
wire  _GEN19096 = io_x[70] ? _GEN7020 : _GEN8474;
wire  _GEN19097 = io_x[33] ? _GEN19096 : _GEN19095;
wire  _GEN19098 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19099 = io_x[0] ? _GEN19098 : _GEN6845;
wire  _GEN19100 = io_x[76] ? _GEN19099 : _GEN6834;
wire  _GEN19101 = io_x[42] ? _GEN19100 : _GEN6874;
wire  _GEN19102 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19103 = io_x[0] ? _GEN19102 : _GEN6845;
wire  _GEN19104 = io_x[76] ? _GEN6833 : _GEN19103;
wire  _GEN19105 = io_x[42] ? _GEN6874 : _GEN19104;
wire  _GEN19106 = io_x[38] ? _GEN19105 : _GEN19101;
wire  _GEN19107 = io_x[10] ? _GEN7044 : _GEN19106;
wire  _GEN19108 = io_x[71] ? _GEN19107 : _GEN7203;
wire  _GEN19109 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19110 = io_x[0] ? _GEN19109 : _GEN6845;
wire  _GEN19111 = io_x[76] ? _GEN19110 : _GEN6834;
wire  _GEN19112 = io_x[42] ? _GEN6874 : _GEN19111;
wire  _GEN19113 = io_x[38] ? _GEN7036 : _GEN19112;
wire  _GEN19114 = io_x[10] ? _GEN7094 : _GEN19113;
wire  _GEN19115 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN19116 = io_x[42] ? _GEN19115 : _GEN6874;
wire  _GEN19117 = io_x[38] ? _GEN6871 : _GEN19116;
wire  _GEN19118 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19119 = io_x[0] ? _GEN6845 : _GEN19118;
wire  _GEN19120 = io_x[76] ? _GEN6834 : _GEN19119;
wire  _GEN19121 = io_x[42] ? _GEN6874 : _GEN19120;
wire  _GEN19122 = io_x[38] ? _GEN19121 : _GEN6871;
wire  _GEN19123 = io_x[10] ? _GEN19122 : _GEN19117;
wire  _GEN19124 = io_x[71] ? _GEN19123 : _GEN19114;
wire  _GEN19125 = io_x[70] ? _GEN19124 : _GEN19108;
wire  _GEN19126 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19127 = io_x[0] ? _GEN19126 : _GEN6845;
wire  _GEN19128 = io_x[76] ? _GEN19127 : _GEN6834;
wire  _GEN19129 = io_x[42] ? _GEN19128 : _GEN6874;
wire  _GEN19130 = io_x[38] ? _GEN6871 : _GEN19129;
wire  _GEN19131 = io_x[10] ? _GEN7044 : _GEN19130;
wire  _GEN19132 = io_x[71] ? _GEN19131 : _GEN7196;
wire  _GEN19133 = io_x[70] ? _GEN8474 : _GEN19132;
wire  _GEN19134 = io_x[33] ? _GEN19133 : _GEN19125;
wire  _GEN19135 = io_x[21] ? _GEN19134 : _GEN19097;
wire  _GEN19136 = io_x[18] ? _GEN19135 : _GEN19017;
wire  _GEN19137 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN19138 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19139 = io_x[0] ? _GEN6845 : _GEN19138;
wire  _GEN19140 = io_x[76] ? _GEN19139 : _GEN6834;
wire  _GEN19141 = io_x[42] ? _GEN19140 : _GEN6874;
wire  _GEN19142 = io_x[38] ? _GEN19141 : _GEN6871;
wire  _GEN19143 = io_x[10] ? _GEN19142 : _GEN19137;
wire  _GEN19144 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN19145 = io_x[76] ? _GEN19144 : _GEN6834;
wire  _GEN19146 = io_x[42] ? _GEN19145 : _GEN6874;
wire  _GEN19147 = io_x[38] ? _GEN19146 : _GEN6871;
wire  _GEN19148 = io_x[10] ? _GEN7044 : _GEN19147;
wire  _GEN19149 = io_x[71] ? _GEN19148 : _GEN19143;
wire  _GEN19150 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19151 = io_x[0] ? _GEN6858 : _GEN19150;
wire  _GEN19152 = io_x[76] ? _GEN19151 : _GEN6834;
wire  _GEN19153 = io_x[42] ? _GEN6874 : _GEN19152;
wire  _GEN19154 = io_x[38] ? _GEN6871 : _GEN19153;
wire  _GEN19155 = io_x[10] ? _GEN19154 : _GEN7044;
wire  _GEN19156 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19157 = io_x[41] ? _GEN6836 : _GEN19156;
wire  _GEN19158 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19159 = io_x[41] ? _GEN6836 : _GEN19158;
wire  _GEN19160 = io_x[14] ? _GEN19159 : _GEN19157;
wire  _GEN19161 = io_x[0] ? _GEN19160 : _GEN6845;
wire  _GEN19162 = io_x[76] ? _GEN19161 : _GEN6834;
wire  _GEN19163 = io_x[42] ? _GEN6874 : _GEN19162;
wire  _GEN19164 = io_x[38] ? _GEN6871 : _GEN19163;
wire  _GEN19165 = io_x[10] ? _GEN7094 : _GEN19164;
wire  _GEN19166 = io_x[71] ? _GEN19165 : _GEN19155;
wire  _GEN19167 = io_x[70] ? _GEN19166 : _GEN19149;
wire  _GEN19168 = io_x[33] ? _GEN12627 : _GEN19167;
wire  _GEN19169 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN19170 = io_x[76] ? _GEN19169 : _GEN6833;
wire  _GEN19171 = io_x[42] ? _GEN19170 : _GEN6863;
wire  _GEN19172 = io_x[38] ? _GEN19171 : _GEN6871;
wire  _GEN19173 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN19174 = io_x[76] ? _GEN19173 : _GEN6833;
wire  _GEN19175 = io_x[42] ? _GEN19174 : _GEN6874;
wire  _GEN19176 = io_x[38] ? _GEN19175 : _GEN6871;
wire  _GEN19177 = io_x[10] ? _GEN19176 : _GEN19172;
wire  _GEN19178 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19179 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19180 = io_x[41] ? _GEN19179 : _GEN6836;
wire  _GEN19181 = io_x[14] ? _GEN6843 : _GEN19180;
wire  _GEN19182 = io_x[0] ? _GEN6858 : _GEN19181;
wire  _GEN19183 = io_x[76] ? _GEN19182 : _GEN6834;
wire  _GEN19184 = io_x[42] ? _GEN19183 : _GEN6874;
wire  _GEN19185 = io_x[38] ? _GEN19184 : _GEN19178;
wire  _GEN19186 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19187 = io_x[41] ? _GEN6836 : _GEN19186;
wire  _GEN19188 = io_x[14] ? _GEN6856 : _GEN19187;
wire  _GEN19189 = io_x[0] ? _GEN19188 : _GEN6845;
wire  _GEN19190 = io_x[76] ? _GEN19189 : _GEN6834;
wire  _GEN19191 = io_x[42] ? _GEN19190 : _GEN6874;
wire  _GEN19192 = io_x[38] ? _GEN19191 : _GEN6871;
wire  _GEN19193 = io_x[10] ? _GEN19192 : _GEN19185;
wire  _GEN19194 = io_x[71] ? _GEN19193 : _GEN19177;
wire  _GEN19195 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19196 = io_x[0] ? _GEN19195 : _GEN6845;
wire  _GEN19197 = io_x[76] ? _GEN19196 : _GEN6834;
wire  _GEN19198 = io_x[42] ? _GEN6874 : _GEN19197;
wire  _GEN19199 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19200 = io_x[41] ? _GEN19199 : _GEN6836;
wire  _GEN19201 = io_x[14] ? _GEN6843 : _GEN19200;
wire  _GEN19202 = io_x[0] ? _GEN19201 : _GEN6845;
wire  _GEN19203 = io_x[76] ? _GEN19202 : _GEN6834;
wire  _GEN19204 = io_x[42] ? _GEN6863 : _GEN19203;
wire  _GEN19205 = io_x[38] ? _GEN19204 : _GEN19198;
wire  _GEN19206 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19207 = io_x[41] ? _GEN6924 : _GEN19206;
wire  _GEN19208 = io_x[14] ? _GEN19207 : _GEN6843;
wire  _GEN19209 = io_x[0] ? _GEN6858 : _GEN19208;
wire  _GEN19210 = io_x[76] ? _GEN6834 : _GEN19209;
wire  _GEN19211 = io_x[42] ? _GEN19210 : _GEN6874;
wire  _GEN19212 = io_x[38] ? _GEN6871 : _GEN19211;
wire  _GEN19213 = io_x[10] ? _GEN19212 : _GEN19205;
wire  _GEN19214 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19215 = io_x[0] ? _GEN19214 : _GEN6845;
wire  _GEN19216 = io_x[76] ? _GEN19215 : _GEN6833;
wire  _GEN19217 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19218 = io_x[41] ? _GEN6836 : _GEN19217;
wire  _GEN19219 = io_x[14] ? _GEN6843 : _GEN19218;
wire  _GEN19220 = io_x[0] ? _GEN6845 : _GEN19219;
wire  _GEN19221 = io_x[76] ? _GEN19220 : _GEN6833;
wire  _GEN19222 = io_x[42] ? _GEN19221 : _GEN19216;
wire  _GEN19223 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19224 = io_x[0] ? _GEN19223 : _GEN6845;
wire  _GEN19225 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN19226 = io_x[76] ? _GEN19225 : _GEN19224;
wire  _GEN19227 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN19228 = io_x[6] ? _GEN6850 : _GEN19227;
wire  _GEN19229 = io_x[41] ? _GEN19228 : _GEN6836;
wire  _GEN19230 = io_x[14] ? _GEN6856 : _GEN19229;
wire  _GEN19231 = io_x[0] ? _GEN6858 : _GEN19230;
wire  _GEN19232 = io_x[76] ? _GEN19231 : _GEN6834;
wire  _GEN19233 = io_x[42] ? _GEN19232 : _GEN19226;
wire  _GEN19234 = io_x[38] ? _GEN19233 : _GEN19222;
wire  _GEN19235 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN19236 = io_x[42] ? _GEN19235 : _GEN6874;
wire  _GEN19237 = io_x[38] ? _GEN7036 : _GEN19236;
wire  _GEN19238 = io_x[10] ? _GEN19237 : _GEN19234;
wire  _GEN19239 = io_x[71] ? _GEN19238 : _GEN19213;
wire  _GEN19240 = io_x[70] ? _GEN19239 : _GEN19194;
wire  _GEN19241 = io_x[33] ? _GEN12627 : _GEN19240;
wire  _GEN19242 = io_x[21] ? _GEN19241 : _GEN19168;
wire  _GEN19243 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19244 = io_x[38] ? _GEN19243 : _GEN6871;
wire  _GEN19245 = io_x[10] ? _GEN7044 : _GEN19244;
wire  _GEN19246 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19247 = io_x[41] ? _GEN6836 : _GEN19246;
wire  _GEN19248 = io_x[14] ? _GEN6843 : _GEN19247;
wire  _GEN19249 = io_x[0] ? _GEN19248 : _GEN6845;
wire  _GEN19250 = io_x[76] ? _GEN19249 : _GEN6833;
wire  _GEN19251 = io_x[42] ? _GEN19250 : _GEN6874;
wire  _GEN19252 = io_x[38] ? _GEN6871 : _GEN19251;
wire  _GEN19253 = io_x[10] ? _GEN7044 : _GEN19252;
wire  _GEN19254 = io_x[71] ? _GEN19253 : _GEN19245;
wire  _GEN19255 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19256 = io_x[41] ? _GEN6836 : _GEN19255;
wire  _GEN19257 = io_x[14] ? _GEN6843 : _GEN19256;
wire  _GEN19258 = io_x[0] ? _GEN6845 : _GEN19257;
wire  _GEN19259 = io_x[76] ? _GEN19258 : _GEN6834;
wire  _GEN19260 = io_x[42] ? _GEN6874 : _GEN19259;
wire  _GEN19261 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN19262 = io_x[42] ? _GEN6874 : _GEN19261;
wire  _GEN19263 = io_x[38] ? _GEN19262 : _GEN19260;
wire  _GEN19264 = io_x[10] ? _GEN7044 : _GEN19263;
wire  _GEN19265 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN19266 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19267 = io_x[41] ? _GEN6836 : _GEN19266;
wire  _GEN19268 = io_x[14] ? _GEN6843 : _GEN19267;
wire  _GEN19269 = io_x[0] ? _GEN19268 : _GEN6845;
wire  _GEN19270 = io_x[76] ? _GEN19269 : _GEN6834;
wire  _GEN19271 = io_x[42] ? _GEN19270 : _GEN19265;
wire  _GEN19272 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN19273 = io_x[14] ? _GEN6843 : _GEN19272;
wire  _GEN19274 = io_x[0] ? _GEN19273 : _GEN6845;
wire  _GEN19275 = io_x[76] ? _GEN19274 : _GEN6834;
wire  _GEN19276 = io_x[42] ? _GEN19275 : _GEN6874;
wire  _GEN19277 = io_x[38] ? _GEN19276 : _GEN19271;
wire  _GEN19278 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19279 = io_x[0] ? _GEN6845 : _GEN19278;
wire  _GEN19280 = io_x[76] ? _GEN19279 : _GEN6834;
wire  _GEN19281 = io_x[42] ? _GEN6874 : _GEN19280;
wire  _GEN19282 = io_x[38] ? _GEN6871 : _GEN19281;
wire  _GEN19283 = io_x[10] ? _GEN19282 : _GEN19277;
wire  _GEN19284 = io_x[71] ? _GEN19283 : _GEN19264;
wire  _GEN19285 = io_x[70] ? _GEN19284 : _GEN19254;
wire  _GEN19286 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19287 = io_x[41] ? _GEN6836 : _GEN19286;
wire  _GEN19288 = io_x[14] ? _GEN6843 : _GEN19287;
wire  _GEN19289 = io_x[0] ? _GEN19288 : _GEN6845;
wire  _GEN19290 = io_x[76] ? _GEN19289 : _GEN6834;
wire  _GEN19291 = io_x[42] ? _GEN19290 : _GEN6874;
wire  _GEN19292 = io_x[38] ? _GEN6871 : _GEN19291;
wire  _GEN19293 = io_x[10] ? _GEN7044 : _GEN19292;
wire  _GEN19294 = io_x[71] ? _GEN19293 : _GEN7196;
wire  _GEN19295 = io_x[70] ? _GEN8474 : _GEN19294;
wire  _GEN19296 = io_x[33] ? _GEN19295 : _GEN19285;
wire  _GEN19297 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19298 = io_x[41] ? _GEN19297 : _GEN6836;
wire  _GEN19299 = io_x[14] ? _GEN19298 : _GEN6856;
wire  _GEN19300 = io_x[0] ? _GEN19299 : _GEN6845;
wire  _GEN19301 = io_x[76] ? _GEN6834 : _GEN19300;
wire  _GEN19302 = io_x[42] ? _GEN6863 : _GEN19301;
wire  _GEN19303 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19304 = io_x[41] ? _GEN19303 : _GEN6836;
wire  _GEN19305 = io_x[14] ? _GEN6843 : _GEN19304;
wire  _GEN19306 = io_x[0] ? _GEN6845 : _GEN19305;
wire  _GEN19307 = io_x[76] ? _GEN6834 : _GEN19306;
wire  _GEN19308 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19309 = io_x[0] ? _GEN6845 : _GEN19308;
wire  _GEN19310 = io_x[76] ? _GEN19309 : _GEN6834;
wire  _GEN19311 = io_x[42] ? _GEN19310 : _GEN19307;
wire  _GEN19312 = io_x[38] ? _GEN19311 : _GEN19302;
wire  _GEN19313 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19314 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN19315 = io_x[14] ? _GEN19314 : _GEN6843;
wire  _GEN19316 = io_x[0] ? _GEN19315 : _GEN6845;
wire  _GEN19317 = io_x[76] ? _GEN19316 : _GEN6834;
wire  _GEN19318 = io_x[42] ? _GEN19317 : _GEN6874;
wire  _GEN19319 = io_x[38] ? _GEN19318 : _GEN19313;
wire  _GEN19320 = io_x[10] ? _GEN19319 : _GEN19312;
wire  _GEN19321 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19322 = io_x[41] ? _GEN6836 : _GEN19321;
wire  _GEN19323 = io_x[14] ? _GEN6843 : _GEN19322;
wire  _GEN19324 = io_x[0] ? _GEN19323 : _GEN6858;
wire  _GEN19325 = io_x[76] ? _GEN19324 : _GEN6834;
wire  _GEN19326 = io_x[42] ? _GEN19325 : _GEN6863;
wire  _GEN19327 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19328 = io_x[41] ? _GEN19327 : _GEN6836;
wire  _GEN19329 = io_x[14] ? _GEN6856 : _GEN19328;
wire  _GEN19330 = io_x[0] ? _GEN19329 : _GEN6845;
wire  _GEN19331 = io_x[76] ? _GEN19330 : _GEN6834;
wire  _GEN19332 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN19333 = io_x[76] ? _GEN19332 : _GEN6834;
wire  _GEN19334 = io_x[42] ? _GEN19333 : _GEN19331;
wire  _GEN19335 = io_x[38] ? _GEN19334 : _GEN19326;
wire  _GEN19336 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN19337 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN19338 = io_x[42] ? _GEN19337 : _GEN19336;
wire  _GEN19339 = io_x[38] ? _GEN19338 : _GEN6871;
wire  _GEN19340 = io_x[10] ? _GEN19339 : _GEN19335;
wire  _GEN19341 = io_x[71] ? _GEN19340 : _GEN19320;
wire  _GEN19342 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN19343 = io_x[6] ? _GEN6850 : _GEN19342;
wire  _GEN19344 = io_x[41] ? _GEN19343 : _GEN6836;
wire  _GEN19345 = io_x[14] ? _GEN6843 : _GEN19344;
wire  _GEN19346 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19347 = io_x[41] ? _GEN19346 : _GEN6836;
wire  _GEN19348 = io_x[14] ? _GEN6843 : _GEN19347;
wire  _GEN19349 = io_x[0] ? _GEN19348 : _GEN19345;
wire  _GEN19350 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN19351 = io_x[76] ? _GEN19350 : _GEN19349;
wire  _GEN19352 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN19353 = io_x[14] ? _GEN6843 : _GEN19352;
wire  _GEN19354 = io_x[0] ? _GEN6858 : _GEN19353;
wire  _GEN19355 = io_x[76] ? _GEN6834 : _GEN19354;
wire  _GEN19356 = io_x[42] ? _GEN19355 : _GEN19351;
wire  _GEN19357 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN19358 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19359 = io_x[0] ? _GEN6845 : _GEN19358;
wire  _GEN19360 = io_x[76] ? _GEN19359 : _GEN19357;
wire  _GEN19361 = io_x[42] ? _GEN19360 : _GEN6874;
wire  _GEN19362 = io_x[38] ? _GEN19361 : _GEN19356;
wire  _GEN19363 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19364 = io_x[0] ? _GEN6845 : _GEN19363;
wire  _GEN19365 = io_x[76] ? _GEN6834 : _GEN19364;
wire  _GEN19366 = io_x[42] ? _GEN6863 : _GEN19365;
wire  _GEN19367 = io_x[38] ? _GEN7036 : _GEN19366;
wire  _GEN19368 = io_x[10] ? _GEN19367 : _GEN19362;
wire  _GEN19369 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19370 = io_x[41] ? _GEN19369 : _GEN6836;
wire  _GEN19371 = io_x[14] ? _GEN6856 : _GEN19370;
wire  _GEN19372 = io_x[0] ? _GEN19371 : _GEN6845;
wire  _GEN19373 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN19374 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19375 = io_x[41] ? _GEN6836 : _GEN19374;
wire  _GEN19376 = io_x[14] ? _GEN19375 : _GEN19373;
wire  _GEN19377 = io_x[0] ? _GEN19376 : _GEN6845;
wire  _GEN19378 = io_x[76] ? _GEN19377 : _GEN19372;
wire  _GEN19379 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN19380 = io_x[14] ? _GEN6843 : _GEN19379;
wire  _GEN19381 = io_x[0] ? _GEN6845 : _GEN19380;
wire  _GEN19382 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN19383 = io_x[14] ? _GEN6843 : _GEN19382;
wire  _GEN19384 = io_x[0] ? _GEN6845 : _GEN19383;
wire  _GEN19385 = io_x[76] ? _GEN19384 : _GEN19381;
wire  _GEN19386 = io_x[42] ? _GEN19385 : _GEN19378;
wire  _GEN19387 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19388 = io_x[41] ? _GEN6836 : _GEN19387;
wire  _GEN19389 = io_x[14] ? _GEN6843 : _GEN19388;
wire  _GEN19390 = io_x[0] ? _GEN19389 : _GEN6858;
wire  _GEN19391 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN19392 = io_x[14] ? _GEN6843 : _GEN19391;
wire  _GEN19393 = io_x[0] ? _GEN6845 : _GEN19392;
wire  _GEN19394 = io_x[76] ? _GEN19393 : _GEN19390;
wire  _GEN19395 = io_x[42] ? _GEN19394 : _GEN6874;
wire  _GEN19396 = io_x[38] ? _GEN19395 : _GEN19386;
wire  _GEN19397 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN19398 = io_x[14] ? _GEN19397 : _GEN6843;
wire  _GEN19399 = io_x[0] ? _GEN19398 : _GEN6845;
wire  _GEN19400 = io_x[76] ? _GEN19399 : _GEN6833;
wire  _GEN19401 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19402 = io_x[0] ? _GEN6845 : _GEN19401;
wire  _GEN19403 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19404 = io_x[0] ? _GEN6845 : _GEN19403;
wire  _GEN19405 = io_x[76] ? _GEN19404 : _GEN19402;
wire  _GEN19406 = io_x[42] ? _GEN19405 : _GEN19400;
wire  _GEN19407 = io_x[38] ? _GEN7036 : _GEN19406;
wire  _GEN19408 = io_x[10] ? _GEN19407 : _GEN19396;
wire  _GEN19409 = io_x[71] ? _GEN19408 : _GEN19368;
wire  _GEN19410 = io_x[70] ? _GEN19409 : _GEN19341;
wire  _GEN19411 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN19412 = io_x[10] ? _GEN7044 : _GEN19411;
wire  _GEN19413 = io_x[71] ? _GEN19412 : _GEN7196;
wire  _GEN19414 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN19415 = io_x[71] ? _GEN7196 : _GEN19414;
wire  _GEN19416 = io_x[70] ? _GEN19415 : _GEN19413;
wire  _GEN19417 = io_x[33] ? _GEN19416 : _GEN19410;
wire  _GEN19418 = io_x[21] ? _GEN19417 : _GEN19296;
wire  _GEN19419 = io_x[18] ? _GEN19418 : _GEN19242;
wire  _GEN19420 = io_x[20] ? _GEN19419 : _GEN19136;
wire  _GEN19421 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN19422 = io_x[76] ? _GEN6834 : _GEN19421;
wire  _GEN19423 = io_x[42] ? _GEN19422 : _GEN6863;
wire  _GEN19424 = io_x[38] ? _GEN7036 : _GEN19423;
wire  _GEN19425 = io_x[10] ? _GEN7044 : _GEN19424;
wire  _GEN19426 = io_x[71] ? _GEN19425 : _GEN7203;
wire  _GEN19427 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN19428 = io_x[10] ? _GEN7094 : _GEN19427;
wire  _GEN19429 = io_x[71] ? _GEN7196 : _GEN19428;
wire  _GEN19430 = io_x[70] ? _GEN19429 : _GEN19426;
wire  _GEN19431 = io_x[33] ? _GEN12627 : _GEN19430;
wire  _GEN19432 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19433 = io_x[41] ? _GEN6836 : _GEN19432;
wire  _GEN19434 = io_x[14] ? _GEN19433 : _GEN6843;
wire  _GEN19435 = io_x[0] ? _GEN19434 : _GEN6845;
wire  _GEN19436 = io_x[76] ? _GEN19435 : _GEN6834;
wire  _GEN19437 = io_x[42] ? _GEN6874 : _GEN19436;
wire  _GEN19438 = io_x[38] ? _GEN19437 : _GEN6871;
wire  _GEN19439 = io_x[10] ? _GEN19438 : _GEN7094;
wire  _GEN19440 = io_x[71] ? _GEN19439 : _GEN7196;
wire  _GEN19441 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN19442 = io_x[71] ? _GEN19441 : _GEN7203;
wire  _GEN19443 = io_x[70] ? _GEN19442 : _GEN19440;
wire  _GEN19444 = io_x[33] ? _GEN12627 : _GEN19443;
wire  _GEN19445 = io_x[21] ? _GEN19444 : _GEN19431;
wire  _GEN19446 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN19447 = io_x[42] ? _GEN6874 : _GEN19446;
wire  _GEN19448 = io_x[38] ? _GEN6871 : _GEN19447;
wire  _GEN19449 = io_x[10] ? _GEN7044 : _GEN19448;
wire  _GEN19450 = io_x[71] ? _GEN19449 : _GEN7196;
wire  _GEN19451 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN19452 = io_x[71] ? _GEN19451 : _GEN7203;
wire  _GEN19453 = io_x[70] ? _GEN19452 : _GEN19450;
wire  _GEN19454 = io_x[33] ? _GEN12641 : _GEN19453;
wire  _GEN19455 = io_x[21] ? _GEN19454 : _GEN12643;
wire  _GEN19456 = io_x[18] ? _GEN19455 : _GEN19445;
wire  _GEN19457 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19458 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN19459 = io_x[76] ? _GEN6834 : _GEN19458;
wire  _GEN19460 = io_x[42] ? _GEN19459 : _GEN6874;
wire  _GEN19461 = io_x[38] ? _GEN19460 : _GEN19457;
wire  _GEN19462 = io_x[10] ? _GEN7094 : _GEN19461;
wire  _GEN19463 = io_x[71] ? _GEN7196 : _GEN19462;
wire  _GEN19464 = io_x[70] ? _GEN19463 : _GEN8474;
wire  _GEN19465 = io_x[33] ? _GEN12641 : _GEN19464;
wire  _GEN19466 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN19467 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19468 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN19469 = io_x[38] ? _GEN19468 : _GEN19467;
wire  _GEN19470 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN19471 = io_x[42] ? _GEN6863 : _GEN19470;
wire  _GEN19472 = io_x[38] ? _GEN6871 : _GEN19471;
wire  _GEN19473 = io_x[10] ? _GEN19472 : _GEN19469;
wire  _GEN19474 = io_x[71] ? _GEN19473 : _GEN19466;
wire  _GEN19475 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN19476 = io_x[14] ? _GEN6843 : _GEN19475;
wire  _GEN19477 = io_x[0] ? _GEN6845 : _GEN19476;
wire  _GEN19478 = io_x[76] ? _GEN19477 : _GEN6834;
wire  _GEN19479 = io_x[42] ? _GEN6863 : _GEN19478;
wire  _GEN19480 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN19481 = io_x[38] ? _GEN19480 : _GEN19479;
wire  _GEN19482 = io_x[10] ? _GEN7094 : _GEN19481;
wire  _GEN19483 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN19484 = io_x[38] ? _GEN19483 : _GEN7036;
wire  _GEN19485 = io_x[10] ? _GEN7094 : _GEN19484;
wire  _GEN19486 = io_x[71] ? _GEN19485 : _GEN19482;
wire  _GEN19487 = io_x[70] ? _GEN19486 : _GEN19474;
wire  _GEN19488 = io_x[33] ? _GEN12627 : _GEN19487;
wire  _GEN19489 = io_x[21] ? _GEN19488 : _GEN19465;
wire  _GEN19490 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN19491 = io_x[42] ? _GEN6874 : _GEN19490;
wire  _GEN19492 = io_x[38] ? _GEN19491 : _GEN6871;
wire  _GEN19493 = io_x[10] ? _GEN7044 : _GEN19492;
wire  _GEN19494 = io_x[71] ? _GEN19493 : _GEN7203;
wire  _GEN19495 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN19496 = io_x[6] ? _GEN6850 : _GEN19495;
wire  _GEN19497 = io_x[41] ? _GEN6836 : _GEN19496;
wire  _GEN19498 = io_x[14] ? _GEN6843 : _GEN19497;
wire  _GEN19499 = io_x[0] ? _GEN6845 : _GEN19498;
wire  _GEN19500 = io_x[76] ? _GEN19499 : _GEN6834;
wire  _GEN19501 = io_x[42] ? _GEN6874 : _GEN19500;
wire  _GEN19502 = io_x[38] ? _GEN19501 : _GEN6871;
wire  _GEN19503 = io_x[10] ? _GEN7044 : _GEN19502;
wire  _GEN19504 = io_x[71] ? _GEN7196 : _GEN19503;
wire  _GEN19505 = io_x[70] ? _GEN19504 : _GEN19494;
wire  _GEN19506 = io_x[33] ? _GEN12627 : _GEN19505;
wire  _GEN19507 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN19508 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19509 = io_x[38] ? _GEN19508 : _GEN19507;
wire  _GEN19510 = io_x[10] ? _GEN7044 : _GEN19509;
wire  _GEN19511 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19512 = io_x[41] ? _GEN6836 : _GEN19511;
wire  _GEN19513 = io_x[14] ? _GEN19512 : _GEN6856;
wire  _GEN19514 = io_x[0] ? _GEN19513 : _GEN6858;
wire  _GEN19515 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19516 = io_x[41] ? _GEN6836 : _GEN19515;
wire  _GEN19517 = io_x[14] ? _GEN6856 : _GEN19516;
wire  _GEN19518 = io_x[0] ? _GEN19517 : _GEN6845;
wire  _GEN19519 = io_x[76] ? _GEN19518 : _GEN19514;
wire  _GEN19520 = io_x[42] ? _GEN6874 : _GEN19519;
wire  _GEN19521 = io_x[38] ? _GEN6871 : _GEN19520;
wire  _GEN19522 = io_x[10] ? _GEN7044 : _GEN19521;
wire  _GEN19523 = io_x[71] ? _GEN19522 : _GEN19510;
wire  _GEN19524 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19525 = io_x[41] ? _GEN6836 : _GEN19524;
wire  _GEN19526 = io_x[14] ? _GEN6856 : _GEN19525;
wire  _GEN19527 = io_x[0] ? _GEN19526 : _GEN6858;
wire  _GEN19528 = io_x[76] ? _GEN19527 : _GEN6834;
wire  _GEN19529 = io_x[42] ? _GEN6874 : _GEN19528;
wire  _GEN19530 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN19531 = io_x[76] ? _GEN19530 : _GEN6833;
wire  _GEN19532 = io_x[42] ? _GEN19531 : _GEN6874;
wire  _GEN19533 = io_x[38] ? _GEN19532 : _GEN19529;
wire  _GEN19534 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19535 = io_x[41] ? _GEN19534 : _GEN6836;
wire  _GEN19536 = io_x[14] ? _GEN19535 : _GEN6843;
wire  _GEN19537 = io_x[0] ? _GEN19536 : _GEN6845;
wire  _GEN19538 = io_x[76] ? _GEN6834 : _GEN19537;
wire  _GEN19539 = io_x[42] ? _GEN6874 : _GEN19538;
wire  _GEN19540 = io_x[38] ? _GEN7036 : _GEN19539;
wire  _GEN19541 = io_x[10] ? _GEN19540 : _GEN19533;
wire  _GEN19542 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19543 = io_x[41] ? _GEN19542 : _GEN6836;
wire  _GEN19544 = io_x[14] ? _GEN6843 : _GEN19543;
wire  _GEN19545 = io_x[0] ? _GEN19544 : _GEN6845;
wire  _GEN19546 = io_x[76] ? _GEN19545 : _GEN6833;
wire  _GEN19547 = io_x[42] ? _GEN6874 : _GEN19546;
wire  _GEN19548 = io_x[38] ? _GEN6871 : _GEN19547;
wire  _GEN19549 = io_x[10] ? _GEN7044 : _GEN19548;
wire  _GEN19550 = io_x[71] ? _GEN19549 : _GEN19541;
wire  _GEN19551 = io_x[70] ? _GEN19550 : _GEN19523;
wire  _GEN19552 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19553 = io_x[41] ? _GEN6836 : _GEN19552;
wire  _GEN19554 = io_x[14] ? _GEN19553 : _GEN6856;
wire  _GEN19555 = io_x[0] ? _GEN19554 : _GEN6845;
wire  _GEN19556 = io_x[76] ? _GEN6834 : _GEN19555;
wire  _GEN19557 = io_x[42] ? _GEN6874 : _GEN19556;
wire  _GEN19558 = io_x[38] ? _GEN6871 : _GEN19557;
wire  _GEN19559 = io_x[10] ? _GEN7044 : _GEN19558;
wire  _GEN19560 = io_x[71] ? _GEN19559 : _GEN7196;
wire  _GEN19561 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN19562 = io_x[10] ? _GEN7044 : _GEN19561;
wire  _GEN19563 = io_x[71] ? _GEN7196 : _GEN19562;
wire  _GEN19564 = io_x[70] ? _GEN19563 : _GEN19560;
wire  _GEN19565 = io_x[33] ? _GEN19564 : _GEN19551;
wire  _GEN19566 = io_x[21] ? _GEN19565 : _GEN19506;
wire  _GEN19567 = io_x[18] ? _GEN19566 : _GEN19489;
wire  _GEN19568 = io_x[20] ? _GEN19567 : _GEN19456;
wire  _GEN19569 = io_x[45] ? _GEN19568 : _GEN19420;
wire  _GEN19570 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19571 = io_x[0] ? _GEN6845 : _GEN19570;
wire  _GEN19572 = io_x[76] ? _GEN19571 : _GEN6834;
wire  _GEN19573 = io_x[42] ? _GEN19572 : _GEN6874;
wire  _GEN19574 = io_x[38] ? _GEN19573 : _GEN6871;
wire  _GEN19575 = io_x[10] ? _GEN19574 : _GEN7094;
wire  _GEN19576 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19577 = io_x[41] ? _GEN6836 : _GEN19576;
wire  _GEN19578 = io_x[14] ? _GEN19577 : _GEN6843;
wire  _GEN19579 = io_x[0] ? _GEN19578 : _GEN6845;
wire  _GEN19580 = io_x[76] ? _GEN19579 : _GEN6834;
wire  _GEN19581 = io_x[42] ? _GEN19580 : _GEN6874;
wire  _GEN19582 = io_x[38] ? _GEN19581 : _GEN6871;
wire  _GEN19583 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19584 = io_x[0] ? _GEN6845 : _GEN19583;
wire  _GEN19585 = io_x[76] ? _GEN19584 : _GEN6834;
wire  _GEN19586 = io_x[42] ? _GEN19585 : _GEN6874;
wire  _GEN19587 = io_x[38] ? _GEN6871 : _GEN19586;
wire  _GEN19588 = io_x[10] ? _GEN19587 : _GEN19582;
wire  _GEN19589 = io_x[71] ? _GEN19588 : _GEN19575;
wire  _GEN19590 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN19591 = io_x[14] ? _GEN6843 : _GEN19590;
wire  _GEN19592 = io_x[0] ? _GEN19591 : _GEN6858;
wire  _GEN19593 = io_x[76] ? _GEN19592 : _GEN6834;
wire  _GEN19594 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN19595 = io_x[42] ? _GEN19594 : _GEN19593;
wire  _GEN19596 = io_x[38] ? _GEN6871 : _GEN19595;
wire  _GEN19597 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN19598 = io_x[14] ? _GEN6843 : _GEN19597;
wire  _GEN19599 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN19600 = io_x[14] ? _GEN19599 : _GEN6843;
wire  _GEN19601 = io_x[0] ? _GEN19600 : _GEN19598;
wire  _GEN19602 = io_x[76] ? _GEN19601 : _GEN6834;
wire  _GEN19603 = io_x[42] ? _GEN6874 : _GEN19602;
wire  _GEN19604 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19605 = io_x[41] ? _GEN19604 : _GEN6836;
wire  _GEN19606 = io_x[14] ? _GEN6843 : _GEN19605;
wire  _GEN19607 = io_x[0] ? _GEN19606 : _GEN6845;
wire  _GEN19608 = io_x[76] ? _GEN19607 : _GEN6834;
wire  _GEN19609 = io_x[42] ? _GEN6874 : _GEN19608;
wire  _GEN19610 = io_x[38] ? _GEN19609 : _GEN19603;
wire  _GEN19611 = io_x[10] ? _GEN19610 : _GEN19596;
wire  _GEN19612 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19613 = io_x[0] ? _GEN6845 : _GEN19612;
wire  _GEN19614 = io_x[76] ? _GEN19613 : _GEN6834;
wire  _GEN19615 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN19616 = io_x[42] ? _GEN19615 : _GEN19614;
wire  _GEN19617 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19618 = io_x[41] ? _GEN6836 : _GEN19617;
wire  _GEN19619 = io_x[14] ? _GEN19618 : _GEN6843;
wire  _GEN19620 = io_x[0] ? _GEN19619 : _GEN6845;
wire  _GEN19621 = io_x[76] ? _GEN19620 : _GEN6834;
wire  _GEN19622 = io_x[42] ? _GEN19621 : _GEN6874;
wire  _GEN19623 = io_x[38] ? _GEN19622 : _GEN19616;
wire  _GEN19624 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19625 = io_x[41] ? _GEN19624 : _GEN6836;
wire  _GEN19626 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19627 = io_x[41] ? _GEN19626 : _GEN6836;
wire  _GEN19628 = io_x[14] ? _GEN19627 : _GEN19625;
wire  _GEN19629 = io_x[0] ? _GEN6845 : _GEN19628;
wire  _GEN19630 = io_x[76] ? _GEN19629 : _GEN6834;
wire  _GEN19631 = io_x[42] ? _GEN19630 : _GEN6874;
wire  _GEN19632 = io_x[38] ? _GEN19631 : _GEN7036;
wire  _GEN19633 = io_x[10] ? _GEN19632 : _GEN19623;
wire  _GEN19634 = io_x[71] ? _GEN19633 : _GEN19611;
wire  _GEN19635 = io_x[70] ? _GEN19634 : _GEN19589;
wire  _GEN19636 = io_x[33] ? _GEN12627 : _GEN19635;
wire  _GEN19637 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN19638 = io_x[6] ? _GEN19637 : _GEN6850;
wire  _GEN19639 = io_x[41] ? _GEN19638 : _GEN6836;
wire  _GEN19640 = io_x[14] ? _GEN19639 : _GEN6843;
wire  _GEN19641 = io_x[0] ? _GEN19640 : _GEN6845;
wire  _GEN19642 = io_x[76] ? _GEN6834 : _GEN19641;
wire  _GEN19643 = io_x[42] ? _GEN6874 : _GEN19642;
wire  _GEN19644 = io_x[38] ? _GEN19643 : _GEN7036;
wire  _GEN19645 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19646 = io_x[38] ? _GEN19645 : _GEN6871;
wire  _GEN19647 = io_x[10] ? _GEN19646 : _GEN19644;
wire  _GEN19648 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN19649 = io_x[42] ? _GEN19648 : _GEN6874;
wire  _GEN19650 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN19651 = io_x[76] ? _GEN19650 : _GEN6834;
wire  _GEN19652 = io_x[42] ? _GEN19651 : _GEN6874;
wire  _GEN19653 = io_x[38] ? _GEN19652 : _GEN19649;
wire  _GEN19654 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN19655 = io_x[6] ? _GEN6840 : _GEN19654;
wire  _GEN19656 = io_x[41] ? _GEN19655 : _GEN6836;
wire  _GEN19657 = io_x[14] ? _GEN6843 : _GEN19656;
wire  _GEN19658 = io_x[0] ? _GEN6845 : _GEN19657;
wire  _GEN19659 = io_x[76] ? _GEN19658 : _GEN6834;
wire  _GEN19660 = io_x[42] ? _GEN19659 : _GEN6874;
wire  _GEN19661 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN19662 = io_x[42] ? _GEN19661 : _GEN6874;
wire  _GEN19663 = io_x[38] ? _GEN19662 : _GEN19660;
wire  _GEN19664 = io_x[10] ? _GEN19663 : _GEN19653;
wire  _GEN19665 = io_x[71] ? _GEN19664 : _GEN19647;
wire  _GEN19666 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19667 = io_x[0] ? _GEN6845 : _GEN19666;
wire  _GEN19668 = io_x[76] ? _GEN19667 : _GEN6834;
wire  _GEN19669 = io_x[42] ? _GEN6874 : _GEN19668;
wire  _GEN19670 = io_x[38] ? _GEN7036 : _GEN19669;
wire  _GEN19671 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19672 = io_x[0] ? _GEN6845 : _GEN19671;
wire  _GEN19673 = io_x[76] ? _GEN19672 : _GEN6834;
wire  _GEN19674 = io_x[42] ? _GEN6863 : _GEN19673;
wire  _GEN19675 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN19676 = io_x[76] ? _GEN6834 : _GEN19675;
wire  _GEN19677 = io_x[42] ? _GEN6863 : _GEN19676;
wire  _GEN19678 = io_x[38] ? _GEN19677 : _GEN19674;
wire  _GEN19679 = io_x[10] ? _GEN19678 : _GEN19670;
wire  _GEN19680 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19681 = io_x[41] ? _GEN19680 : _GEN6836;
wire  _GEN19682 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19683 = io_x[41] ? _GEN19682 : _GEN6836;
wire  _GEN19684 = io_x[14] ? _GEN19683 : _GEN19681;
wire  _GEN19685 = io_x[0] ? _GEN6845 : _GEN19684;
wire  _GEN19686 = io_x[76] ? _GEN19685 : _GEN6834;
wire  _GEN19687 = io_x[42] ? _GEN19686 : _GEN6874;
wire  _GEN19688 = io_x[38] ? _GEN19687 : _GEN6871;
wire  _GEN19689 = io_x[10] ? _GEN19688 : _GEN7044;
wire  _GEN19690 = io_x[71] ? _GEN19689 : _GEN19679;
wire  _GEN19691 = io_x[70] ? _GEN19690 : _GEN19665;
wire  _GEN19692 = io_x[33] ? _GEN12627 : _GEN19691;
wire  _GEN19693 = io_x[21] ? _GEN19692 : _GEN19636;
wire  _GEN19694 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN19695 = io_x[42] ? _GEN19694 : _GEN6874;
wire  _GEN19696 = io_x[38] ? _GEN19695 : _GEN6871;
wire  _GEN19697 = io_x[10] ? _GEN19696 : _GEN7044;
wire  _GEN19698 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19699 = io_x[41] ? _GEN19698 : _GEN6836;
wire  _GEN19700 = io_x[14] ? _GEN6856 : _GEN19699;
wire  _GEN19701 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19702 = io_x[0] ? _GEN19701 : _GEN19700;
wire  _GEN19703 = io_x[76] ? _GEN19702 : _GEN6834;
wire  _GEN19704 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19705 = io_x[41] ? _GEN6836 : _GEN19704;
wire  _GEN19706 = io_x[14] ? _GEN19705 : _GEN6843;
wire  _GEN19707 = io_x[0] ? _GEN19706 : _GEN6845;
wire  _GEN19708 = io_x[76] ? _GEN6834 : _GEN19707;
wire  _GEN19709 = io_x[42] ? _GEN19708 : _GEN19703;
wire  _GEN19710 = io_x[38] ? _GEN19709 : _GEN6871;
wire  _GEN19711 = io_x[10] ? _GEN19710 : _GEN7044;
wire  _GEN19712 = io_x[71] ? _GEN19711 : _GEN19697;
wire  _GEN19713 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19714 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN19715 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19716 = io_x[41] ? _GEN6836 : _GEN19715;
wire  _GEN19717 = io_x[14] ? _GEN19716 : _GEN19714;
wire  _GEN19718 = io_x[0] ? _GEN19717 : _GEN19713;
wire  _GEN19719 = io_x[76] ? _GEN19718 : _GEN6834;
wire  _GEN19720 = io_x[42] ? _GEN6874 : _GEN19719;
wire  _GEN19721 = io_x[38] ? _GEN6871 : _GEN19720;
wire  _GEN19722 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN19723 = io_x[76] ? _GEN19722 : _GEN6834;
wire  _GEN19724 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19725 = io_x[41] ? _GEN19724 : _GEN6836;
wire  _GEN19726 = io_x[14] ? _GEN6843 : _GEN19725;
wire  _GEN19727 = io_x[0] ? _GEN6845 : _GEN19726;
wire  _GEN19728 = io_x[76] ? _GEN6834 : _GEN19727;
wire  _GEN19729 = io_x[42] ? _GEN19728 : _GEN19723;
wire  _GEN19730 = io_x[38] ? _GEN6871 : _GEN19729;
wire  _GEN19731 = io_x[10] ? _GEN19730 : _GEN19721;
wire  _GEN19732 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19733 = io_x[38] ? _GEN19732 : _GEN6871;
wire  _GEN19734 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19735 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN19736 = io_x[76] ? _GEN6834 : _GEN19735;
wire  _GEN19737 = io_x[42] ? _GEN19736 : _GEN6874;
wire  _GEN19738 = io_x[38] ? _GEN19737 : _GEN19734;
wire  _GEN19739 = io_x[10] ? _GEN19738 : _GEN19733;
wire  _GEN19740 = io_x[71] ? _GEN19739 : _GEN19731;
wire  _GEN19741 = io_x[70] ? _GEN19740 : _GEN19712;
wire  _GEN19742 = io_x[33] ? _GEN12627 : _GEN19741;
wire  _GEN19743 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN19744 = io_x[38] ? _GEN19743 : _GEN6871;
wire  _GEN19745 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19746 = io_x[38] ? _GEN19745 : _GEN7036;
wire  _GEN19747 = io_x[10] ? _GEN19746 : _GEN19744;
wire  _GEN19748 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN19749 = io_x[38] ? _GEN19748 : _GEN7036;
wire  _GEN19750 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN19751 = io_x[6] ? _GEN19750 : _GEN6850;
wire  _GEN19752 = io_x[41] ? _GEN6836 : _GEN19751;
wire  _GEN19753 = io_x[14] ? _GEN19752 : _GEN6843;
wire  _GEN19754 = io_x[0] ? _GEN19753 : _GEN6845;
wire  _GEN19755 = io_x[76] ? _GEN6834 : _GEN19754;
wire  _GEN19756 = io_x[42] ? _GEN19755 : _GEN6874;
wire  _GEN19757 = io_x[38] ? _GEN19756 : _GEN6871;
wire  _GEN19758 = io_x[10] ? _GEN19757 : _GEN19749;
wire  _GEN19759 = io_x[71] ? _GEN19758 : _GEN19747;
wire  _GEN19760 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19761 = io_x[0] ? _GEN19760 : _GEN6845;
wire  _GEN19762 = io_x[76] ? _GEN6834 : _GEN19761;
wire  _GEN19763 = io_x[42] ? _GEN6874 : _GEN19762;
wire  _GEN19764 = io_x[38] ? _GEN19763 : _GEN6871;
wire  _GEN19765 = io_x[10] ? _GEN19764 : _GEN7044;
wire  _GEN19766 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN19767 = io_x[42] ? _GEN19766 : _GEN6874;
wire  _GEN19768 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN19769 = io_x[6] ? _GEN19768 : _GEN6850;
wire  _GEN19770 = io_x[41] ? _GEN19769 : _GEN6836;
wire  _GEN19771 = io_x[14] ? _GEN19770 : _GEN6843;
wire  _GEN19772 = io_x[0] ? _GEN19771 : _GEN6845;
wire  _GEN19773 = io_x[76] ? _GEN6834 : _GEN19772;
wire  _GEN19774 = io_x[42] ? _GEN6863 : _GEN19773;
wire  _GEN19775 = io_x[38] ? _GEN19774 : _GEN19767;
wire  _GEN19776 = io_x[10] ? _GEN19775 : _GEN7094;
wire  _GEN19777 = io_x[71] ? _GEN19776 : _GEN19765;
wire  _GEN19778 = io_x[70] ? _GEN19777 : _GEN19759;
wire  _GEN19779 = io_x[33] ? _GEN12627 : _GEN19778;
wire  _GEN19780 = io_x[21] ? _GEN19779 : _GEN19742;
wire  _GEN19781 = io_x[18] ? _GEN19780 : _GEN19693;
wire  _GEN19782 = io_x[10] ? _GEN7094 : _GEN7044;
wire  _GEN19783 = io_x[71] ? _GEN19782 : _GEN7203;
wire  _GEN19784 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19785 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19786 = io_x[0] ? _GEN19785 : _GEN19784;
wire  _GEN19787 = io_x[76] ? _GEN19786 : _GEN6834;
wire  _GEN19788 = io_x[42] ? _GEN6874 : _GEN19787;
wire  _GEN19789 = io_x[38] ? _GEN6871 : _GEN19788;
wire  _GEN19790 = io_x[10] ? _GEN7094 : _GEN19789;
wire  _GEN19791 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19792 = io_x[38] ? _GEN19791 : _GEN6871;
wire  _GEN19793 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN19794 = io_x[76] ? _GEN6834 : _GEN19793;
wire  _GEN19795 = io_x[42] ? _GEN19794 : _GEN6863;
wire  _GEN19796 = io_x[38] ? _GEN19795 : _GEN7036;
wire  _GEN19797 = io_x[10] ? _GEN19796 : _GEN19792;
wire  _GEN19798 = io_x[71] ? _GEN19797 : _GEN19790;
wire  _GEN19799 = io_x[70] ? _GEN19798 : _GEN19783;
wire  _GEN19800 = io_x[33] ? _GEN12627 : _GEN19799;
wire  _GEN19801 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19802 = io_x[0] ? _GEN6845 : _GEN19801;
wire  _GEN19803 = io_x[76] ? _GEN19802 : _GEN6834;
wire  _GEN19804 = io_x[42] ? _GEN19803 : _GEN6874;
wire  _GEN19805 = io_x[38] ? _GEN19804 : _GEN7036;
wire  _GEN19806 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19807 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN19808 = io_x[76] ? _GEN19807 : _GEN6833;
wire  _GEN19809 = io_x[42] ? _GEN19808 : _GEN6863;
wire  _GEN19810 = io_x[38] ? _GEN19809 : _GEN19806;
wire  _GEN19811 = io_x[10] ? _GEN19810 : _GEN19805;
wire  _GEN19812 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19813 = io_x[41] ? _GEN19812 : _GEN6836;
wire  _GEN19814 = io_x[14] ? _GEN6843 : _GEN19813;
wire  _GEN19815 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19816 = io_x[0] ? _GEN19815 : _GEN19814;
wire  _GEN19817 = io_x[76] ? _GEN19816 : _GEN6834;
wire  _GEN19818 = io_x[42] ? _GEN19817 : _GEN6874;
wire  _GEN19819 = io_x[38] ? _GEN19818 : _GEN6871;
wire  _GEN19820 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19821 = io_x[0] ? _GEN19820 : _GEN6845;
wire  _GEN19822 = io_x[76] ? _GEN6833 : _GEN19821;
wire  _GEN19823 = io_x[42] ? _GEN6874 : _GEN19822;
wire  _GEN19824 = io_x[38] ? _GEN19823 : _GEN6871;
wire  _GEN19825 = io_x[10] ? _GEN19824 : _GEN19819;
wire  _GEN19826 = io_x[71] ? _GEN19825 : _GEN19811;
wire  _GEN19827 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN19828 = io_x[14] ? _GEN6843 : _GEN19827;
wire  _GEN19829 = io_x[0] ? _GEN6858 : _GEN19828;
wire  _GEN19830 = io_x[76] ? _GEN19829 : _GEN6834;
wire  _GEN19831 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN19832 = io_x[42] ? _GEN19831 : _GEN19830;
wire  _GEN19833 = io_x[38] ? _GEN7036 : _GEN19832;
wire  _GEN19834 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19835 = io_x[0] ? _GEN6845 : _GEN19834;
wire  _GEN19836 = io_x[76] ? _GEN19835 : _GEN6834;
wire  _GEN19837 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN19838 = io_x[42] ? _GEN19837 : _GEN19836;
wire  _GEN19839 = io_x[38] ? _GEN6871 : _GEN19838;
wire  _GEN19840 = io_x[10] ? _GEN19839 : _GEN19833;
wire  _GEN19841 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19842 = io_x[41] ? _GEN6836 : _GEN19841;
wire  _GEN19843 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19844 = io_x[41] ? _GEN6836 : _GEN19843;
wire  _GEN19845 = io_x[14] ? _GEN19844 : _GEN19842;
wire  _GEN19846 = io_x[0] ? _GEN19845 : _GEN6845;
wire  _GEN19847 = io_x[76] ? _GEN19846 : _GEN6833;
wire  _GEN19848 = io_x[42] ? _GEN6874 : _GEN19847;
wire  _GEN19849 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN19850 = io_x[42] ? _GEN19849 : _GEN6874;
wire  _GEN19851 = io_x[38] ? _GEN19850 : _GEN19848;
wire  _GEN19852 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN19853 = io_x[6] ? _GEN19852 : _GEN6850;
wire  _GEN19854 = io_x[41] ? _GEN6836 : _GEN19853;
wire  _GEN19855 = io_x[14] ? _GEN19854 : _GEN6843;
wire  _GEN19856 = io_x[0] ? _GEN6845 : _GEN19855;
wire  _GEN19857 = io_x[76] ? _GEN6834 : _GEN19856;
wire  _GEN19858 = io_x[42] ? _GEN19857 : _GEN6874;
wire  _GEN19859 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19860 = io_x[41] ? _GEN19859 : _GEN6836;
wire  _GEN19861 = io_x[14] ? _GEN6843 : _GEN19860;
wire  _GEN19862 = io_x[0] ? _GEN6845 : _GEN19861;
wire  _GEN19863 = io_x[76] ? _GEN6834 : _GEN19862;
wire  _GEN19864 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN19865 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN19866 = io_x[6] ? _GEN19865 : _GEN6850;
wire  _GEN19867 = io_x[41] ? _GEN6836 : _GEN19866;
wire  _GEN19868 = io_x[14] ? _GEN19867 : _GEN6843;
wire  _GEN19869 = io_x[0] ? _GEN6845 : _GEN19868;
wire  _GEN19870 = io_x[76] ? _GEN19869 : _GEN19864;
wire  _GEN19871 = io_x[42] ? _GEN19870 : _GEN19863;
wire  _GEN19872 = io_x[38] ? _GEN19871 : _GEN19858;
wire  _GEN19873 = io_x[10] ? _GEN19872 : _GEN19851;
wire  _GEN19874 = io_x[71] ? _GEN19873 : _GEN19840;
wire  _GEN19875 = io_x[70] ? _GEN19874 : _GEN19826;
wire  _GEN19876 = io_x[71] ? _GEN7196 : _GEN7203;
wire  _GEN19877 = io_x[70] ? _GEN8474 : _GEN19876;
wire  _GEN19878 = io_x[33] ? _GEN19877 : _GEN19875;
wire  _GEN19879 = io_x[21] ? _GEN19878 : _GEN19800;
wire  _GEN19880 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19881 = io_x[0] ? _GEN6858 : _GEN19880;
wire  _GEN19882 = io_x[76] ? _GEN6834 : _GEN19881;
wire  _GEN19883 = io_x[42] ? _GEN6863 : _GEN19882;
wire  _GEN19884 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN19885 = io_x[6] ? _GEN19884 : _GEN6850;
wire  _GEN19886 = io_x[41] ? _GEN19885 : _GEN6836;
wire  _GEN19887 = io_x[14] ? _GEN19886 : _GEN6843;
wire  _GEN19888 = io_x[0] ? _GEN19887 : _GEN6845;
wire  _GEN19889 = io_x[76] ? _GEN6834 : _GEN19888;
wire  _GEN19890 = io_x[42] ? _GEN6863 : _GEN19889;
wire  _GEN19891 = io_x[38] ? _GEN19890 : _GEN19883;
wire  _GEN19892 = io_x[10] ? _GEN19891 : _GEN7044;
wire  _GEN19893 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN19894 = io_x[10] ? _GEN19893 : _GEN7044;
wire  _GEN19895 = io_x[71] ? _GEN19894 : _GEN19892;
wire  _GEN19896 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN19897 = io_x[38] ? _GEN19896 : _GEN6871;
wire  _GEN19898 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19899 = io_x[0] ? _GEN6845 : _GEN19898;
wire  _GEN19900 = io_x[76] ? _GEN6834 : _GEN19899;
wire  _GEN19901 = io_x[42] ? _GEN19900 : _GEN6874;
wire  _GEN19902 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN19903 = io_x[38] ? _GEN19902 : _GEN19901;
wire  _GEN19904 = io_x[10] ? _GEN19903 : _GEN19897;
wire  _GEN19905 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN19906 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19907 = io_x[0] ? _GEN6845 : _GEN19906;
wire  _GEN19908 = io_x[76] ? _GEN6834 : _GEN19907;
wire  _GEN19909 = io_x[42] ? _GEN19908 : _GEN6874;
wire  _GEN19910 = io_x[38] ? _GEN19909 : _GEN19905;
wire  _GEN19911 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19912 = io_x[0] ? _GEN19911 : _GEN6845;
wire  _GEN19913 = io_x[76] ? _GEN6834 : _GEN19912;
wire  _GEN19914 = io_x[42] ? _GEN19913 : _GEN6863;
wire  _GEN19915 = io_x[38] ? _GEN19914 : _GEN7036;
wire  _GEN19916 = io_x[10] ? _GEN19915 : _GEN19910;
wire  _GEN19917 = io_x[71] ? _GEN19916 : _GEN19904;
wire  _GEN19918 = io_x[70] ? _GEN19917 : _GEN19895;
wire  _GEN19919 = io_x[33] ? _GEN12641 : _GEN19918;
wire  _GEN19920 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN19921 = io_x[76] ? _GEN6834 : _GEN19920;
wire  _GEN19922 = io_x[42] ? _GEN6863 : _GEN19921;
wire  _GEN19923 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19924 = io_x[0] ? _GEN6845 : _GEN19923;
wire  _GEN19925 = io_x[76] ? _GEN19924 : _GEN6834;
wire  _GEN19926 = io_x[42] ? _GEN19925 : _GEN6874;
wire  _GEN19927 = io_x[38] ? _GEN19926 : _GEN19922;
wire  _GEN19928 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN19929 = io_x[6] ? _GEN19928 : _GEN6850;
wire  _GEN19930 = io_x[41] ? _GEN19929 : _GEN6836;
wire  _GEN19931 = io_x[14] ? _GEN19930 : _GEN6843;
wire  _GEN19932 = io_x[0] ? _GEN6858 : _GEN19931;
wire  _GEN19933 = io_x[76] ? _GEN6834 : _GEN19932;
wire  _GEN19934 = io_x[42] ? _GEN6863 : _GEN19933;
wire  _GEN19935 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19936 = io_x[41] ? _GEN19935 : _GEN6836;
wire  _GEN19937 = io_x[14] ? _GEN6856 : _GEN19936;
wire  _GEN19938 = io_x[0] ? _GEN19937 : _GEN6858;
wire  _GEN19939 = io_x[76] ? _GEN6834 : _GEN19938;
wire  _GEN19940 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19941 = io_x[41] ? _GEN6836 : _GEN19940;
wire  _GEN19942 = io_x[14] ? _GEN19941 : _GEN6843;
wire  _GEN19943 = io_x[0] ? _GEN19942 : _GEN6845;
wire  _GEN19944 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN19945 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19946 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19947 = io_x[41] ? _GEN19946 : _GEN19945;
wire  _GEN19948 = io_x[14] ? _GEN19947 : _GEN19944;
wire  _GEN19949 = io_x[0] ? _GEN19948 : _GEN6845;
wire  _GEN19950 = io_x[76] ? _GEN19949 : _GEN19943;
wire  _GEN19951 = io_x[42] ? _GEN19950 : _GEN19939;
wire  _GEN19952 = io_x[38] ? _GEN19951 : _GEN19934;
wire  _GEN19953 = io_x[10] ? _GEN19952 : _GEN19927;
wire  _GEN19954 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN19955 = io_x[0] ? _GEN19954 : _GEN6845;
wire  _GEN19956 = io_x[76] ? _GEN6834 : _GEN19955;
wire  _GEN19957 = io_x[42] ? _GEN6874 : _GEN19956;
wire  _GEN19958 = io_x[38] ? _GEN19957 : _GEN7036;
wire  _GEN19959 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19960 = io_x[41] ? _GEN6836 : _GEN19959;
wire  _GEN19961 = io_x[14] ? _GEN6843 : _GEN19960;
wire  _GEN19962 = io_x[0] ? _GEN19961 : _GEN6845;
wire  _GEN19963 = io_x[76] ? _GEN19962 : _GEN6834;
wire  _GEN19964 = io_x[42] ? _GEN19963 : _GEN6874;
wire  _GEN19965 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19966 = io_x[41] ? _GEN6836 : _GEN19965;
wire  _GEN19967 = io_x[14] ? _GEN19966 : _GEN6843;
wire  _GEN19968 = io_x[0] ? _GEN19967 : _GEN6858;
wire  _GEN19969 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN19970 = io_x[6] ? _GEN19969 : _GEN6840;
wire  _GEN19971 = io_x[41] ? _GEN6836 : _GEN19970;
wire  _GEN19972 = io_x[14] ? _GEN19971 : _GEN6843;
wire  _GEN19973 = io_x[0] ? _GEN19972 : _GEN6858;
wire  _GEN19974 = io_x[76] ? _GEN19973 : _GEN19968;
wire  _GEN19975 = io_x[42] ? _GEN19974 : _GEN6874;
wire  _GEN19976 = io_x[38] ? _GEN19975 : _GEN19964;
wire  _GEN19977 = io_x[10] ? _GEN19976 : _GEN19958;
wire  _GEN19978 = io_x[71] ? _GEN19977 : _GEN19953;
wire  _GEN19979 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN19980 = io_x[0] ? _GEN6845 : _GEN19979;
wire  _GEN19981 = io_x[76] ? _GEN19980 : _GEN6834;
wire  _GEN19982 = io_x[42] ? _GEN19981 : _GEN6874;
wire  _GEN19983 = io_x[38] ? _GEN6871 : _GEN19982;
wire  _GEN19984 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN19985 = io_x[41] ? _GEN19984 : _GEN6836;
wire  _GEN19986 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19987 = io_x[41] ? _GEN19986 : _GEN6836;
wire  _GEN19988 = io_x[14] ? _GEN19987 : _GEN19985;
wire  _GEN19989 = io_x[0] ? _GEN19988 : _GEN6845;
wire  _GEN19990 = io_x[76] ? _GEN6834 : _GEN19989;
wire  _GEN19991 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19992 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN19993 = io_x[41] ? _GEN19992 : _GEN19991;
wire  _GEN19994 = io_x[14] ? _GEN19993 : _GEN6843;
wire  _GEN19995 = io_x[0] ? _GEN6845 : _GEN19994;
wire  _GEN19996 = io_x[76] ? _GEN6834 : _GEN19995;
wire  _GEN19997 = io_x[42] ? _GEN19996 : _GEN19990;
wire  _GEN19998 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN19999 = io_x[6] ? _GEN19998 : _GEN6850;
wire  _GEN20000 = io_x[41] ? _GEN19999 : _GEN6836;
wire  _GEN20001 = io_x[14] ? _GEN20000 : _GEN6843;
wire  _GEN20002 = io_x[0] ? _GEN20001 : _GEN6845;
wire  _GEN20003 = io_x[76] ? _GEN6834 : _GEN20002;
wire  _GEN20004 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN20005 = io_x[41] ? _GEN6836 : _GEN20004;
wire  _GEN20006 = io_x[14] ? _GEN20005 : _GEN6843;
wire  _GEN20007 = io_x[0] ? _GEN20006 : _GEN6858;
wire  _GEN20008 = io_x[76] ? _GEN6834 : _GEN20007;
wire  _GEN20009 = io_x[42] ? _GEN20008 : _GEN20003;
wire  _GEN20010 = io_x[38] ? _GEN20009 : _GEN19997;
wire  _GEN20011 = io_x[10] ? _GEN20010 : _GEN19983;
wire  _GEN20012 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN20013 = io_x[0] ? _GEN20012 : _GEN6845;
wire  _GEN20014 = io_x[76] ? _GEN6833 : _GEN20013;
wire  _GEN20015 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN20016 = io_x[0] ? _GEN6845 : _GEN20015;
wire  _GEN20017 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN20018 = io_x[0] ? _GEN6845 : _GEN20017;
wire  _GEN20019 = io_x[76] ? _GEN20018 : _GEN20016;
wire  _GEN20020 = io_x[42] ? _GEN20019 : _GEN20014;
wire  _GEN20021 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN20022 = io_x[0] ? _GEN6845 : _GEN20021;
wire  _GEN20023 = io_x[76] ? _GEN6834 : _GEN20022;
wire  _GEN20024 = io_x[42] ? _GEN20023 : _GEN6874;
wire  _GEN20025 = io_x[38] ? _GEN20024 : _GEN20020;
wire  _GEN20026 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN20027 = io_x[6] ? _GEN20026 : _GEN6850;
wire  _GEN20028 = io_x[41] ? _GEN20027 : _GEN6836;
wire  _GEN20029 = io_x[14] ? _GEN20028 : _GEN6856;
wire  _GEN20030 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN20031 = io_x[6] ? _GEN20030 : _GEN6840;
wire  _GEN20032 = io_x[41] ? _GEN6836 : _GEN20031;
wire  _GEN20033 = io_x[14] ? _GEN20032 : _GEN6856;
wire  _GEN20034 = io_x[0] ? _GEN20033 : _GEN20029;
wire  _GEN20035 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN20036 = io_x[14] ? _GEN20035 : _GEN6856;
wire  _GEN20037 = io_x[0] ? _GEN20036 : _GEN6845;
wire  _GEN20038 = io_x[76] ? _GEN20037 : _GEN20034;
wire  _GEN20039 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN20040 = io_x[41] ? _GEN6836 : _GEN20039;
wire  _GEN20041 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN20042 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN20043 = io_x[41] ? _GEN20042 : _GEN20041;
wire  _GEN20044 = io_x[14] ? _GEN20043 : _GEN20040;
wire  _GEN20045 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN20046 = io_x[41] ? _GEN6836 : _GEN20045;
wire  _GEN20047 = io_x[14] ? _GEN20046 : _GEN6843;
wire  _GEN20048 = io_x[0] ? _GEN20047 : _GEN20044;
wire  _GEN20049 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN20050 = io_x[6] ? _GEN20049 : _GEN6840;
wire  _GEN20051 = io_x[41] ? _GEN6836 : _GEN20050;
wire  _GEN20052 = io_x[14] ? _GEN20051 : _GEN6856;
wire  _GEN20053 = io_x[0] ? _GEN6845 : _GEN20052;
wire  _GEN20054 = io_x[76] ? _GEN20053 : _GEN20048;
wire  _GEN20055 = io_x[42] ? _GEN20054 : _GEN20038;
wire  _GEN20056 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN20057 = io_x[6] ? _GEN20056 : _GEN6840;
wire  _GEN20058 = io_x[41] ? _GEN20057 : _GEN6836;
wire  _GEN20059 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN20060 = io_x[41] ? _GEN20059 : _GEN6836;
wire  _GEN20061 = io_x[14] ? _GEN20060 : _GEN20058;
wire  _GEN20062 = io_x[0] ? _GEN20061 : _GEN6845;
wire  _GEN20063 = io_x[76] ? _GEN6834 : _GEN20062;
wire  _GEN20064 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN20065 = io_x[41] ? _GEN6836 : _GEN20064;
wire  _GEN20066 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN20067 = io_x[41] ? _GEN6836 : _GEN20066;
wire  _GEN20068 = io_x[14] ? _GEN20067 : _GEN20065;
wire  _GEN20069 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN20070 = io_x[41] ? _GEN6836 : _GEN20069;
wire  _GEN20071 = io_x[14] ? _GEN20070 : _GEN6843;
wire  _GEN20072 = io_x[0] ? _GEN20071 : _GEN20068;
wire  _GEN20073 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN20074 = io_x[14] ? _GEN20073 : _GEN6856;
wire  _GEN20075 = io_x[0] ? _GEN20074 : _GEN6845;
wire  _GEN20076 = io_x[76] ? _GEN20075 : _GEN20072;
wire  _GEN20077 = io_x[42] ? _GEN20076 : _GEN20063;
wire  _GEN20078 = io_x[38] ? _GEN20077 : _GEN20055;
wire  _GEN20079 = io_x[10] ? _GEN20078 : _GEN20025;
wire  _GEN20080 = io_x[71] ? _GEN20079 : _GEN20011;
wire  _GEN20081 = io_x[70] ? _GEN20080 : _GEN19978;
wire  _GEN20082 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN20083 = io_x[41] ? _GEN20082 : _GEN6836;
wire  _GEN20084 = io_x[14] ? _GEN6843 : _GEN20083;
wire  _GEN20085 = io_x[0] ? _GEN20084 : _GEN6845;
wire  _GEN20086 = io_x[76] ? _GEN6834 : _GEN20085;
wire  _GEN20087 = io_x[42] ? _GEN6863 : _GEN20086;
wire  _GEN20088 = io_x[38] ? _GEN20087 : _GEN7036;
wire  _GEN20089 = io_x[10] ? _GEN20088 : _GEN7044;
wire  _GEN20090 = io_x[71] ? _GEN7196 : _GEN20089;
wire  _GEN20091 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN20092 = io_x[10] ? _GEN20091 : _GEN7044;
wire  _GEN20093 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN20094 = io_x[0] ? _GEN20093 : _GEN6845;
wire  _GEN20095 = io_x[76] ? _GEN6834 : _GEN20094;
wire  _GEN20096 = io_x[42] ? _GEN20095 : _GEN6874;
wire  _GEN20097 = io_x[38] ? _GEN20096 : _GEN7036;
wire  _GEN20098 = io_x[10] ? _GEN20097 : _GEN7044;
wire  _GEN20099 = io_x[71] ? _GEN20098 : _GEN20092;
wire  _GEN20100 = io_x[70] ? _GEN20099 : _GEN20090;
wire  _GEN20101 = io_x[33] ? _GEN20100 : _GEN20081;
wire  _GEN20102 = io_x[21] ? _GEN20101 : _GEN19919;
wire  _GEN20103 = io_x[18] ? _GEN20102 : _GEN19879;
wire  _GEN20104 = io_x[20] ? _GEN20103 : _GEN19781;
wire  _GEN20105 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN20106 = io_x[0] ? _GEN20105 : _GEN6845;
wire  _GEN20107 = io_x[76] ? _GEN6834 : _GEN20106;
wire  _GEN20108 = io_x[42] ? _GEN6874 : _GEN20107;
wire  _GEN20109 = io_x[38] ? _GEN20108 : _GEN7036;
wire  _GEN20110 = io_x[10] ? _GEN20109 : _GEN7094;
wire  _GEN20111 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN20112 = io_x[10] ? _GEN7044 : _GEN20111;
wire  _GEN20113 = io_x[71] ? _GEN20112 : _GEN20110;
wire  _GEN20114 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN20115 = io_x[42] ? _GEN6874 : _GEN20114;
wire  _GEN20116 = io_x[38] ? _GEN20115 : _GEN6871;
wire  _GEN20117 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN20118 = io_x[41] ? _GEN6924 : _GEN20117;
wire  _GEN20119 = io_x[14] ? _GEN20118 : _GEN6843;
wire  _GEN20120 = io_x[0] ? _GEN6845 : _GEN20119;
wire  _GEN20121 = io_x[76] ? _GEN20120 : _GEN6834;
wire  _GEN20122 = io_x[42] ? _GEN6874 : _GEN20121;
wire  _GEN20123 = io_x[38] ? _GEN20122 : _GEN6871;
wire  _GEN20124 = io_x[10] ? _GEN20123 : _GEN20116;
wire  _GEN20125 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN20126 = io_x[10] ? _GEN7044 : _GEN20125;
wire  _GEN20127 = io_x[71] ? _GEN20126 : _GEN20124;
wire  _GEN20128 = io_x[70] ? _GEN20127 : _GEN20113;
wire  _GEN20129 = io_x[33] ? _GEN12641 : _GEN20128;
wire  _GEN20130 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN20131 = io_x[38] ? _GEN20130 : _GEN6871;
wire  _GEN20132 = io_x[10] ? _GEN7044 : _GEN20131;
wire  _GEN20133 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN20134 = io_x[42] ? _GEN20133 : _GEN6874;
wire  _GEN20135 = io_x[38] ? _GEN20134 : _GEN6871;
wire  _GEN20136 = io_x[10] ? _GEN20135 : _GEN7094;
wire  _GEN20137 = io_x[71] ? _GEN20136 : _GEN20132;
wire  _GEN20138 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN20139 = io_x[41] ? _GEN20138 : _GEN6836;
wire  _GEN20140 = io_x[14] ? _GEN20139 : _GEN6843;
wire  _GEN20141 = io_x[0] ? _GEN20140 : _GEN6845;
wire  _GEN20142 = io_x[76] ? _GEN20141 : _GEN6834;
wire  _GEN20143 = io_x[42] ? _GEN20142 : _GEN6863;
wire  _GEN20144 = io_x[38] ? _GEN20143 : _GEN6871;
wire  _GEN20145 = io_x[10] ? _GEN20144 : _GEN7094;
wire  _GEN20146 = io_x[71] ? _GEN20145 : _GEN7203;
wire  _GEN20147 = io_x[70] ? _GEN20146 : _GEN20137;
wire  _GEN20148 = io_x[33] ? _GEN12641 : _GEN20147;
wire  _GEN20149 = io_x[21] ? _GEN20148 : _GEN20129;
wire  _GEN20150 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN20151 = io_x[42] ? _GEN20150 : _GEN6863;
wire  _GEN20152 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN20153 = io_x[76] ? _GEN6834 : _GEN20152;
wire  _GEN20154 = io_x[42] ? _GEN6874 : _GEN20153;
wire  _GEN20155 = io_x[38] ? _GEN20154 : _GEN20151;
wire  _GEN20156 = io_x[10] ? _GEN20155 : _GEN7044;
wire  _GEN20157 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN20158 = io_x[38] ? _GEN20157 : _GEN6871;
wire  _GEN20159 = io_x[10] ? _GEN20158 : _GEN7094;
wire  _GEN20160 = io_x[71] ? _GEN20159 : _GEN20156;
wire  _GEN20161 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN20162 = io_x[38] ? _GEN7036 : _GEN20161;
wire  _GEN20163 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN20164 = io_x[0] ? _GEN20163 : _GEN6845;
wire  _GEN20165 = io_x[76] ? _GEN6834 : _GEN20164;
wire  _GEN20166 = io_x[42] ? _GEN6874 : _GEN20165;
wire  _GEN20167 = io_x[38] ? _GEN7036 : _GEN20166;
wire  _GEN20168 = io_x[10] ? _GEN20167 : _GEN20162;
wire  _GEN20169 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN20170 = io_x[10] ? _GEN20169 : _GEN7044;
wire  _GEN20171 = io_x[71] ? _GEN20170 : _GEN20168;
wire  _GEN20172 = io_x[70] ? _GEN20171 : _GEN20160;
wire  _GEN20173 = io_x[33] ? _GEN12641 : _GEN20172;
wire  _GEN20174 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN20175 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN20176 = io_x[41] ? _GEN6836 : _GEN20175;
wire  _GEN20177 = io_x[14] ? _GEN20176 : _GEN6843;
wire  _GEN20178 = io_x[0] ? _GEN20177 : _GEN6845;
wire  _GEN20179 = io_x[76] ? _GEN6834 : _GEN20178;
wire  _GEN20180 = io_x[42] ? _GEN6874 : _GEN20179;
wire  _GEN20181 = io_x[38] ? _GEN6871 : _GEN20180;
wire  _GEN20182 = io_x[10] ? _GEN20181 : _GEN20174;
wire  _GEN20183 = io_x[71] ? _GEN20182 : _GEN7196;
wire  _GEN20184 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN20185 = io_x[14] ? _GEN20184 : _GEN6843;
wire  _GEN20186 = io_x[0] ? _GEN20185 : _GEN6845;
wire  _GEN20187 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN20188 = io_x[0] ? _GEN6845 : _GEN20187;
wire  _GEN20189 = io_x[76] ? _GEN20188 : _GEN20186;
wire  _GEN20190 = io_x[42] ? _GEN6874 : _GEN20189;
wire  _GEN20191 = io_x[38] ? _GEN6871 : _GEN20190;
wire  _GEN20192 = io_x[10] ? _GEN20191 : _GEN7094;
wire  _GEN20193 = io_x[2] ? _GEN6837 : _GEN6838;
wire  _GEN20194 = io_x[6] ? _GEN20193 : _GEN6850;
wire  _GEN20195 = io_x[41] ? _GEN6836 : _GEN20194;
wire  _GEN20196 = io_x[14] ? _GEN20195 : _GEN6843;
wire  _GEN20197 = io_x[0] ? _GEN20196 : _GEN6845;
wire  _GEN20198 = io_x[76] ? _GEN20197 : _GEN6834;
wire  _GEN20199 = io_x[42] ? _GEN6874 : _GEN20198;
wire  _GEN20200 = io_x[38] ? _GEN20199 : _GEN7036;
wire  _GEN20201 = io_x[10] ? _GEN20200 : _GEN7044;
wire  _GEN20202 = io_x[71] ? _GEN20201 : _GEN20192;
wire  _GEN20203 = io_x[70] ? _GEN20202 : _GEN20183;
wire  _GEN20204 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN20205 = io_x[41] ? _GEN6836 : _GEN20204;
wire  _GEN20206 = io_x[14] ? _GEN20205 : _GEN6843;
wire  _GEN20207 = io_x[0] ? _GEN20206 : _GEN6845;
wire  _GEN20208 = io_x[76] ? _GEN6834 : _GEN20207;
wire  _GEN20209 = io_x[42] ? _GEN6874 : _GEN20208;
wire  _GEN20210 = io_x[38] ? _GEN6871 : _GEN20209;
wire  _GEN20211 = io_x[10] ? _GEN20210 : _GEN7044;
wire  _GEN20212 = io_x[71] ? _GEN20211 : _GEN7196;
wire  _GEN20213 = io_x[70] ? _GEN8474 : _GEN20212;
wire  _GEN20214 = io_x[33] ? _GEN20213 : _GEN20203;
wire  _GEN20215 = io_x[21] ? _GEN20214 : _GEN20173;
wire  _GEN20216 = io_x[18] ? _GEN20215 : _GEN20149;
wire  _GEN20217 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN20218 = io_x[38] ? _GEN6871 : _GEN7036;
wire  _GEN20219 = io_x[10] ? _GEN20218 : _GEN20217;
wire  _GEN20220 = io_x[2] ? _GEN6838 : _GEN6837;
wire  _GEN20221 = io_x[6] ? _GEN20220 : _GEN6850;
wire  _GEN20222 = io_x[41] ? _GEN6836 : _GEN20221;
wire  _GEN20223 = io_x[14] ? _GEN20222 : _GEN6843;
wire  _GEN20224 = io_x[0] ? _GEN6845 : _GEN20223;
wire  _GEN20225 = io_x[76] ? _GEN6834 : _GEN20224;
wire  _GEN20226 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN20227 = io_x[42] ? _GEN20226 : _GEN20225;
wire  _GEN20228 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN20229 = io_x[42] ? _GEN6863 : _GEN20228;
wire  _GEN20230 = io_x[38] ? _GEN20229 : _GEN20227;
wire  _GEN20231 = io_x[10] ? _GEN20230 : _GEN7094;
wire  _GEN20232 = io_x[71] ? _GEN20231 : _GEN20219;
wire  _GEN20233 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN20234 = io_x[0] ? _GEN6845 : _GEN6858;
wire  _GEN20235 = io_x[76] ? _GEN20234 : _GEN6833;
wire  _GEN20236 = io_x[42] ? _GEN20235 : _GEN20233;
wire  _GEN20237 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN20238 = io_x[38] ? _GEN20237 : _GEN20236;
wire  _GEN20239 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN20240 = io_x[10] ? _GEN20239 : _GEN20238;
wire  _GEN20241 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN20242 = io_x[14] ? _GEN6843 : _GEN20241;
wire  _GEN20243 = io_x[0] ? _GEN6845 : _GEN20242;
wire  _GEN20244 = io_x[76] ? _GEN6834 : _GEN20243;
wire  _GEN20245 = io_x[42] ? _GEN6874 : _GEN20244;
wire  _GEN20246 = io_x[38] ? _GEN20245 : _GEN7036;
wire  _GEN20247 = io_x[42] ? _GEN6874 : _GEN6863;
wire  _GEN20248 = io_x[38] ? _GEN6871 : _GEN20247;
wire  _GEN20249 = io_x[10] ? _GEN20248 : _GEN20246;
wire  _GEN20250 = io_x[71] ? _GEN20249 : _GEN20240;
wire  _GEN20251 = io_x[70] ? _GEN20250 : _GEN20232;
wire  _GEN20252 = io_x[33] ? _GEN12641 : _GEN20251;
wire  _GEN20253 = io_x[21] ? _GEN20252 : _GEN12643;
wire  _GEN20254 = io_x[38] ? _GEN7036 : _GEN6871;
wire  _GEN20255 = io_x[10] ? _GEN7044 : _GEN20254;
wire  _GEN20256 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN20257 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN20258 = io_x[0] ? _GEN20257 : _GEN20256;
wire  _GEN20259 = io_x[76] ? _GEN6833 : _GEN20258;
wire  _GEN20260 = io_x[42] ? _GEN6874 : _GEN20259;
wire  _GEN20261 = io_x[41] ? _GEN6836 : _GEN6924;
wire  _GEN20262 = io_x[14] ? _GEN20261 : _GEN6856;
wire  _GEN20263 = io_x[0] ? _GEN20262 : _GEN6858;
wire  _GEN20264 = io_x[76] ? _GEN20263 : _GEN6833;
wire  _GEN20265 = io_x[42] ? _GEN20264 : _GEN6874;
wire  _GEN20266 = io_x[38] ? _GEN20265 : _GEN20260;
wire  _GEN20267 = io_x[10] ? _GEN20266 : _GEN7094;
wire  _GEN20268 = io_x[71] ? _GEN20267 : _GEN20255;
wire  _GEN20269 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN20270 = io_x[0] ? _GEN20269 : _GEN6845;
wire  _GEN20271 = io_x[76] ? _GEN20270 : _GEN6834;
wire  _GEN20272 = io_x[42] ? _GEN20271 : _GEN6863;
wire  _GEN20273 = io_x[38] ? _GEN7036 : _GEN20272;
wire  _GEN20274 = io_x[10] ? _GEN20273 : _GEN7094;
wire  _GEN20275 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN20276 = io_x[0] ? _GEN20275 : _GEN6845;
wire  _GEN20277 = io_x[76] ? _GEN6834 : _GEN20276;
wire  _GEN20278 = io_x[42] ? _GEN6874 : _GEN20277;
wire  _GEN20279 = io_x[38] ? _GEN6871 : _GEN20278;
wire  _GEN20280 = io_x[10] ? _GEN20279 : _GEN7044;
wire  _GEN20281 = io_x[71] ? _GEN20280 : _GEN20274;
wire  _GEN20282 = io_x[70] ? _GEN20281 : _GEN20268;
wire  _GEN20283 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN20284 = io_x[0] ? _GEN20283 : _GEN6845;
wire  _GEN20285 = io_x[76] ? _GEN6834 : _GEN20284;
wire  _GEN20286 = io_x[42] ? _GEN6874 : _GEN20285;
wire  _GEN20287 = io_x[38] ? _GEN6871 : _GEN20286;
wire  _GEN20288 = io_x[10] ? _GEN20287 : _GEN7044;
wire  _GEN20289 = io_x[71] ? _GEN20288 : _GEN7196;
wire  _GEN20290 = io_x[70] ? _GEN7020 : _GEN20289;
wire  _GEN20291 = io_x[33] ? _GEN20290 : _GEN20282;
wire  _GEN20292 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN20293 = io_x[0] ? _GEN6845 : _GEN20292;
wire  _GEN20294 = io_x[76] ? _GEN6834 : _GEN20293;
wire  _GEN20295 = io_x[42] ? _GEN6874 : _GEN20294;
wire  _GEN20296 = io_x[38] ? _GEN20295 : _GEN6871;
wire  _GEN20297 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN20298 = io_x[14] ? _GEN20297 : _GEN6843;
wire  _GEN20299 = io_x[0] ? _GEN6845 : _GEN20298;
wire  _GEN20300 = io_x[76] ? _GEN6834 : _GEN20299;
wire  _GEN20301 = io_x[42] ? _GEN20300 : _GEN6874;
wire  _GEN20302 = io_x[38] ? _GEN6871 : _GEN20301;
wire  _GEN20303 = io_x[10] ? _GEN20302 : _GEN20296;
wire  _GEN20304 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN20305 = io_x[42] ? _GEN6874 : _GEN20304;
wire  _GEN20306 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN20307 = io_x[0] ? _GEN6858 : _GEN20306;
wire  _GEN20308 = io_x[76] ? _GEN6834 : _GEN20307;
wire  _GEN20309 = io_x[42] ? _GEN6874 : _GEN20308;
wire  _GEN20310 = io_x[38] ? _GEN20309 : _GEN20305;
wire  _GEN20311 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN20312 = io_x[41] ? _GEN6836 : _GEN20311;
wire  _GEN20313 = io_x[14] ? _GEN20312 : _GEN6843;
wire  _GEN20314 = io_x[0] ? _GEN20313 : _GEN6858;
wire  _GEN20315 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN20316 = io_x[41] ? _GEN6836 : _GEN20315;
wire  _GEN20317 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN20318 = io_x[41] ? _GEN6836 : _GEN20317;
wire  _GEN20319 = io_x[14] ? _GEN20318 : _GEN20316;
wire  _GEN20320 = io_x[0] ? _GEN20319 : _GEN6845;
wire  _GEN20321 = io_x[76] ? _GEN20320 : _GEN20314;
wire  _GEN20322 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN20323 = io_x[76] ? _GEN6833 : _GEN20322;
wire  _GEN20324 = io_x[42] ? _GEN20323 : _GEN20321;
wire  _GEN20325 = io_x[76] ? _GEN6833 : _GEN6834;
wire  _GEN20326 = io_x[42] ? _GEN6874 : _GEN20325;
wire  _GEN20327 = io_x[38] ? _GEN20326 : _GEN20324;
wire  _GEN20328 = io_x[10] ? _GEN20327 : _GEN20310;
wire  _GEN20329 = io_x[71] ? _GEN20328 : _GEN20303;
wire  _GEN20330 = io_x[14] ? _GEN6843 : _GEN6856;
wire  _GEN20331 = io_x[0] ? _GEN6845 : _GEN20330;
wire  _GEN20332 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN20333 = io_x[0] ? _GEN6845 : _GEN20332;
wire  _GEN20334 = io_x[76] ? _GEN20333 : _GEN20331;
wire  _GEN20335 = io_x[42] ? _GEN6863 : _GEN20334;
wire  _GEN20336 = io_x[42] ? _GEN6863 : _GEN6874;
wire  _GEN20337 = io_x[38] ? _GEN20336 : _GEN20335;
wire  _GEN20338 = io_x[0] ? _GEN6858 : _GEN6845;
wire  _GEN20339 = io_x[6] ? _GEN6840 : _GEN6850;
wire  _GEN20340 = io_x[41] ? _GEN6836 : _GEN20339;
wire  _GEN20341 = io_x[6] ? _GEN6850 : _GEN6840;
wire  _GEN20342 = io_x[41] ? _GEN6836 : _GEN20341;
wire  _GEN20343 = io_x[14] ? _GEN20342 : _GEN20340;
wire  _GEN20344 = io_x[0] ? _GEN20343 : _GEN6845;
wire  _GEN20345 = io_x[76] ? _GEN20344 : _GEN20338;
wire  _GEN20346 = io_x[41] ? _GEN6924 : _GEN6836;
wire  _GEN20347 = io_x[14] ? _GEN20346 : _GEN6843;
wire  _GEN20348 = io_x[0] ? _GEN20347 : _GEN6845;
wire  _GEN20349 = io_x[76] ? _GEN20348 : _GEN6834;
wire  _GEN20350 = io_x[42] ? _GEN20349 : _GEN20345;
wire  _GEN20351 = io_x[38] ? _GEN7036 : _GEN20350;
wire  _GEN20352 = io_x[10] ? _GEN20351 : _GEN20337;
wire  _GEN20353 = io_x[76] ? _GEN6834 : _GEN6833;
wire  _GEN20354 = io_x[42] ? _GEN20353 : _GEN6874;
wire  _GEN20355 = io_x[38] ? _GEN20354 : _GEN6871;
wire  _GEN20356 = io_x[14] ? _GEN6856 : _GEN6843;
wire  _GEN20357 = io_x[0] ? _GEN6845 : _GEN20356;
wire  _GEN20358 = io_x[76] ? _GEN6834 : _GEN20357;
wire  _GEN20359 = io_x[42] ? _GEN6863 : _GEN20358;
wire  _GEN20360 = io_x[38] ? _GEN20359 : _GEN7036;
wire  _GEN20361 = io_x[10] ? _GEN20360 : _GEN20355;
wire  _GEN20362 = io_x[71] ? _GEN20361 : _GEN20352;
wire  _GEN20363 = io_x[70] ? _GEN20362 : _GEN20329;
wire  _GEN20364 = io_x[10] ? _GEN7044 : _GEN7094;
wire  _GEN20365 = io_x[71] ? _GEN20364 : _GEN7196;
wire  _GEN20366 = io_x[71] ? _GEN7196 : _GEN7203;
wire  _GEN20367 = io_x[70] ? _GEN20366 : _GEN20365;
wire  _GEN20368 = io_x[33] ? _GEN20367 : _GEN20363;
wire  _GEN20369 = io_x[21] ? _GEN20368 : _GEN20291;
wire  _GEN20370 = io_x[18] ? _GEN20369 : _GEN20253;
wire  _GEN20371 = io_x[20] ? _GEN20370 : _GEN20216;
wire  _GEN20372 = io_x[45] ? _GEN20371 : _GEN20104;
wire  _GEN20373 = io_x[28] ? _GEN20372 : _GEN19569;
wire  _GEN20374 = io_x[79] ? _GEN20373 : _GEN18836;
wire  _GEN20375 = io_x[48] ? _GEN20374 : _GEN18749;
wire  _GEN20376 = io_x[47] ? _GEN20375 : _GEN14309;
assign io_y[8] = _GEN20376;
wire  _GEN20377 = 1'b0;
wire  _GEN20378 = 1'b1;
wire  _GEN20379 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20380 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20381 = io_x[5] ? _GEN20380 : _GEN20379;
wire  _GEN20382 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20383 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20384 = io_x[5] ? _GEN20383 : _GEN20382;
wire  _GEN20385 = io_x[1] ? _GEN20384 : _GEN20381;
wire  _GEN20386 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20387 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20388 = io_x[5] ? _GEN20387 : _GEN20386;
wire  _GEN20389 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20390 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20391 = io_x[5] ? _GEN20390 : _GEN20389;
wire  _GEN20392 = io_x[1] ? _GEN20391 : _GEN20388;
wire  _GEN20393 = io_x[9] ? _GEN20392 : _GEN20385;
wire  _GEN20394 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20395 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20396 = io_x[5] ? _GEN20395 : _GEN20394;
wire  _GEN20397 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20398 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20399 = io_x[5] ? _GEN20398 : _GEN20397;
wire  _GEN20400 = io_x[1] ? _GEN20399 : _GEN20396;
wire  _GEN20401 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20402 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20403 = io_x[5] ? _GEN20402 : _GEN20401;
wire  _GEN20404 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20405 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20406 = io_x[5] ? _GEN20405 : _GEN20404;
wire  _GEN20407 = io_x[1] ? _GEN20406 : _GEN20403;
wire  _GEN20408 = io_x[9] ? _GEN20407 : _GEN20400;
wire  _GEN20409 = io_x[13] ? _GEN20408 : _GEN20393;
wire  _GEN20410 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20411 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20412 = io_x[5] ? _GEN20411 : _GEN20410;
wire  _GEN20413 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20414 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20415 = io_x[5] ? _GEN20414 : _GEN20413;
wire  _GEN20416 = io_x[1] ? _GEN20415 : _GEN20412;
wire  _GEN20417 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20418 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20419 = io_x[5] ? _GEN20418 : _GEN20417;
wire  _GEN20420 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20421 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20422 = io_x[5] ? _GEN20421 : _GEN20420;
wire  _GEN20423 = io_x[1] ? _GEN20422 : _GEN20419;
wire  _GEN20424 = io_x[9] ? _GEN20423 : _GEN20416;
wire  _GEN20425 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20426 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20427 = io_x[5] ? _GEN20426 : _GEN20425;
wire  _GEN20428 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20429 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20430 = io_x[5] ? _GEN20429 : _GEN20428;
wire  _GEN20431 = io_x[1] ? _GEN20430 : _GEN20427;
wire  _GEN20432 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20433 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20434 = io_x[5] ? _GEN20433 : _GEN20432;
wire  _GEN20435 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20436 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20437 = io_x[5] ? _GEN20436 : _GEN20435;
wire  _GEN20438 = io_x[1] ? _GEN20437 : _GEN20434;
wire  _GEN20439 = io_x[9] ? _GEN20438 : _GEN20431;
wire  _GEN20440 = io_x[13] ? _GEN20439 : _GEN20424;
wire  _GEN20441 = io_x[44] ? _GEN20440 : _GEN20409;
wire  _GEN20442 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20443 = 1'b1;
wire  _GEN20444 = io_x[5] ? _GEN20443 : _GEN20442;
wire  _GEN20445 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20446 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20447 = io_x[5] ? _GEN20446 : _GEN20445;
wire  _GEN20448 = io_x[1] ? _GEN20447 : _GEN20444;
wire  _GEN20449 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20450 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20451 = io_x[5] ? _GEN20450 : _GEN20449;
wire  _GEN20452 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20453 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20454 = io_x[5] ? _GEN20453 : _GEN20452;
wire  _GEN20455 = io_x[1] ? _GEN20454 : _GEN20451;
wire  _GEN20456 = io_x[9] ? _GEN20455 : _GEN20448;
wire  _GEN20457 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20458 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20459 = io_x[5] ? _GEN20458 : _GEN20457;
wire  _GEN20460 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20461 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20462 = io_x[5] ? _GEN20461 : _GEN20460;
wire  _GEN20463 = io_x[1] ? _GEN20462 : _GEN20459;
wire  _GEN20464 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20465 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20466 = io_x[5] ? _GEN20465 : _GEN20464;
wire  _GEN20467 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20468 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20469 = io_x[5] ? _GEN20468 : _GEN20467;
wire  _GEN20470 = io_x[1] ? _GEN20469 : _GEN20466;
wire  _GEN20471 = io_x[9] ? _GEN20470 : _GEN20463;
wire  _GEN20472 = io_x[13] ? _GEN20471 : _GEN20456;
wire  _GEN20473 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20474 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20475 = io_x[5] ? _GEN20474 : _GEN20473;
wire  _GEN20476 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20477 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20478 = io_x[5] ? _GEN20477 : _GEN20476;
wire  _GEN20479 = io_x[1] ? _GEN20478 : _GEN20475;
wire  _GEN20480 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20481 = 1'b0;
wire  _GEN20482 = io_x[5] ? _GEN20481 : _GEN20480;
wire  _GEN20483 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20484 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20485 = io_x[5] ? _GEN20484 : _GEN20483;
wire  _GEN20486 = io_x[1] ? _GEN20485 : _GEN20482;
wire  _GEN20487 = io_x[9] ? _GEN20486 : _GEN20479;
wire  _GEN20488 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20489 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20490 = io_x[5] ? _GEN20489 : _GEN20488;
wire  _GEN20491 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20492 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20493 = io_x[5] ? _GEN20492 : _GEN20491;
wire  _GEN20494 = io_x[1] ? _GEN20493 : _GEN20490;
wire  _GEN20495 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20496 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20497 = io_x[5] ? _GEN20496 : _GEN20495;
wire  _GEN20498 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20499 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20500 = io_x[5] ? _GEN20499 : _GEN20498;
wire  _GEN20501 = io_x[1] ? _GEN20500 : _GEN20497;
wire  _GEN20502 = io_x[9] ? _GEN20501 : _GEN20494;
wire  _GEN20503 = io_x[13] ? _GEN20502 : _GEN20487;
wire  _GEN20504 = io_x[44] ? _GEN20503 : _GEN20472;
wire  _GEN20505 = io_x[37] ? _GEN20504 : _GEN20441;
wire  _GEN20506 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20507 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20508 = io_x[5] ? _GEN20507 : _GEN20506;
wire  _GEN20509 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20510 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20511 = io_x[5] ? _GEN20510 : _GEN20509;
wire  _GEN20512 = io_x[1] ? _GEN20511 : _GEN20508;
wire  _GEN20513 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20514 = io_x[5] ? _GEN20513 : _GEN20443;
wire  _GEN20515 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20516 = io_x[5] ? _GEN20515 : _GEN20481;
wire  _GEN20517 = io_x[1] ? _GEN20516 : _GEN20514;
wire  _GEN20518 = io_x[9] ? _GEN20517 : _GEN20512;
wire  _GEN20519 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20520 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20521 = io_x[5] ? _GEN20520 : _GEN20519;
wire  _GEN20522 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20523 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20524 = io_x[5] ? _GEN20523 : _GEN20522;
wire  _GEN20525 = io_x[1] ? _GEN20524 : _GEN20521;
wire  _GEN20526 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20527 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20528 = io_x[5] ? _GEN20527 : _GEN20526;
wire  _GEN20529 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20530 = io_x[5] ? _GEN20481 : _GEN20529;
wire  _GEN20531 = io_x[1] ? _GEN20530 : _GEN20528;
wire  _GEN20532 = io_x[9] ? _GEN20531 : _GEN20525;
wire  _GEN20533 = io_x[13] ? _GEN20532 : _GEN20518;
wire  _GEN20534 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20535 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20536 = io_x[5] ? _GEN20535 : _GEN20534;
wire  _GEN20537 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20538 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20539 = io_x[5] ? _GEN20538 : _GEN20537;
wire  _GEN20540 = io_x[1] ? _GEN20539 : _GEN20536;
wire  _GEN20541 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20542 = io_x[5] ? _GEN20481 : _GEN20541;
wire  _GEN20543 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20544 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20545 = io_x[5] ? _GEN20544 : _GEN20543;
wire  _GEN20546 = io_x[1] ? _GEN20545 : _GEN20542;
wire  _GEN20547 = io_x[9] ? _GEN20546 : _GEN20540;
wire  _GEN20548 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20549 = io_x[5] ? _GEN20481 : _GEN20548;
wire  _GEN20550 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20551 = io_x[5] ? _GEN20443 : _GEN20550;
wire  _GEN20552 = io_x[1] ? _GEN20551 : _GEN20549;
wire  _GEN20553 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20554 = io_x[5] ? _GEN20443 : _GEN20553;
wire  _GEN20555 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20556 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20557 = io_x[5] ? _GEN20556 : _GEN20555;
wire  _GEN20558 = io_x[1] ? _GEN20557 : _GEN20554;
wire  _GEN20559 = io_x[9] ? _GEN20558 : _GEN20552;
wire  _GEN20560 = io_x[13] ? _GEN20559 : _GEN20547;
wire  _GEN20561 = io_x[44] ? _GEN20560 : _GEN20533;
wire  _GEN20562 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20563 = io_x[5] ? _GEN20443 : _GEN20562;
wire  _GEN20564 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20565 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20566 = io_x[5] ? _GEN20565 : _GEN20564;
wire  _GEN20567 = io_x[1] ? _GEN20566 : _GEN20563;
wire  _GEN20568 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20569 = io_x[5] ? _GEN20568 : _GEN20443;
wire  _GEN20570 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20571 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20572 = io_x[5] ? _GEN20571 : _GEN20570;
wire  _GEN20573 = io_x[1] ? _GEN20572 : _GEN20569;
wire  _GEN20574 = io_x[9] ? _GEN20573 : _GEN20567;
wire  _GEN20575 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20576 = io_x[5] ? _GEN20481 : _GEN20575;
wire  _GEN20577 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20578 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20579 = io_x[5] ? _GEN20578 : _GEN20577;
wire  _GEN20580 = io_x[1] ? _GEN20579 : _GEN20576;
wire  _GEN20581 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20582 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20583 = io_x[5] ? _GEN20582 : _GEN20581;
wire  _GEN20584 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20585 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20586 = io_x[5] ? _GEN20585 : _GEN20584;
wire  _GEN20587 = io_x[1] ? _GEN20586 : _GEN20583;
wire  _GEN20588 = io_x[9] ? _GEN20587 : _GEN20580;
wire  _GEN20589 = io_x[13] ? _GEN20588 : _GEN20574;
wire  _GEN20590 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20591 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20592 = io_x[5] ? _GEN20591 : _GEN20590;
wire  _GEN20593 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20594 = io_x[5] ? _GEN20593 : _GEN20443;
wire  _GEN20595 = io_x[1] ? _GEN20594 : _GEN20592;
wire  _GEN20596 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20597 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20598 = io_x[5] ? _GEN20597 : _GEN20596;
wire  _GEN20599 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20600 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20601 = io_x[5] ? _GEN20600 : _GEN20599;
wire  _GEN20602 = io_x[1] ? _GEN20601 : _GEN20598;
wire  _GEN20603 = io_x[9] ? _GEN20602 : _GEN20595;
wire  _GEN20604 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20605 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20606 = io_x[5] ? _GEN20605 : _GEN20604;
wire  _GEN20607 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20608 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20609 = io_x[5] ? _GEN20608 : _GEN20607;
wire  _GEN20610 = io_x[1] ? _GEN20609 : _GEN20606;
wire  _GEN20611 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20612 = io_x[5] ? _GEN20611 : _GEN20481;
wire  _GEN20613 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20614 = io_x[5] ? _GEN20613 : _GEN20443;
wire  _GEN20615 = io_x[1] ? _GEN20614 : _GEN20612;
wire  _GEN20616 = io_x[9] ? _GEN20615 : _GEN20610;
wire  _GEN20617 = io_x[13] ? _GEN20616 : _GEN20603;
wire  _GEN20618 = io_x[44] ? _GEN20617 : _GEN20589;
wire  _GEN20619 = io_x[37] ? _GEN20618 : _GEN20561;
wire  _GEN20620 = io_x[38] ? _GEN20619 : _GEN20505;
wire  _GEN20621 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20622 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20623 = io_x[5] ? _GEN20622 : _GEN20621;
wire  _GEN20624 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20625 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20626 = io_x[5] ? _GEN20625 : _GEN20624;
wire  _GEN20627 = io_x[1] ? _GEN20626 : _GEN20623;
wire  _GEN20628 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20629 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20630 = io_x[5] ? _GEN20629 : _GEN20628;
wire  _GEN20631 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20632 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20633 = io_x[5] ? _GEN20632 : _GEN20631;
wire  _GEN20634 = io_x[1] ? _GEN20633 : _GEN20630;
wire  _GEN20635 = io_x[9] ? _GEN20634 : _GEN20627;
wire  _GEN20636 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20637 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20638 = io_x[5] ? _GEN20637 : _GEN20636;
wire  _GEN20639 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20640 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20641 = io_x[5] ? _GEN20640 : _GEN20639;
wire  _GEN20642 = io_x[1] ? _GEN20641 : _GEN20638;
wire  _GEN20643 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20644 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20645 = io_x[5] ? _GEN20644 : _GEN20643;
wire  _GEN20646 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20647 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20648 = io_x[5] ? _GEN20647 : _GEN20646;
wire  _GEN20649 = io_x[1] ? _GEN20648 : _GEN20645;
wire  _GEN20650 = io_x[9] ? _GEN20649 : _GEN20642;
wire  _GEN20651 = io_x[13] ? _GEN20650 : _GEN20635;
wire  _GEN20652 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20653 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20654 = io_x[5] ? _GEN20653 : _GEN20652;
wire  _GEN20655 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20656 = io_x[5] ? _GEN20655 : _GEN20443;
wire  _GEN20657 = io_x[1] ? _GEN20656 : _GEN20654;
wire  _GEN20658 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20659 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20660 = io_x[5] ? _GEN20659 : _GEN20658;
wire  _GEN20661 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20662 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20663 = io_x[5] ? _GEN20662 : _GEN20661;
wire  _GEN20664 = io_x[1] ? _GEN20663 : _GEN20660;
wire  _GEN20665 = io_x[9] ? _GEN20664 : _GEN20657;
wire  _GEN20666 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20667 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20668 = io_x[5] ? _GEN20667 : _GEN20666;
wire  _GEN20669 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20670 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20671 = io_x[5] ? _GEN20670 : _GEN20669;
wire  _GEN20672 = io_x[1] ? _GEN20671 : _GEN20668;
wire  _GEN20673 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20674 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20675 = io_x[5] ? _GEN20674 : _GEN20673;
wire  _GEN20676 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20677 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20678 = io_x[5] ? _GEN20677 : _GEN20676;
wire  _GEN20679 = io_x[1] ? _GEN20678 : _GEN20675;
wire  _GEN20680 = io_x[9] ? _GEN20679 : _GEN20672;
wire  _GEN20681 = io_x[13] ? _GEN20680 : _GEN20665;
wire  _GEN20682 = io_x[44] ? _GEN20681 : _GEN20651;
wire  _GEN20683 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20684 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20685 = io_x[5] ? _GEN20684 : _GEN20683;
wire  _GEN20686 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20687 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20688 = io_x[5] ? _GEN20687 : _GEN20686;
wire  _GEN20689 = io_x[1] ? _GEN20688 : _GEN20685;
wire  _GEN20690 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20691 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20692 = io_x[5] ? _GEN20691 : _GEN20690;
wire  _GEN20693 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20694 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20695 = io_x[5] ? _GEN20694 : _GEN20693;
wire  _GEN20696 = io_x[1] ? _GEN20695 : _GEN20692;
wire  _GEN20697 = io_x[9] ? _GEN20696 : _GEN20689;
wire  _GEN20698 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20699 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20700 = io_x[5] ? _GEN20699 : _GEN20698;
wire  _GEN20701 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20702 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20703 = io_x[5] ? _GEN20702 : _GEN20701;
wire  _GEN20704 = io_x[1] ? _GEN20703 : _GEN20700;
wire  _GEN20705 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20706 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20707 = io_x[5] ? _GEN20706 : _GEN20705;
wire  _GEN20708 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20709 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20710 = io_x[5] ? _GEN20709 : _GEN20708;
wire  _GEN20711 = io_x[1] ? _GEN20710 : _GEN20707;
wire  _GEN20712 = io_x[9] ? _GEN20711 : _GEN20704;
wire  _GEN20713 = io_x[13] ? _GEN20712 : _GEN20697;
wire  _GEN20714 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20715 = io_x[5] ? _GEN20443 : _GEN20714;
wire  _GEN20716 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20717 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20718 = io_x[5] ? _GEN20717 : _GEN20716;
wire  _GEN20719 = io_x[1] ? _GEN20718 : _GEN20715;
wire  _GEN20720 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20721 = io_x[5] ? _GEN20720 : _GEN20443;
wire  _GEN20722 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20723 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20724 = io_x[5] ? _GEN20723 : _GEN20722;
wire  _GEN20725 = io_x[1] ? _GEN20724 : _GEN20721;
wire  _GEN20726 = io_x[9] ? _GEN20725 : _GEN20719;
wire  _GEN20727 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20728 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20729 = io_x[5] ? _GEN20728 : _GEN20727;
wire  _GEN20730 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20731 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20732 = io_x[5] ? _GEN20731 : _GEN20730;
wire  _GEN20733 = io_x[1] ? _GEN20732 : _GEN20729;
wire  _GEN20734 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20735 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20736 = io_x[5] ? _GEN20735 : _GEN20734;
wire  _GEN20737 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20738 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20739 = io_x[5] ? _GEN20738 : _GEN20737;
wire  _GEN20740 = io_x[1] ? _GEN20739 : _GEN20736;
wire  _GEN20741 = io_x[9] ? _GEN20740 : _GEN20733;
wire  _GEN20742 = io_x[13] ? _GEN20741 : _GEN20726;
wire  _GEN20743 = io_x[44] ? _GEN20742 : _GEN20713;
wire  _GEN20744 = io_x[37] ? _GEN20743 : _GEN20682;
wire  _GEN20745 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20746 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20747 = io_x[5] ? _GEN20746 : _GEN20745;
wire  _GEN20748 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20749 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20750 = io_x[5] ? _GEN20749 : _GEN20748;
wire  _GEN20751 = io_x[1] ? _GEN20750 : _GEN20747;
wire  _GEN20752 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20753 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20754 = io_x[5] ? _GEN20753 : _GEN20752;
wire  _GEN20755 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20756 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20757 = io_x[5] ? _GEN20756 : _GEN20755;
wire  _GEN20758 = io_x[1] ? _GEN20757 : _GEN20754;
wire  _GEN20759 = io_x[9] ? _GEN20758 : _GEN20751;
wire  _GEN20760 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20761 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20762 = io_x[5] ? _GEN20761 : _GEN20760;
wire  _GEN20763 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20764 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20765 = io_x[5] ? _GEN20764 : _GEN20763;
wire  _GEN20766 = io_x[1] ? _GEN20765 : _GEN20762;
wire  _GEN20767 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20768 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20769 = io_x[5] ? _GEN20768 : _GEN20767;
wire  _GEN20770 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20771 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20772 = io_x[5] ? _GEN20771 : _GEN20770;
wire  _GEN20773 = io_x[1] ? _GEN20772 : _GEN20769;
wire  _GEN20774 = io_x[9] ? _GEN20773 : _GEN20766;
wire  _GEN20775 = io_x[13] ? _GEN20774 : _GEN20759;
wire  _GEN20776 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20777 = io_x[5] ? _GEN20443 : _GEN20776;
wire  _GEN20778 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20779 = io_x[5] ? _GEN20778 : _GEN20443;
wire  _GEN20780 = io_x[1] ? _GEN20779 : _GEN20777;
wire  _GEN20781 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20782 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20783 = io_x[5] ? _GEN20782 : _GEN20781;
wire  _GEN20784 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20785 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20786 = io_x[5] ? _GEN20785 : _GEN20784;
wire  _GEN20787 = io_x[1] ? _GEN20786 : _GEN20783;
wire  _GEN20788 = io_x[9] ? _GEN20787 : _GEN20780;
wire  _GEN20789 = io_x[5] ? _GEN20481 : _GEN20443;
wire  _GEN20790 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20791 = io_x[5] ? _GEN20790 : _GEN20481;
wire  _GEN20792 = io_x[1] ? _GEN20791 : _GEN20789;
wire  _GEN20793 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20794 = io_x[5] ? _GEN20793 : _GEN20481;
wire  _GEN20795 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20796 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20797 = io_x[5] ? _GEN20796 : _GEN20795;
wire  _GEN20798 = io_x[1] ? _GEN20797 : _GEN20794;
wire  _GEN20799 = io_x[9] ? _GEN20798 : _GEN20792;
wire  _GEN20800 = io_x[13] ? _GEN20799 : _GEN20788;
wire  _GEN20801 = io_x[44] ? _GEN20800 : _GEN20775;
wire  _GEN20802 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20803 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20804 = io_x[5] ? _GEN20803 : _GEN20802;
wire  _GEN20805 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20806 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20807 = io_x[5] ? _GEN20806 : _GEN20805;
wire  _GEN20808 = io_x[1] ? _GEN20807 : _GEN20804;
wire  _GEN20809 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20810 = io_x[5] ? _GEN20481 : _GEN20809;
wire  _GEN20811 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20812 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20813 = io_x[5] ? _GEN20812 : _GEN20811;
wire  _GEN20814 = io_x[1] ? _GEN20813 : _GEN20810;
wire  _GEN20815 = io_x[9] ? _GEN20814 : _GEN20808;
wire  _GEN20816 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20817 = io_x[5] ? _GEN20816 : _GEN20443;
wire  _GEN20818 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20819 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20820 = io_x[5] ? _GEN20819 : _GEN20818;
wire  _GEN20821 = io_x[1] ? _GEN20820 : _GEN20817;
wire  _GEN20822 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20823 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20824 = io_x[5] ? _GEN20823 : _GEN20822;
wire  _GEN20825 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20826 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20827 = io_x[5] ? _GEN20826 : _GEN20825;
wire  _GEN20828 = io_x[1] ? _GEN20827 : _GEN20824;
wire  _GEN20829 = io_x[9] ? _GEN20828 : _GEN20821;
wire  _GEN20830 = io_x[13] ? _GEN20829 : _GEN20815;
wire  _GEN20831 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20832 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20833 = io_x[5] ? _GEN20832 : _GEN20831;
wire  _GEN20834 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20835 = io_x[5] ? _GEN20834 : _GEN20443;
wire  _GEN20836 = io_x[1] ? _GEN20835 : _GEN20833;
wire  _GEN20837 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20838 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20839 = io_x[5] ? _GEN20838 : _GEN20837;
wire  _GEN20840 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20841 = io_x[5] ? _GEN20840 : _GEN20481;
wire  _GEN20842 = io_x[1] ? _GEN20841 : _GEN20839;
wire  _GEN20843 = io_x[9] ? _GEN20842 : _GEN20836;
wire  _GEN20844 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20845 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20846 = io_x[5] ? _GEN20845 : _GEN20844;
wire  _GEN20847 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20848 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20849 = io_x[5] ? _GEN20848 : _GEN20847;
wire  _GEN20850 = io_x[1] ? _GEN20849 : _GEN20846;
wire  _GEN20851 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20852 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20853 = io_x[5] ? _GEN20852 : _GEN20851;
wire  _GEN20854 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20855 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20856 = io_x[5] ? _GEN20855 : _GEN20854;
wire  _GEN20857 = io_x[1] ? _GEN20856 : _GEN20853;
wire  _GEN20858 = io_x[9] ? _GEN20857 : _GEN20850;
wire  _GEN20859 = io_x[13] ? _GEN20858 : _GEN20843;
wire  _GEN20860 = io_x[44] ? _GEN20859 : _GEN20830;
wire  _GEN20861 = io_x[37] ? _GEN20860 : _GEN20801;
wire  _GEN20862 = io_x[38] ? _GEN20861 : _GEN20744;
wire  _GEN20863 = io_x[24] ? _GEN20862 : _GEN20620;
wire  _GEN20864 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20865 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20866 = io_x[5] ? _GEN20865 : _GEN20864;
wire  _GEN20867 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20868 = io_x[5] ? _GEN20443 : _GEN20867;
wire  _GEN20869 = io_x[1] ? _GEN20868 : _GEN20866;
wire  _GEN20870 = io_x[5] ? _GEN20443 : _GEN20481;
wire  _GEN20871 = io_x[5] ? _GEN20481 : _GEN20443;
wire  _GEN20872 = io_x[1] ? _GEN20871 : _GEN20870;
wire  _GEN20873 = io_x[9] ? _GEN20872 : _GEN20869;
wire  _GEN20874 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20875 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20876 = io_x[5] ? _GEN20875 : _GEN20874;
wire  _GEN20877 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20878 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20879 = io_x[5] ? _GEN20878 : _GEN20877;
wire  _GEN20880 = io_x[1] ? _GEN20879 : _GEN20876;
wire  _GEN20881 = io_x[5] ? _GEN20481 : _GEN20443;
wire  _GEN20882 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20883 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20884 = io_x[5] ? _GEN20883 : _GEN20882;
wire  _GEN20885 = io_x[1] ? _GEN20884 : _GEN20881;
wire  _GEN20886 = io_x[9] ? _GEN20885 : _GEN20880;
wire  _GEN20887 = io_x[13] ? _GEN20886 : _GEN20873;
wire  _GEN20888 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20889 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20890 = io_x[5] ? _GEN20889 : _GEN20888;
wire  _GEN20891 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20892 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20893 = io_x[5] ? _GEN20892 : _GEN20891;
wire  _GEN20894 = io_x[1] ? _GEN20893 : _GEN20890;
wire  _GEN20895 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20896 = io_x[5] ? _GEN20895 : _GEN20481;
wire  _GEN20897 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20898 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20899 = io_x[5] ? _GEN20898 : _GEN20897;
wire  _GEN20900 = io_x[1] ? _GEN20899 : _GEN20896;
wire  _GEN20901 = io_x[9] ? _GEN20900 : _GEN20894;
wire  _GEN20902 = io_x[5] ? _GEN20443 : _GEN20481;
wire  _GEN20903 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20904 = io_x[5] ? _GEN20481 : _GEN20903;
wire  _GEN20905 = io_x[1] ? _GEN20904 : _GEN20902;
wire  _GEN20906 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20907 = io_x[5] ? _GEN20906 : _GEN20443;
wire  _GEN20908 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20909 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20910 = io_x[5] ? _GEN20909 : _GEN20908;
wire  _GEN20911 = io_x[1] ? _GEN20910 : _GEN20907;
wire  _GEN20912 = io_x[9] ? _GEN20911 : _GEN20905;
wire  _GEN20913 = io_x[13] ? _GEN20912 : _GEN20901;
wire  _GEN20914 = io_x[44] ? _GEN20913 : _GEN20887;
wire  _GEN20915 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20916 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20917 = io_x[5] ? _GEN20916 : _GEN20915;
wire  _GEN20918 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20919 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20920 = io_x[5] ? _GEN20919 : _GEN20918;
wire  _GEN20921 = io_x[1] ? _GEN20920 : _GEN20917;
wire  _GEN20922 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20923 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20924 = io_x[5] ? _GEN20923 : _GEN20922;
wire  _GEN20925 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20926 = io_x[5] ? _GEN20481 : _GEN20925;
wire  _GEN20927 = io_x[1] ? _GEN20926 : _GEN20924;
wire  _GEN20928 = io_x[9] ? _GEN20927 : _GEN20921;
wire  _GEN20929 = io_x[5] ? _GEN20443 : _GEN20481;
wire  _GEN20930 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20931 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20932 = io_x[5] ? _GEN20931 : _GEN20930;
wire  _GEN20933 = io_x[1] ? _GEN20932 : _GEN20929;
wire  _GEN20934 = io_x[5] ? _GEN20481 : _GEN20443;
wire  _GEN20935 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20936 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20937 = io_x[5] ? _GEN20936 : _GEN20935;
wire  _GEN20938 = io_x[1] ? _GEN20937 : _GEN20934;
wire  _GEN20939 = io_x[9] ? _GEN20938 : _GEN20933;
wire  _GEN20940 = io_x[13] ? _GEN20939 : _GEN20928;
wire  _GEN20941 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20942 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20943 = io_x[5] ? _GEN20942 : _GEN20941;
wire  _GEN20944 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20945 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20946 = io_x[5] ? _GEN20945 : _GEN20944;
wire  _GEN20947 = io_x[1] ? _GEN20946 : _GEN20943;
wire  _GEN20948 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20949 = io_x[5] ? _GEN20948 : _GEN20481;
wire  _GEN20950 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20951 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20952 = io_x[5] ? _GEN20951 : _GEN20950;
wire  _GEN20953 = io_x[1] ? _GEN20952 : _GEN20949;
wire  _GEN20954 = io_x[9] ? _GEN20953 : _GEN20947;
wire  _GEN20955 = io_x[5] ? _GEN20443 : _GEN20481;
wire  _GEN20956 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20957 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20958 = io_x[5] ? _GEN20957 : _GEN20956;
wire  _GEN20959 = io_x[1] ? _GEN20958 : _GEN20955;
wire  _GEN20960 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20961 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20962 = io_x[5] ? _GEN20961 : _GEN20960;
wire  _GEN20963 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20964 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20965 = io_x[5] ? _GEN20964 : _GEN20963;
wire  _GEN20966 = io_x[1] ? _GEN20965 : _GEN20962;
wire  _GEN20967 = io_x[9] ? _GEN20966 : _GEN20959;
wire  _GEN20968 = io_x[13] ? _GEN20967 : _GEN20954;
wire  _GEN20969 = io_x[44] ? _GEN20968 : _GEN20940;
wire  _GEN20970 = io_x[37] ? _GEN20969 : _GEN20914;
wire  _GEN20971 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20972 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20973 = io_x[5] ? _GEN20972 : _GEN20971;
wire  _GEN20974 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20975 = io_x[5] ? _GEN20443 : _GEN20974;
wire  _GEN20976 = io_x[1] ? _GEN20975 : _GEN20973;
wire  _GEN20977 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20978 = io_x[5] ? _GEN20443 : _GEN20977;
wire  _GEN20979 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20980 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20981 = io_x[5] ? _GEN20980 : _GEN20979;
wire  _GEN20982 = io_x[1] ? _GEN20981 : _GEN20978;
wire  _GEN20983 = io_x[9] ? _GEN20982 : _GEN20976;
wire  _GEN20984 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20985 = io_x[5] ? _GEN20443 : _GEN20984;
wire  _GEN20986 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20987 = io_x[5] ? _GEN20481 : _GEN20986;
wire  _GEN20988 = io_x[1] ? _GEN20987 : _GEN20985;
wire  _GEN20989 = io_x[5] ? _GEN20481 : _GEN20443;
wire  _GEN20990 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20991 = io_x[5] ? _GEN20990 : _GEN20481;
wire  _GEN20992 = io_x[1] ? _GEN20991 : _GEN20989;
wire  _GEN20993 = io_x[9] ? _GEN20992 : _GEN20988;
wire  _GEN20994 = io_x[13] ? _GEN20993 : _GEN20983;
wire  _GEN20995 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN20996 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20997 = io_x[5] ? _GEN20996 : _GEN20995;
wire  _GEN20998 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN20999 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21000 = io_x[5] ? _GEN20999 : _GEN20998;
wire  _GEN21001 = io_x[1] ? _GEN21000 : _GEN20997;
wire  _GEN21002 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21003 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21004 = io_x[5] ? _GEN21003 : _GEN21002;
wire  _GEN21005 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21006 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21007 = io_x[5] ? _GEN21006 : _GEN21005;
wire  _GEN21008 = io_x[1] ? _GEN21007 : _GEN21004;
wire  _GEN21009 = io_x[9] ? _GEN21008 : _GEN21001;
wire  _GEN21010 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21011 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21012 = io_x[5] ? _GEN21011 : _GEN21010;
wire  _GEN21013 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21014 = io_x[5] ? _GEN20481 : _GEN21013;
wire  _GEN21015 = io_x[1] ? _GEN21014 : _GEN21012;
wire  _GEN21016 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21017 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21018 = io_x[5] ? _GEN21017 : _GEN21016;
wire  _GEN21019 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21020 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21021 = io_x[5] ? _GEN21020 : _GEN21019;
wire  _GEN21022 = io_x[1] ? _GEN21021 : _GEN21018;
wire  _GEN21023 = io_x[9] ? _GEN21022 : _GEN21015;
wire  _GEN21024 = io_x[13] ? _GEN21023 : _GEN21009;
wire  _GEN21025 = io_x[44] ? _GEN21024 : _GEN20994;
wire  _GEN21026 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21027 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21028 = io_x[5] ? _GEN21027 : _GEN21026;
wire  _GEN21029 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21030 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21031 = io_x[5] ? _GEN21030 : _GEN21029;
wire  _GEN21032 = io_x[1] ? _GEN21031 : _GEN21028;
wire  _GEN21033 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21034 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21035 = io_x[5] ? _GEN21034 : _GEN21033;
wire  _GEN21036 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21037 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21038 = io_x[5] ? _GEN21037 : _GEN21036;
wire  _GEN21039 = io_x[1] ? _GEN21038 : _GEN21035;
wire  _GEN21040 = io_x[9] ? _GEN21039 : _GEN21032;
wire  _GEN21041 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21042 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21043 = io_x[5] ? _GEN21042 : _GEN21041;
wire  _GEN21044 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21045 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21046 = io_x[5] ? _GEN21045 : _GEN21044;
wire  _GEN21047 = io_x[1] ? _GEN21046 : _GEN21043;
wire  _GEN21048 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21049 = io_x[5] ? _GEN21048 : _GEN20443;
wire  _GEN21050 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21051 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21052 = io_x[5] ? _GEN21051 : _GEN21050;
wire  _GEN21053 = io_x[1] ? _GEN21052 : _GEN21049;
wire  _GEN21054 = io_x[9] ? _GEN21053 : _GEN21047;
wire  _GEN21055 = io_x[13] ? _GEN21054 : _GEN21040;
wire  _GEN21056 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21057 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21058 = io_x[5] ? _GEN21057 : _GEN21056;
wire  _GEN21059 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21060 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21061 = io_x[5] ? _GEN21060 : _GEN21059;
wire  _GEN21062 = io_x[1] ? _GEN21061 : _GEN21058;
wire  _GEN21063 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21064 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21065 = io_x[5] ? _GEN21064 : _GEN21063;
wire  _GEN21066 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21067 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21068 = io_x[5] ? _GEN21067 : _GEN21066;
wire  _GEN21069 = io_x[1] ? _GEN21068 : _GEN21065;
wire  _GEN21070 = io_x[9] ? _GEN21069 : _GEN21062;
wire  _GEN21071 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21072 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21073 = io_x[5] ? _GEN21072 : _GEN21071;
wire  _GEN21074 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21075 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21076 = io_x[5] ? _GEN21075 : _GEN21074;
wire  _GEN21077 = io_x[1] ? _GEN21076 : _GEN21073;
wire  _GEN21078 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21079 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21080 = io_x[5] ? _GEN21079 : _GEN21078;
wire  _GEN21081 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21082 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21083 = io_x[5] ? _GEN21082 : _GEN21081;
wire  _GEN21084 = io_x[1] ? _GEN21083 : _GEN21080;
wire  _GEN21085 = io_x[9] ? _GEN21084 : _GEN21077;
wire  _GEN21086 = io_x[13] ? _GEN21085 : _GEN21070;
wire  _GEN21087 = io_x[44] ? _GEN21086 : _GEN21055;
wire  _GEN21088 = io_x[37] ? _GEN21087 : _GEN21025;
wire  _GEN21089 = io_x[38] ? _GEN21088 : _GEN20970;
wire  _GEN21090 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21091 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21092 = io_x[5] ? _GEN21091 : _GEN21090;
wire  _GEN21093 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21094 = io_x[5] ? _GEN21093 : _GEN20481;
wire  _GEN21095 = io_x[1] ? _GEN21094 : _GEN21092;
wire  _GEN21096 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21097 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21098 = io_x[5] ? _GEN21097 : _GEN21096;
wire  _GEN21099 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21100 = io_x[5] ? _GEN20481 : _GEN21099;
wire  _GEN21101 = io_x[1] ? _GEN21100 : _GEN21098;
wire  _GEN21102 = io_x[9] ? _GEN21101 : _GEN21095;
wire  _GEN21103 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21104 = io_x[5] ? _GEN20443 : _GEN21103;
wire  _GEN21105 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21106 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21107 = io_x[5] ? _GEN21106 : _GEN21105;
wire  _GEN21108 = io_x[1] ? _GEN21107 : _GEN21104;
wire  _GEN21109 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21110 = io_x[5] ? _GEN21109 : _GEN20443;
wire  _GEN21111 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21112 = io_x[5] ? _GEN21111 : _GEN20481;
wire  _GEN21113 = io_x[1] ? _GEN21112 : _GEN21110;
wire  _GEN21114 = io_x[9] ? _GEN21113 : _GEN21108;
wire  _GEN21115 = io_x[13] ? _GEN21114 : _GEN21102;
wire  _GEN21116 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21117 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21118 = io_x[5] ? _GEN21117 : _GEN21116;
wire  _GEN21119 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21120 = io_x[5] ? _GEN21119 : _GEN20443;
wire  _GEN21121 = io_x[1] ? _GEN21120 : _GEN21118;
wire  _GEN21122 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21123 = io_x[5] ? _GEN21122 : _GEN20481;
wire  _GEN21124 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21125 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21126 = io_x[5] ? _GEN21125 : _GEN21124;
wire  _GEN21127 = io_x[1] ? _GEN21126 : _GEN21123;
wire  _GEN21128 = io_x[9] ? _GEN21127 : _GEN21121;
wire  _GEN21129 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21130 = io_x[5] ? _GEN21129 : _GEN20481;
wire  _GEN21131 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21132 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21133 = io_x[5] ? _GEN21132 : _GEN21131;
wire  _GEN21134 = io_x[1] ? _GEN21133 : _GEN21130;
wire  _GEN21135 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21136 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21137 = io_x[5] ? _GEN21136 : _GEN21135;
wire  _GEN21138 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21139 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21140 = io_x[5] ? _GEN21139 : _GEN21138;
wire  _GEN21141 = io_x[1] ? _GEN21140 : _GEN21137;
wire  _GEN21142 = io_x[9] ? _GEN21141 : _GEN21134;
wire  _GEN21143 = io_x[13] ? _GEN21142 : _GEN21128;
wire  _GEN21144 = io_x[44] ? _GEN21143 : _GEN21115;
wire  _GEN21145 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21146 = io_x[5] ? _GEN20481 : _GEN21145;
wire  _GEN21147 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21148 = io_x[5] ? _GEN21147 : _GEN20481;
wire  _GEN21149 = io_x[1] ? _GEN21148 : _GEN21146;
wire  _GEN21150 = io_x[5] ? _GEN20443 : _GEN20481;
wire  _GEN21151 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21152 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21153 = io_x[5] ? _GEN21152 : _GEN21151;
wire  _GEN21154 = io_x[1] ? _GEN21153 : _GEN21150;
wire  _GEN21155 = io_x[9] ? _GEN21154 : _GEN21149;
wire  _GEN21156 = io_x[5] ? _GEN20443 : _GEN20481;
wire  _GEN21157 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21158 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21159 = io_x[5] ? _GEN21158 : _GEN21157;
wire  _GEN21160 = io_x[1] ? _GEN21159 : _GEN21156;
wire  _GEN21161 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21162 = io_x[5] ? _GEN21161 : _GEN20443;
wire  _GEN21163 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21164 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21165 = io_x[5] ? _GEN21164 : _GEN21163;
wire  _GEN21166 = io_x[1] ? _GEN21165 : _GEN21162;
wire  _GEN21167 = io_x[9] ? _GEN21166 : _GEN21160;
wire  _GEN21168 = io_x[13] ? _GEN21167 : _GEN21155;
wire  _GEN21169 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21170 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21171 = io_x[5] ? _GEN21170 : _GEN21169;
wire  _GEN21172 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21173 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21174 = io_x[5] ? _GEN21173 : _GEN21172;
wire  _GEN21175 = io_x[1] ? _GEN21174 : _GEN21171;
wire  _GEN21176 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21177 = io_x[5] ? _GEN21176 : _GEN20481;
wire  _GEN21178 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21179 = io_x[5] ? _GEN21178 : _GEN20481;
wire  _GEN21180 = io_x[1] ? _GEN21179 : _GEN21177;
wire  _GEN21181 = io_x[9] ? _GEN21180 : _GEN21175;
wire  _GEN21182 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21183 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21184 = io_x[5] ? _GEN21183 : _GEN21182;
wire  _GEN21185 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21186 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21187 = io_x[5] ? _GEN21186 : _GEN21185;
wire  _GEN21188 = io_x[1] ? _GEN21187 : _GEN21184;
wire  _GEN21189 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21190 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21191 = io_x[5] ? _GEN21190 : _GEN21189;
wire  _GEN21192 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21193 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21194 = io_x[5] ? _GEN21193 : _GEN21192;
wire  _GEN21195 = io_x[1] ? _GEN21194 : _GEN21191;
wire  _GEN21196 = io_x[9] ? _GEN21195 : _GEN21188;
wire  _GEN21197 = io_x[13] ? _GEN21196 : _GEN21181;
wire  _GEN21198 = io_x[44] ? _GEN21197 : _GEN21168;
wire  _GEN21199 = io_x[37] ? _GEN21198 : _GEN21144;
wire  _GEN21200 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21201 = io_x[5] ? _GEN20481 : _GEN21200;
wire  _GEN21202 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21203 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21204 = io_x[5] ? _GEN21203 : _GEN21202;
wire  _GEN21205 = io_x[1] ? _GEN21204 : _GEN21201;
wire  _GEN21206 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21207 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21208 = io_x[5] ? _GEN21207 : _GEN21206;
wire  _GEN21209 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21210 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21211 = io_x[5] ? _GEN21210 : _GEN21209;
wire  _GEN21212 = io_x[1] ? _GEN21211 : _GEN21208;
wire  _GEN21213 = io_x[9] ? _GEN21212 : _GEN21205;
wire  _GEN21214 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21215 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21216 = io_x[5] ? _GEN21215 : _GEN21214;
wire  _GEN21217 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21218 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21219 = io_x[5] ? _GEN21218 : _GEN21217;
wire  _GEN21220 = io_x[1] ? _GEN21219 : _GEN21216;
wire  _GEN21221 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21222 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21223 = io_x[5] ? _GEN21222 : _GEN21221;
wire  _GEN21224 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21225 = io_x[5] ? _GEN21224 : _GEN20481;
wire  _GEN21226 = io_x[1] ? _GEN21225 : _GEN21223;
wire  _GEN21227 = io_x[9] ? _GEN21226 : _GEN21220;
wire  _GEN21228 = io_x[13] ? _GEN21227 : _GEN21213;
wire  _GEN21229 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21230 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21231 = io_x[5] ? _GEN21230 : _GEN21229;
wire  _GEN21232 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21233 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21234 = io_x[5] ? _GEN21233 : _GEN21232;
wire  _GEN21235 = io_x[1] ? _GEN21234 : _GEN21231;
wire  _GEN21236 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21237 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21238 = io_x[5] ? _GEN21237 : _GEN21236;
wire  _GEN21239 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21240 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21241 = io_x[5] ? _GEN21240 : _GEN21239;
wire  _GEN21242 = io_x[1] ? _GEN21241 : _GEN21238;
wire  _GEN21243 = io_x[9] ? _GEN21242 : _GEN21235;
wire  _GEN21244 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21245 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21246 = io_x[5] ? _GEN21245 : _GEN21244;
wire  _GEN21247 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21248 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21249 = io_x[5] ? _GEN21248 : _GEN21247;
wire  _GEN21250 = io_x[1] ? _GEN21249 : _GEN21246;
wire  _GEN21251 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21252 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21253 = io_x[5] ? _GEN21252 : _GEN21251;
wire  _GEN21254 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21255 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21256 = io_x[5] ? _GEN21255 : _GEN21254;
wire  _GEN21257 = io_x[1] ? _GEN21256 : _GEN21253;
wire  _GEN21258 = io_x[9] ? _GEN21257 : _GEN21250;
wire  _GEN21259 = io_x[13] ? _GEN21258 : _GEN21243;
wire  _GEN21260 = io_x[44] ? _GEN21259 : _GEN21228;
wire  _GEN21261 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21262 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21263 = io_x[5] ? _GEN21262 : _GEN21261;
wire  _GEN21264 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21265 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21266 = io_x[5] ? _GEN21265 : _GEN21264;
wire  _GEN21267 = io_x[1] ? _GEN21266 : _GEN21263;
wire  _GEN21268 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21269 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21270 = io_x[5] ? _GEN21269 : _GEN21268;
wire  _GEN21271 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21272 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21273 = io_x[5] ? _GEN21272 : _GEN21271;
wire  _GEN21274 = io_x[1] ? _GEN21273 : _GEN21270;
wire  _GEN21275 = io_x[9] ? _GEN21274 : _GEN21267;
wire  _GEN21276 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21277 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21278 = io_x[5] ? _GEN21277 : _GEN21276;
wire  _GEN21279 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21280 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21281 = io_x[5] ? _GEN21280 : _GEN21279;
wire  _GEN21282 = io_x[1] ? _GEN21281 : _GEN21278;
wire  _GEN21283 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21284 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21285 = io_x[5] ? _GEN21284 : _GEN21283;
wire  _GEN21286 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21287 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21288 = io_x[5] ? _GEN21287 : _GEN21286;
wire  _GEN21289 = io_x[1] ? _GEN21288 : _GEN21285;
wire  _GEN21290 = io_x[9] ? _GEN21289 : _GEN21282;
wire  _GEN21291 = io_x[13] ? _GEN21290 : _GEN21275;
wire  _GEN21292 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21293 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21294 = io_x[5] ? _GEN21293 : _GEN21292;
wire  _GEN21295 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21296 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21297 = io_x[5] ? _GEN21296 : _GEN21295;
wire  _GEN21298 = io_x[1] ? _GEN21297 : _GEN21294;
wire  _GEN21299 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21300 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21301 = io_x[5] ? _GEN21300 : _GEN21299;
wire  _GEN21302 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21303 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21304 = io_x[5] ? _GEN21303 : _GEN21302;
wire  _GEN21305 = io_x[1] ? _GEN21304 : _GEN21301;
wire  _GEN21306 = io_x[9] ? _GEN21305 : _GEN21298;
wire  _GEN21307 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21308 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21309 = io_x[5] ? _GEN21308 : _GEN21307;
wire  _GEN21310 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21311 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21312 = io_x[5] ? _GEN21311 : _GEN21310;
wire  _GEN21313 = io_x[1] ? _GEN21312 : _GEN21309;
wire  _GEN21314 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21315 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21316 = io_x[5] ? _GEN21315 : _GEN21314;
wire  _GEN21317 = io_x[43] ? _GEN20377 : _GEN20378;
wire  _GEN21318 = io_x[43] ? _GEN20378 : _GEN20377;
wire  _GEN21319 = io_x[5] ? _GEN21318 : _GEN21317;
wire  _GEN21320 = io_x[1] ? _GEN21319 : _GEN21316;
wire  _GEN21321 = io_x[9] ? _GEN21320 : _GEN21313;
wire  _GEN21322 = io_x[13] ? _GEN21321 : _GEN21306;
wire  _GEN21323 = io_x[44] ? _GEN21322 : _GEN21291;
wire  _GEN21324 = io_x[37] ? _GEN21323 : _GEN21260;
wire  _GEN21325 = io_x[38] ? _GEN21324 : _GEN21199;
wire  _GEN21326 = io_x[24] ? _GEN21325 : _GEN21089;
wire  _GEN21327 = io_x[75] ? _GEN21326 : _GEN20863;
assign io_y[7] = _GEN21327;
wire  _GEN21328 = 1'b0;
wire  _GEN21329 = 1'b1;
wire  _GEN21330 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21331 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21332 = io_x[8] ? _GEN21331 : _GEN21330;
wire  _GEN21333 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21334 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21335 = io_x[8] ? _GEN21334 : _GEN21333;
wire  _GEN21336 = io_x[12] ? _GEN21335 : _GEN21332;
wire  _GEN21337 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21338 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21339 = io_x[8] ? _GEN21338 : _GEN21337;
wire  _GEN21340 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21341 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21342 = io_x[8] ? _GEN21341 : _GEN21340;
wire  _GEN21343 = io_x[12] ? _GEN21342 : _GEN21339;
wire  _GEN21344 = io_x[0] ? _GEN21343 : _GEN21336;
wire  _GEN21345 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21346 = 1'b0;
wire  _GEN21347 = io_x[8] ? _GEN21346 : _GEN21345;
wire  _GEN21348 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21349 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21350 = io_x[8] ? _GEN21349 : _GEN21348;
wire  _GEN21351 = io_x[12] ? _GEN21350 : _GEN21347;
wire  _GEN21352 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21353 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21354 = io_x[8] ? _GEN21353 : _GEN21352;
wire  _GEN21355 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21356 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21357 = io_x[8] ? _GEN21356 : _GEN21355;
wire  _GEN21358 = io_x[12] ? _GEN21357 : _GEN21354;
wire  _GEN21359 = io_x[0] ? _GEN21358 : _GEN21351;
wire  _GEN21360 = io_x[32] ? _GEN21359 : _GEN21344;
wire  _GEN21361 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21362 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21363 = io_x[8] ? _GEN21362 : _GEN21361;
wire  _GEN21364 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21365 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21366 = io_x[8] ? _GEN21365 : _GEN21364;
wire  _GEN21367 = io_x[12] ? _GEN21366 : _GEN21363;
wire  _GEN21368 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21369 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21370 = io_x[8] ? _GEN21369 : _GEN21368;
wire  _GEN21371 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21372 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21373 = io_x[8] ? _GEN21372 : _GEN21371;
wire  _GEN21374 = io_x[12] ? _GEN21373 : _GEN21370;
wire  _GEN21375 = io_x[0] ? _GEN21374 : _GEN21367;
wire  _GEN21376 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21377 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21378 = io_x[8] ? _GEN21377 : _GEN21376;
wire  _GEN21379 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21380 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21381 = io_x[8] ? _GEN21380 : _GEN21379;
wire  _GEN21382 = io_x[12] ? _GEN21381 : _GEN21378;
wire  _GEN21383 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21384 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21385 = io_x[8] ? _GEN21384 : _GEN21383;
wire  _GEN21386 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21387 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21388 = io_x[8] ? _GEN21387 : _GEN21386;
wire  _GEN21389 = io_x[12] ? _GEN21388 : _GEN21385;
wire  _GEN21390 = io_x[0] ? _GEN21389 : _GEN21382;
wire  _GEN21391 = io_x[32] ? _GEN21390 : _GEN21375;
wire  _GEN21392 = io_x[42] ? _GEN21391 : _GEN21360;
wire  _GEN21393 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21394 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21395 = io_x[8] ? _GEN21394 : _GEN21393;
wire  _GEN21396 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21397 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21398 = io_x[8] ? _GEN21397 : _GEN21396;
wire  _GEN21399 = io_x[12] ? _GEN21398 : _GEN21395;
wire  _GEN21400 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21401 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21402 = io_x[8] ? _GEN21401 : _GEN21400;
wire  _GEN21403 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21404 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21405 = io_x[8] ? _GEN21404 : _GEN21403;
wire  _GEN21406 = io_x[12] ? _GEN21405 : _GEN21402;
wire  _GEN21407 = io_x[0] ? _GEN21406 : _GEN21399;
wire  _GEN21408 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21409 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21410 = io_x[8] ? _GEN21409 : _GEN21408;
wire  _GEN21411 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21412 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21413 = io_x[8] ? _GEN21412 : _GEN21411;
wire  _GEN21414 = io_x[12] ? _GEN21413 : _GEN21410;
wire  _GEN21415 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21416 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21417 = io_x[8] ? _GEN21416 : _GEN21415;
wire  _GEN21418 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21419 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21420 = io_x[8] ? _GEN21419 : _GEN21418;
wire  _GEN21421 = io_x[12] ? _GEN21420 : _GEN21417;
wire  _GEN21422 = io_x[0] ? _GEN21421 : _GEN21414;
wire  _GEN21423 = io_x[32] ? _GEN21422 : _GEN21407;
wire  _GEN21424 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21425 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21426 = io_x[8] ? _GEN21425 : _GEN21424;
wire  _GEN21427 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21428 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21429 = io_x[8] ? _GEN21428 : _GEN21427;
wire  _GEN21430 = io_x[12] ? _GEN21429 : _GEN21426;
wire  _GEN21431 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21432 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21433 = io_x[8] ? _GEN21432 : _GEN21431;
wire  _GEN21434 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21435 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21436 = io_x[8] ? _GEN21435 : _GEN21434;
wire  _GEN21437 = io_x[12] ? _GEN21436 : _GEN21433;
wire  _GEN21438 = io_x[0] ? _GEN21437 : _GEN21430;
wire  _GEN21439 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21440 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21441 = io_x[8] ? _GEN21440 : _GEN21439;
wire  _GEN21442 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21443 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21444 = io_x[8] ? _GEN21443 : _GEN21442;
wire  _GEN21445 = io_x[12] ? _GEN21444 : _GEN21441;
wire  _GEN21446 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21447 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21448 = io_x[8] ? _GEN21447 : _GEN21446;
wire  _GEN21449 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21450 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21451 = io_x[8] ? _GEN21450 : _GEN21449;
wire  _GEN21452 = io_x[12] ? _GEN21451 : _GEN21448;
wire  _GEN21453 = io_x[0] ? _GEN21452 : _GEN21445;
wire  _GEN21454 = io_x[32] ? _GEN21453 : _GEN21438;
wire  _GEN21455 = io_x[42] ? _GEN21454 : _GEN21423;
wire  _GEN21456 = io_x[69] ? _GEN21455 : _GEN21392;
wire  _GEN21457 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21458 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21459 = io_x[8] ? _GEN21458 : _GEN21457;
wire  _GEN21460 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21461 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21462 = io_x[8] ? _GEN21461 : _GEN21460;
wire  _GEN21463 = io_x[12] ? _GEN21462 : _GEN21459;
wire  _GEN21464 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21465 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21466 = io_x[8] ? _GEN21465 : _GEN21464;
wire  _GEN21467 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21468 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21469 = io_x[8] ? _GEN21468 : _GEN21467;
wire  _GEN21470 = io_x[12] ? _GEN21469 : _GEN21466;
wire  _GEN21471 = io_x[0] ? _GEN21470 : _GEN21463;
wire  _GEN21472 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21473 = io_x[8] ? _GEN21346 : _GEN21472;
wire  _GEN21474 = 1'b1;
wire  _GEN21475 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21476 = io_x[8] ? _GEN21475 : _GEN21474;
wire  _GEN21477 = io_x[12] ? _GEN21476 : _GEN21473;
wire  _GEN21478 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21479 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21480 = io_x[8] ? _GEN21479 : _GEN21478;
wire  _GEN21481 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21482 = io_x[8] ? _GEN21481 : _GEN21474;
wire  _GEN21483 = io_x[12] ? _GEN21482 : _GEN21480;
wire  _GEN21484 = io_x[0] ? _GEN21483 : _GEN21477;
wire  _GEN21485 = io_x[32] ? _GEN21484 : _GEN21471;
wire  _GEN21486 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21487 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21488 = io_x[8] ? _GEN21487 : _GEN21486;
wire  _GEN21489 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21490 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21491 = io_x[8] ? _GEN21490 : _GEN21489;
wire  _GEN21492 = io_x[12] ? _GEN21491 : _GEN21488;
wire  _GEN21493 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21494 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21495 = io_x[8] ? _GEN21494 : _GEN21493;
wire  _GEN21496 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21497 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21498 = io_x[8] ? _GEN21497 : _GEN21496;
wire  _GEN21499 = io_x[12] ? _GEN21498 : _GEN21495;
wire  _GEN21500 = io_x[0] ? _GEN21499 : _GEN21492;
wire  _GEN21501 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21502 = io_x[8] ? _GEN21474 : _GEN21501;
wire  _GEN21503 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21504 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21505 = io_x[8] ? _GEN21504 : _GEN21503;
wire  _GEN21506 = io_x[12] ? _GEN21505 : _GEN21502;
wire  _GEN21507 = io_x[8] ? _GEN21474 : _GEN21346;
wire  _GEN21508 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21509 = io_x[8] ? _GEN21508 : _GEN21346;
wire  _GEN21510 = io_x[12] ? _GEN21509 : _GEN21507;
wire  _GEN21511 = io_x[0] ? _GEN21510 : _GEN21506;
wire  _GEN21512 = io_x[32] ? _GEN21511 : _GEN21500;
wire  _GEN21513 = io_x[42] ? _GEN21512 : _GEN21485;
wire  _GEN21514 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21515 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21516 = io_x[8] ? _GEN21515 : _GEN21514;
wire  _GEN21517 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21518 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21519 = io_x[8] ? _GEN21518 : _GEN21517;
wire  _GEN21520 = io_x[12] ? _GEN21519 : _GEN21516;
wire  _GEN21521 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21522 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21523 = io_x[8] ? _GEN21522 : _GEN21521;
wire  _GEN21524 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21525 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21526 = io_x[8] ? _GEN21525 : _GEN21524;
wire  _GEN21527 = io_x[12] ? _GEN21526 : _GEN21523;
wire  _GEN21528 = io_x[0] ? _GEN21527 : _GEN21520;
wire  _GEN21529 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21530 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21531 = io_x[8] ? _GEN21530 : _GEN21529;
wire  _GEN21532 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21533 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21534 = io_x[8] ? _GEN21533 : _GEN21532;
wire  _GEN21535 = io_x[12] ? _GEN21534 : _GEN21531;
wire  _GEN21536 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21537 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21538 = io_x[8] ? _GEN21537 : _GEN21536;
wire  _GEN21539 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21540 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21541 = io_x[8] ? _GEN21540 : _GEN21539;
wire  _GEN21542 = io_x[12] ? _GEN21541 : _GEN21538;
wire  _GEN21543 = io_x[0] ? _GEN21542 : _GEN21535;
wire  _GEN21544 = io_x[32] ? _GEN21543 : _GEN21528;
wire  _GEN21545 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21546 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21547 = io_x[8] ? _GEN21546 : _GEN21545;
wire  _GEN21548 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21549 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21550 = io_x[8] ? _GEN21549 : _GEN21548;
wire  _GEN21551 = io_x[12] ? _GEN21550 : _GEN21547;
wire  _GEN21552 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21553 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21554 = io_x[8] ? _GEN21553 : _GEN21552;
wire  _GEN21555 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21556 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21557 = io_x[8] ? _GEN21556 : _GEN21555;
wire  _GEN21558 = io_x[12] ? _GEN21557 : _GEN21554;
wire  _GEN21559 = io_x[0] ? _GEN21558 : _GEN21551;
wire  _GEN21560 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21561 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21562 = io_x[8] ? _GEN21561 : _GEN21560;
wire  _GEN21563 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21564 = io_x[4] ? _GEN21328 : _GEN21329;
wire  _GEN21565 = io_x[8] ? _GEN21564 : _GEN21563;
wire  _GEN21566 = io_x[12] ? _GEN21565 : _GEN21562;
wire  _GEN21567 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21568 = io_x[8] ? _GEN21346 : _GEN21567;
wire  _GEN21569 = io_x[4] ? _GEN21329 : _GEN21328;
wire  _GEN21570 = io_x[8] ? _GEN21569 : _GEN21346;
wire  _GEN21571 = io_x[12] ? _GEN21570 : _GEN21568;
wire  _GEN21572 = io_x[0] ? _GEN21571 : _GEN21566;
wire  _GEN21573 = io_x[32] ? _GEN21572 : _GEN21559;
wire  _GEN21574 = io_x[42] ? _GEN21573 : _GEN21544;
wire  _GEN21575 = io_x[69] ? _GEN21574 : _GEN21513;
wire  _GEN21576 = io_x[75] ? _GEN21575 : _GEN21456;
assign io_y[6] = _GEN21576;
wire  _GEN21577 = 1'b0;
wire  _GEN21578 = 1'b1;
wire  _GEN21579 = io_x[41] ? _GEN21578 : _GEN21577;
wire  _GEN21580 = io_x[41] ? _GEN21578 : _GEN21577;
wire  _GEN21581 = io_x[40] ? _GEN21580 : _GEN21579;
wire  _GEN21582 = io_x[41] ? _GEN21578 : _GEN21577;
wire  _GEN21583 = io_x[41] ? _GEN21578 : _GEN21577;
wire  _GEN21584 = io_x[40] ? _GEN21583 : _GEN21582;
wire  _GEN21585 = io_x[38] ? _GEN21584 : _GEN21581;
assign io_y[5] = _GEN21585;
wire  _GEN21586 = 1'b0;
wire  _GEN21587 = 1'b1;
wire  _GEN21588 = io_x[40] ? _GEN21587 : _GEN21586;
wire  _GEN21589 = io_x[40] ? _GEN21587 : _GEN21586;
wire  _GEN21590 = io_x[38] ? _GEN21589 : _GEN21588;
wire  _GEN21591 = io_x[40] ? _GEN21587 : _GEN21586;
wire  _GEN21592 = io_x[40] ? _GEN21587 : _GEN21586;
wire  _GEN21593 = io_x[38] ? _GEN21592 : _GEN21591;
wire  _GEN21594 = io_x[37] ? _GEN21593 : _GEN21590;
wire  _GEN21595 = io_x[40] ? _GEN21587 : _GEN21586;
wire  _GEN21596 = io_x[40] ? _GEN21587 : _GEN21586;
wire  _GEN21597 = io_x[38] ? _GEN21596 : _GEN21595;
wire  _GEN21598 = io_x[40] ? _GEN21587 : _GEN21586;
wire  _GEN21599 = io_x[40] ? _GEN21587 : _GEN21586;
wire  _GEN21600 = io_x[38] ? _GEN21599 : _GEN21598;
wire  _GEN21601 = io_x[37] ? _GEN21600 : _GEN21597;
wire  _GEN21602 = io_x[4] ? _GEN21601 : _GEN21594;
assign io_y[4] = _GEN21602;
wire  _GEN21603 = 1'b0;
wire  _GEN21604 = 1'b1;
wire  _GEN21605 = io_x[39] ? _GEN21604 : _GEN21603;
wire  _GEN21606 = io_x[39] ? _GEN21604 : _GEN21603;
wire  _GEN21607 = io_x[76] ? _GEN21606 : _GEN21605;
assign io_y[3] = _GEN21607;
wire  _GEN21608 = 1'b0;
wire  _GEN21609 = 1'b1;
wire  _GEN21610 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21611 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21612 = io_x[44] ? _GEN21611 : _GEN21610;
wire  _GEN21613 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21614 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21615 = io_x[44] ? _GEN21614 : _GEN21613;
wire  _GEN21616 = io_x[80] ? _GEN21615 : _GEN21612;
wire  _GEN21617 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21618 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21619 = io_x[44] ? _GEN21618 : _GEN21617;
wire  _GEN21620 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21621 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21622 = io_x[44] ? _GEN21621 : _GEN21620;
wire  _GEN21623 = io_x[80] ? _GEN21622 : _GEN21619;
wire  _GEN21624 = io_x[28] ? _GEN21623 : _GEN21616;
wire  _GEN21625 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21626 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21627 = io_x[44] ? _GEN21626 : _GEN21625;
wire  _GEN21628 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21629 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21630 = io_x[44] ? _GEN21629 : _GEN21628;
wire  _GEN21631 = io_x[80] ? _GEN21630 : _GEN21627;
wire  _GEN21632 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21633 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21634 = io_x[44] ? _GEN21633 : _GEN21632;
wire  _GEN21635 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21636 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21637 = io_x[44] ? _GEN21636 : _GEN21635;
wire  _GEN21638 = io_x[80] ? _GEN21637 : _GEN21634;
wire  _GEN21639 = io_x[28] ? _GEN21638 : _GEN21631;
wire  _GEN21640 = io_x[32] ? _GEN21639 : _GEN21624;
wire  _GEN21641 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21642 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21643 = io_x[44] ? _GEN21642 : _GEN21641;
wire  _GEN21644 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21645 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21646 = io_x[44] ? _GEN21645 : _GEN21644;
wire  _GEN21647 = io_x[80] ? _GEN21646 : _GEN21643;
wire  _GEN21648 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21649 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21650 = io_x[44] ? _GEN21649 : _GEN21648;
wire  _GEN21651 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21652 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21653 = io_x[44] ? _GEN21652 : _GEN21651;
wire  _GEN21654 = io_x[80] ? _GEN21653 : _GEN21650;
wire  _GEN21655 = io_x[28] ? _GEN21654 : _GEN21647;
wire  _GEN21656 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21657 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21658 = io_x[44] ? _GEN21657 : _GEN21656;
wire  _GEN21659 = 1'b1;
wire  _GEN21660 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21661 = io_x[44] ? _GEN21660 : _GEN21659;
wire  _GEN21662 = io_x[80] ? _GEN21661 : _GEN21658;
wire  _GEN21663 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21664 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21665 = io_x[44] ? _GEN21664 : _GEN21663;
wire  _GEN21666 = 1'b0;
wire  _GEN21667 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21668 = io_x[44] ? _GEN21667 : _GEN21666;
wire  _GEN21669 = io_x[80] ? _GEN21668 : _GEN21665;
wire  _GEN21670 = io_x[28] ? _GEN21669 : _GEN21662;
wire  _GEN21671 = io_x[32] ? _GEN21670 : _GEN21655;
wire  _GEN21672 = io_x[46] ? _GEN21671 : _GEN21640;
wire  _GEN21673 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21674 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21675 = io_x[44] ? _GEN21674 : _GEN21673;
wire  _GEN21676 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21677 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21678 = io_x[44] ? _GEN21677 : _GEN21676;
wire  _GEN21679 = io_x[80] ? _GEN21678 : _GEN21675;
wire  _GEN21680 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21681 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21682 = io_x[44] ? _GEN21681 : _GEN21680;
wire  _GEN21683 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21684 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21685 = io_x[44] ? _GEN21684 : _GEN21683;
wire  _GEN21686 = io_x[80] ? _GEN21685 : _GEN21682;
wire  _GEN21687 = io_x[28] ? _GEN21686 : _GEN21679;
wire  _GEN21688 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21689 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21690 = io_x[44] ? _GEN21689 : _GEN21688;
wire  _GEN21691 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21692 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21693 = io_x[44] ? _GEN21692 : _GEN21691;
wire  _GEN21694 = io_x[80] ? _GEN21693 : _GEN21690;
wire  _GEN21695 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21696 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21697 = io_x[44] ? _GEN21696 : _GEN21695;
wire  _GEN21698 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21699 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21700 = io_x[44] ? _GEN21699 : _GEN21698;
wire  _GEN21701 = io_x[80] ? _GEN21700 : _GEN21697;
wire  _GEN21702 = io_x[28] ? _GEN21701 : _GEN21694;
wire  _GEN21703 = io_x[32] ? _GEN21702 : _GEN21687;
wire  _GEN21704 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21705 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21706 = io_x[44] ? _GEN21705 : _GEN21704;
wire  _GEN21707 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21708 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21709 = io_x[44] ? _GEN21708 : _GEN21707;
wire  _GEN21710 = io_x[80] ? _GEN21709 : _GEN21706;
wire  _GEN21711 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21712 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21713 = io_x[44] ? _GEN21712 : _GEN21711;
wire  _GEN21714 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21715 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21716 = io_x[44] ? _GEN21715 : _GEN21714;
wire  _GEN21717 = io_x[80] ? _GEN21716 : _GEN21713;
wire  _GEN21718 = io_x[28] ? _GEN21717 : _GEN21710;
wire  _GEN21719 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21720 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21721 = io_x[44] ? _GEN21720 : _GEN21719;
wire  _GEN21722 = io_x[44] ? _GEN21659 : _GEN21666;
wire  _GEN21723 = io_x[80] ? _GEN21722 : _GEN21721;
wire  _GEN21724 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21725 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21726 = io_x[44] ? _GEN21725 : _GEN21724;
wire  _GEN21727 = io_x[38] ? _GEN21609 : _GEN21608;
wire  _GEN21728 = io_x[44] ? _GEN21659 : _GEN21727;
wire  _GEN21729 = io_x[80] ? _GEN21728 : _GEN21726;
wire  _GEN21730 = io_x[28] ? _GEN21729 : _GEN21723;
wire  _GEN21731 = io_x[32] ? _GEN21730 : _GEN21718;
wire  _GEN21732 = io_x[46] ? _GEN21731 : _GEN21703;
wire  _GEN21733 = io_x[41] ? _GEN21732 : _GEN21672;
assign io_y[2] = _GEN21733;
wire  _GEN21734 = 1'b0;
wire  _GEN21735 = 1'b1;
wire  _GEN21736 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21737 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21738 = io_x[27] ? _GEN21737 : _GEN21736;
wire  _GEN21739 = 1'b1;
wire  _GEN21740 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21741 = io_x[27] ? _GEN21740 : _GEN21739;
wire  _GEN21742 = io_x[29] ? _GEN21741 : _GEN21738;
wire  _GEN21743 = 1'b1;
wire  _GEN21744 = 1'b0;
wire  _GEN21745 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN21746 = io_x[75] ? _GEN21745 : _GEN21742;
wire  _GEN21747 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21748 = io_x[27] ? _GEN21747 : _GEN21739;
wire  _GEN21749 = io_x[29] ? _GEN21748 : _GEN21744;
wire  _GEN21750 = 1'b0;
wire  _GEN21751 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN21752 = io_x[29] ? _GEN21743 : _GEN21751;
wire  _GEN21753 = io_x[75] ? _GEN21752 : _GEN21749;
wire  _GEN21754 = io_x[38] ? _GEN21753 : _GEN21746;
wire  _GEN21755 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21756 = io_x[27] ? _GEN21739 : _GEN21755;
wire  _GEN21757 = io_x[29] ? _GEN21743 : _GEN21756;
wire  _GEN21758 = 1'b1;
wire  _GEN21759 = io_x[75] ? _GEN21758 : _GEN21757;
wire  _GEN21760 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21761 = io_x[27] ? _GEN21750 : _GEN21760;
wire  _GEN21762 = io_x[29] ? _GEN21744 : _GEN21761;
wire  _GEN21763 = io_x[75] ? _GEN21758 : _GEN21762;
wire  _GEN21764 = io_x[38] ? _GEN21763 : _GEN21759;
wire  _GEN21765 = io_x[34] ? _GEN21764 : _GEN21754;
wire  _GEN21766 = 1'b0;
wire  _GEN21767 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21768 = io_x[27] ? _GEN21739 : _GEN21767;
wire  _GEN21769 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21770 = io_x[27] ? _GEN21769 : _GEN21739;
wire  _GEN21771 = io_x[29] ? _GEN21770 : _GEN21768;
wire  _GEN21772 = 1'b0;
wire  _GEN21773 = io_x[75] ? _GEN21772 : _GEN21771;
wire  _GEN21774 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN21775 = io_x[38] ? _GEN21774 : _GEN21773;
wire  _GEN21776 = io_x[34] ? _GEN21775 : _GEN21766;
wire  _GEN21777 = io_x[39] ? _GEN21776 : _GEN21765;
wire  _GEN21778 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21779 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21780 = io_x[27] ? _GEN21779 : _GEN21778;
wire  _GEN21781 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21782 = io_x[27] ? _GEN21750 : _GEN21781;
wire  _GEN21783 = io_x[29] ? _GEN21782 : _GEN21780;
wire  _GEN21784 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21785 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21786 = io_x[27] ? _GEN21785 : _GEN21784;
wire  _GEN21787 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21788 = io_x[27] ? _GEN21787 : _GEN21750;
wire  _GEN21789 = io_x[29] ? _GEN21788 : _GEN21786;
wire  _GEN21790 = io_x[75] ? _GEN21789 : _GEN21783;
wire  _GEN21791 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21792 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21793 = io_x[27] ? _GEN21792 : _GEN21791;
wire  _GEN21794 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21795 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21796 = io_x[27] ? _GEN21795 : _GEN21794;
wire  _GEN21797 = io_x[29] ? _GEN21796 : _GEN21793;
wire  _GEN21798 = io_x[75] ? _GEN21758 : _GEN21797;
wire  _GEN21799 = io_x[38] ? _GEN21798 : _GEN21790;
wire  _GEN21800 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21801 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21802 = io_x[27] ? _GEN21801 : _GEN21800;
wire  _GEN21803 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21804 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21805 = io_x[27] ? _GEN21804 : _GEN21803;
wire  _GEN21806 = io_x[29] ? _GEN21805 : _GEN21802;
wire  _GEN21807 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21808 = io_x[27] ? _GEN21807 : _GEN21739;
wire  _GEN21809 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21810 = io_x[27] ? _GEN21809 : _GEN21739;
wire  _GEN21811 = io_x[29] ? _GEN21810 : _GEN21808;
wire  _GEN21812 = io_x[75] ? _GEN21811 : _GEN21806;
wire  _GEN21813 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21814 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21815 = io_x[27] ? _GEN21814 : _GEN21813;
wire  _GEN21816 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21817 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21818 = io_x[27] ? _GEN21817 : _GEN21816;
wire  _GEN21819 = io_x[29] ? _GEN21818 : _GEN21815;
wire  _GEN21820 = io_x[75] ? _GEN21758 : _GEN21819;
wire  _GEN21821 = io_x[38] ? _GEN21820 : _GEN21812;
wire  _GEN21822 = io_x[34] ? _GEN21821 : _GEN21799;
wire  _GEN21823 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN21824 = io_x[29] ? _GEN21743 : _GEN21823;
wire  _GEN21825 = io_x[75] ? _GEN21758 : _GEN21824;
wire  _GEN21826 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21827 = io_x[27] ? _GEN21750 : _GEN21826;
wire  _GEN21828 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21829 = io_x[27] ? _GEN21750 : _GEN21828;
wire  _GEN21830 = io_x[29] ? _GEN21829 : _GEN21827;
wire  _GEN21831 = io_x[75] ? _GEN21830 : _GEN21758;
wire  _GEN21832 = io_x[38] ? _GEN21831 : _GEN21825;
wire  _GEN21833 = 1'b1;
wire  _GEN21834 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21835 = io_x[27] ? _GEN21834 : _GEN21739;
wire  _GEN21836 = io_x[29] ? _GEN21743 : _GEN21835;
wire  _GEN21837 = io_x[75] ? _GEN21836 : _GEN21758;
wire  _GEN21838 = io_x[38] ? _GEN21837 : _GEN21833;
wire  _GEN21839 = io_x[34] ? _GEN21838 : _GEN21832;
wire  _GEN21840 = io_x[39] ? _GEN21839 : _GEN21822;
wire  _GEN21841 = io_x[46] ? _GEN21840 : _GEN21777;
wire  _GEN21842 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN21843 = io_x[75] ? _GEN21842 : _GEN21758;
wire  _GEN21844 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21845 = io_x[27] ? _GEN21750 : _GEN21844;
wire  _GEN21846 = io_x[29] ? _GEN21744 : _GEN21845;
wire  _GEN21847 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21848 = io_x[27] ? _GEN21739 : _GEN21847;
wire  _GEN21849 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21850 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21851 = io_x[27] ? _GEN21850 : _GEN21849;
wire  _GEN21852 = io_x[29] ? _GEN21851 : _GEN21848;
wire  _GEN21853 = io_x[75] ? _GEN21852 : _GEN21846;
wire  _GEN21854 = io_x[38] ? _GEN21853 : _GEN21843;
wire  _GEN21855 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN21856 = io_x[75] ? _GEN21758 : _GEN21855;
wire  _GEN21857 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21858 = io_x[27] ? _GEN21750 : _GEN21857;
wire  _GEN21859 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN21860 = io_x[29] ? _GEN21859 : _GEN21858;
wire  _GEN21861 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21862 = io_x[27] ? _GEN21739 : _GEN21861;
wire  _GEN21863 = io_x[29] ? _GEN21743 : _GEN21862;
wire  _GEN21864 = io_x[75] ? _GEN21863 : _GEN21860;
wire  _GEN21865 = io_x[38] ? _GEN21864 : _GEN21856;
wire  _GEN21866 = io_x[34] ? _GEN21865 : _GEN21854;
wire  _GEN21867 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21868 = io_x[27] ? _GEN21867 : _GEN21739;
wire  _GEN21869 = io_x[29] ? _GEN21868 : _GEN21744;
wire  _GEN21870 = io_x[75] ? _GEN21772 : _GEN21869;
wire  _GEN21871 = 1'b0;
wire  _GEN21872 = io_x[38] ? _GEN21871 : _GEN21870;
wire  _GEN21873 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21874 = io_x[27] ? _GEN21739 : _GEN21873;
wire  _GEN21875 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21876 = io_x[27] ? _GEN21875 : _GEN21739;
wire  _GEN21877 = io_x[29] ? _GEN21876 : _GEN21874;
wire  _GEN21878 = io_x[75] ? _GEN21772 : _GEN21877;
wire  _GEN21879 = io_x[38] ? _GEN21833 : _GEN21878;
wire  _GEN21880 = io_x[34] ? _GEN21879 : _GEN21872;
wire  _GEN21881 = io_x[39] ? _GEN21880 : _GEN21866;
wire  _GEN21882 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21883 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21884 = io_x[27] ? _GEN21883 : _GEN21882;
wire  _GEN21885 = io_x[29] ? _GEN21884 : _GEN21743;
wire  _GEN21886 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21887 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21888 = io_x[27] ? _GEN21887 : _GEN21886;
wire  _GEN21889 = io_x[29] ? _GEN21743 : _GEN21888;
wire  _GEN21890 = io_x[75] ? _GEN21889 : _GEN21885;
wire  _GEN21891 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21892 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21893 = io_x[27] ? _GEN21892 : _GEN21891;
wire  _GEN21894 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21895 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21896 = io_x[27] ? _GEN21895 : _GEN21894;
wire  _GEN21897 = io_x[29] ? _GEN21896 : _GEN21893;
wire  _GEN21898 = io_x[75] ? _GEN21758 : _GEN21897;
wire  _GEN21899 = io_x[38] ? _GEN21898 : _GEN21890;
wire  _GEN21900 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21901 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21902 = io_x[27] ? _GEN21901 : _GEN21900;
wire  _GEN21903 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21904 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21905 = io_x[27] ? _GEN21904 : _GEN21903;
wire  _GEN21906 = io_x[29] ? _GEN21905 : _GEN21902;
wire  _GEN21907 = io_x[75] ? _GEN21758 : _GEN21906;
wire  _GEN21908 = io_x[38] ? _GEN21833 : _GEN21907;
wire  _GEN21909 = io_x[34] ? _GEN21908 : _GEN21899;
wire  _GEN21910 = 1'b1;
wire  _GEN21911 = io_x[39] ? _GEN21910 : _GEN21909;
wire  _GEN21912 = io_x[46] ? _GEN21911 : _GEN21881;
wire  _GEN21913 = io_x[18] ? _GEN21912 : _GEN21841;
wire  _GEN21914 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21915 = io_x[27] ? _GEN21739 : _GEN21914;
wire  _GEN21916 = io_x[29] ? _GEN21743 : _GEN21915;
wire  _GEN21917 = io_x[75] ? _GEN21758 : _GEN21916;
wire  _GEN21918 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN21919 = io_x[75] ? _GEN21758 : _GEN21918;
wire  _GEN21920 = io_x[38] ? _GEN21919 : _GEN21917;
wire  _GEN21921 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21922 = io_x[27] ? _GEN21739 : _GEN21921;
wire  _GEN21923 = io_x[29] ? _GEN21743 : _GEN21922;
wire  _GEN21924 = io_x[75] ? _GEN21923 : _GEN21772;
wire  _GEN21925 = io_x[38] ? _GEN21833 : _GEN21924;
wire  _GEN21926 = io_x[34] ? _GEN21925 : _GEN21920;
wire  _GEN21927 = 1'b1;
wire  _GEN21928 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN21929 = io_x[75] ? _GEN21928 : _GEN21758;
wire  _GEN21930 = io_x[38] ? _GEN21833 : _GEN21929;
wire  _GEN21931 = io_x[34] ? _GEN21930 : _GEN21927;
wire  _GEN21932 = io_x[39] ? _GEN21931 : _GEN21926;
wire  _GEN21933 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21934 = io_x[27] ? _GEN21739 : _GEN21933;
wire  _GEN21935 = io_x[29] ? _GEN21743 : _GEN21934;
wire  _GEN21936 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21937 = io_x[27] ? _GEN21739 : _GEN21936;
wire  _GEN21938 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21939 = io_x[27] ? _GEN21739 : _GEN21938;
wire  _GEN21940 = io_x[29] ? _GEN21939 : _GEN21937;
wire  _GEN21941 = io_x[75] ? _GEN21940 : _GEN21935;
wire  _GEN21942 = io_x[38] ? _GEN21871 : _GEN21941;
wire  _GEN21943 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21944 = io_x[27] ? _GEN21739 : _GEN21943;
wire  _GEN21945 = io_x[29] ? _GEN21743 : _GEN21944;
wire  _GEN21946 = io_x[75] ? _GEN21758 : _GEN21945;
wire  _GEN21947 = io_x[38] ? _GEN21833 : _GEN21946;
wire  _GEN21948 = io_x[34] ? _GEN21947 : _GEN21942;
wire  _GEN21949 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN21950 = io_x[38] ? _GEN21833 : _GEN21949;
wire  _GEN21951 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21952 = io_x[27] ? _GEN21739 : _GEN21951;
wire  _GEN21953 = io_x[29] ? _GEN21743 : _GEN21952;
wire  _GEN21954 = io_x[75] ? _GEN21953 : _GEN21758;
wire  _GEN21955 = io_x[38] ? _GEN21833 : _GEN21954;
wire  _GEN21956 = io_x[34] ? _GEN21955 : _GEN21950;
wire  _GEN21957 = io_x[39] ? _GEN21956 : _GEN21948;
wire  _GEN21958 = io_x[46] ? _GEN21957 : _GEN21932;
wire  _GEN21959 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN21960 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21961 = io_x[27] ? _GEN21739 : _GEN21960;
wire  _GEN21962 = io_x[29] ? _GEN21743 : _GEN21961;
wire  _GEN21963 = io_x[75] ? _GEN21758 : _GEN21962;
wire  _GEN21964 = io_x[38] ? _GEN21963 : _GEN21959;
wire  _GEN21965 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN21966 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21967 = io_x[27] ? _GEN21739 : _GEN21966;
wire  _GEN21968 = io_x[29] ? _GEN21743 : _GEN21967;
wire  _GEN21969 = io_x[75] ? _GEN21772 : _GEN21968;
wire  _GEN21970 = io_x[38] ? _GEN21969 : _GEN21965;
wire  _GEN21971 = io_x[34] ? _GEN21970 : _GEN21964;
wire  _GEN21972 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21973 = io_x[27] ? _GEN21739 : _GEN21972;
wire  _GEN21974 = io_x[29] ? _GEN21743 : _GEN21973;
wire  _GEN21975 = io_x[75] ? _GEN21974 : _GEN21758;
wire  _GEN21976 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN21977 = io_x[38] ? _GEN21976 : _GEN21975;
wire  _GEN21978 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21979 = io_x[27] ? _GEN21739 : _GEN21978;
wire  _GEN21980 = io_x[29] ? _GEN21744 : _GEN21979;
wire  _GEN21981 = io_x[75] ? _GEN21980 : _GEN21772;
wire  _GEN21982 = io_x[38] ? _GEN21871 : _GEN21981;
wire  _GEN21983 = io_x[34] ? _GEN21982 : _GEN21977;
wire  _GEN21984 = io_x[39] ? _GEN21983 : _GEN21971;
wire  _GEN21985 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN21986 = io_x[38] ? _GEN21871 : _GEN21985;
wire  _GEN21987 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21988 = io_x[27] ? _GEN21739 : _GEN21987;
wire  _GEN21989 = io_x[29] ? _GEN21743 : _GEN21988;
wire  _GEN21990 = io_x[75] ? _GEN21989 : _GEN21758;
wire  _GEN21991 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN21992 = io_x[38] ? _GEN21991 : _GEN21990;
wire  _GEN21993 = io_x[34] ? _GEN21992 : _GEN21986;
wire  _GEN21994 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN21995 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN21996 = io_x[27] ? _GEN21739 : _GEN21995;
wire  _GEN21997 = io_x[29] ? _GEN21743 : _GEN21996;
wire  _GEN21998 = io_x[75] ? _GEN21997 : _GEN21758;
wire  _GEN21999 = io_x[38] ? _GEN21998 : _GEN21994;
wire  _GEN22000 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22001 = io_x[27] ? _GEN21739 : _GEN22000;
wire  _GEN22002 = io_x[29] ? _GEN21743 : _GEN22001;
wire  _GEN22003 = io_x[75] ? _GEN22002 : _GEN21758;
wire  _GEN22004 = io_x[38] ? _GEN21833 : _GEN22003;
wire  _GEN22005 = io_x[34] ? _GEN22004 : _GEN21999;
wire  _GEN22006 = io_x[39] ? _GEN22005 : _GEN21993;
wire  _GEN22007 = io_x[46] ? _GEN22006 : _GEN21984;
wire  _GEN22008 = io_x[18] ? _GEN22007 : _GEN21958;
wire  _GEN22009 = io_x[49] ? _GEN22008 : _GEN21913;
wire  _GEN22010 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22011 = io_x[27] ? _GEN22010 : _GEN21739;
wire  _GEN22012 = io_x[29] ? _GEN22011 : _GEN21743;
wire  _GEN22013 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22014 = io_x[27] ? _GEN22013 : _GEN21739;
wire  _GEN22015 = io_x[29] ? _GEN22014 : _GEN21743;
wire  _GEN22016 = io_x[75] ? _GEN22015 : _GEN22012;
wire  _GEN22017 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22018 = io_x[27] ? _GEN22017 : _GEN21750;
wire  _GEN22019 = io_x[29] ? _GEN22018 : _GEN21743;
wire  _GEN22020 = io_x[75] ? _GEN21758 : _GEN22019;
wire  _GEN22021 = io_x[38] ? _GEN22020 : _GEN22016;
wire  _GEN22022 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22023 = io_x[27] ? _GEN21750 : _GEN22022;
wire  _GEN22024 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22025 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22026 = io_x[27] ? _GEN22025 : _GEN22024;
wire  _GEN22027 = io_x[29] ? _GEN22026 : _GEN22023;
wire  _GEN22028 = io_x[75] ? _GEN21758 : _GEN22027;
wire  _GEN22029 = io_x[38] ? _GEN22028 : _GEN21833;
wire  _GEN22030 = io_x[34] ? _GEN22029 : _GEN22021;
wire  _GEN22031 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22032 = io_x[27] ? _GEN21750 : _GEN22031;
wire  _GEN22033 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22034 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22035 = io_x[27] ? _GEN22034 : _GEN22033;
wire  _GEN22036 = io_x[29] ? _GEN22035 : _GEN22032;
wire  _GEN22037 = io_x[75] ? _GEN21772 : _GEN22036;
wire  _GEN22038 = io_x[38] ? _GEN21871 : _GEN22037;
wire  _GEN22039 = io_x[34] ? _GEN22038 : _GEN21766;
wire  _GEN22040 = io_x[39] ? _GEN22039 : _GEN22030;
wire  _GEN22041 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22042 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22043 = io_x[27] ? _GEN22042 : _GEN22041;
wire  _GEN22044 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22045 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22046 = io_x[27] ? _GEN22045 : _GEN22044;
wire  _GEN22047 = io_x[29] ? _GEN22046 : _GEN22043;
wire  _GEN22048 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22049 = io_x[27] ? _GEN21739 : _GEN22048;
wire  _GEN22050 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22051 = io_x[27] ? _GEN22050 : _GEN21739;
wire  _GEN22052 = io_x[29] ? _GEN22051 : _GEN22049;
wire  _GEN22053 = io_x[75] ? _GEN22052 : _GEN22047;
wire  _GEN22054 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22055 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22056 = io_x[27] ? _GEN22055 : _GEN22054;
wire  _GEN22057 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22058 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22059 = io_x[27] ? _GEN22058 : _GEN22057;
wire  _GEN22060 = io_x[29] ? _GEN22059 : _GEN22056;
wire  _GEN22061 = io_x[75] ? _GEN21758 : _GEN22060;
wire  _GEN22062 = io_x[38] ? _GEN22061 : _GEN22053;
wire  _GEN22063 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22064 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22065 = io_x[27] ? _GEN22064 : _GEN22063;
wire  _GEN22066 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22067 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22068 = io_x[27] ? _GEN22067 : _GEN22066;
wire  _GEN22069 = io_x[29] ? _GEN22068 : _GEN22065;
wire  _GEN22070 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22071 = io_x[27] ? _GEN22070 : _GEN21739;
wire  _GEN22072 = io_x[29] ? _GEN22071 : _GEN21743;
wire  _GEN22073 = io_x[75] ? _GEN22072 : _GEN22069;
wire  _GEN22074 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22075 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22076 = io_x[27] ? _GEN22075 : _GEN22074;
wire  _GEN22077 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22078 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22079 = io_x[27] ? _GEN22078 : _GEN22077;
wire  _GEN22080 = io_x[29] ? _GEN22079 : _GEN22076;
wire  _GEN22081 = io_x[75] ? _GEN21758 : _GEN22080;
wire  _GEN22082 = io_x[38] ? _GEN22081 : _GEN22073;
wire  _GEN22083 = io_x[34] ? _GEN22082 : _GEN22062;
wire  _GEN22084 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22085 = io_x[27] ? _GEN22084 : _GEN21750;
wire  _GEN22086 = io_x[29] ? _GEN22085 : _GEN21744;
wire  _GEN22087 = io_x[75] ? _GEN22086 : _GEN21758;
wire  _GEN22088 = io_x[38] ? _GEN22087 : _GEN21833;
wire  _GEN22089 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN22090 = io_x[29] ? _GEN22089 : _GEN21743;
wire  _GEN22091 = io_x[75] ? _GEN22090 : _GEN21758;
wire  _GEN22092 = io_x[38] ? _GEN22091 : _GEN21833;
wire  _GEN22093 = io_x[34] ? _GEN22092 : _GEN22088;
wire  _GEN22094 = io_x[39] ? _GEN22093 : _GEN22083;
wire  _GEN22095 = io_x[46] ? _GEN22094 : _GEN22040;
wire  _GEN22096 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22097 = io_x[27] ? _GEN22096 : _GEN21750;
wire  _GEN22098 = io_x[29] ? _GEN21743 : _GEN22097;
wire  _GEN22099 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22100 = io_x[27] ? _GEN22099 : _GEN21739;
wire  _GEN22101 = io_x[29] ? _GEN21743 : _GEN22100;
wire  _GEN22102 = io_x[75] ? _GEN22101 : _GEN22098;
wire  _GEN22103 = io_x[38] ? _GEN22102 : _GEN21833;
wire  _GEN22104 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22105 = io_x[27] ? _GEN21750 : _GEN22104;
wire  _GEN22106 = io_x[29] ? _GEN21744 : _GEN22105;
wire  _GEN22107 = io_x[75] ? _GEN21758 : _GEN22106;
wire  _GEN22108 = io_x[38] ? _GEN22107 : _GEN21833;
wire  _GEN22109 = io_x[34] ? _GEN22108 : _GEN22103;
wire  _GEN22110 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22111 = io_x[38] ? _GEN21871 : _GEN22110;
wire  _GEN22112 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22113 = io_x[27] ? _GEN21750 : _GEN22112;
wire  _GEN22114 = io_x[29] ? _GEN22113 : _GEN21743;
wire  _GEN22115 = io_x[75] ? _GEN21758 : _GEN22114;
wire  _GEN22116 = io_x[38] ? _GEN21833 : _GEN22115;
wire  _GEN22117 = io_x[34] ? _GEN22116 : _GEN22111;
wire  _GEN22118 = io_x[39] ? _GEN22117 : _GEN22109;
wire  _GEN22119 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22120 = io_x[27] ? _GEN22119 : _GEN21739;
wire  _GEN22121 = io_x[29] ? _GEN22120 : _GEN21743;
wire  _GEN22122 = io_x[75] ? _GEN21758 : _GEN22121;
wire  _GEN22123 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22124 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22125 = io_x[27] ? _GEN22124 : _GEN22123;
wire  _GEN22126 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22127 = io_x[27] ? _GEN21750 : _GEN22126;
wire  _GEN22128 = io_x[29] ? _GEN22127 : _GEN22125;
wire  _GEN22129 = io_x[75] ? _GEN21772 : _GEN22128;
wire  _GEN22130 = io_x[38] ? _GEN22129 : _GEN22122;
wire  _GEN22131 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22132 = io_x[27] ? _GEN21750 : _GEN22131;
wire  _GEN22133 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22134 = io_x[27] ? _GEN21739 : _GEN22133;
wire  _GEN22135 = io_x[29] ? _GEN22134 : _GEN22132;
wire  _GEN22136 = io_x[75] ? _GEN21758 : _GEN22135;
wire  _GEN22137 = io_x[38] ? _GEN21833 : _GEN22136;
wire  _GEN22138 = io_x[34] ? _GEN22137 : _GEN22130;
wire  _GEN22139 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22140 = io_x[38] ? _GEN22139 : _GEN21833;
wire  _GEN22141 = io_x[34] ? _GEN22140 : _GEN21927;
wire  _GEN22142 = io_x[39] ? _GEN22141 : _GEN22138;
wire  _GEN22143 = io_x[46] ? _GEN22142 : _GEN22118;
wire  _GEN22144 = io_x[18] ? _GEN22143 : _GEN22095;
wire  _GEN22145 = 1'b1;
wire  _GEN22146 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22147 = io_x[27] ? _GEN22146 : _GEN21750;
wire  _GEN22148 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22149 = io_x[27] ? _GEN21750 : _GEN22148;
wire  _GEN22150 = io_x[29] ? _GEN22149 : _GEN22147;
wire  _GEN22151 = io_x[75] ? _GEN22150 : _GEN21758;
wire  _GEN22152 = io_x[38] ? _GEN21871 : _GEN22151;
wire  _GEN22153 = io_x[34] ? _GEN21927 : _GEN22152;
wire  _GEN22154 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22155 = io_x[27] ? _GEN22154 : _GEN21739;
wire  _GEN22156 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22157 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22158 = io_x[27] ? _GEN22157 : _GEN22156;
wire  _GEN22159 = io_x[29] ? _GEN22158 : _GEN22155;
wire  _GEN22160 = io_x[75] ? _GEN22159 : _GEN21758;
wire  _GEN22161 = io_x[38] ? _GEN21833 : _GEN22160;
wire  _GEN22162 = io_x[34] ? _GEN22161 : _GEN21927;
wire  _GEN22163 = io_x[39] ? _GEN22162 : _GEN22153;
wire  _GEN22164 = io_x[46] ? _GEN22163 : _GEN22145;
wire  _GEN22165 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN22166 = io_x[34] ? _GEN22165 : _GEN21927;
wire  _GEN22167 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN22168 = io_x[38] ? _GEN22167 : _GEN21833;
wire  _GEN22169 = io_x[34] ? _GEN21766 : _GEN22168;
wire  _GEN22170 = io_x[39] ? _GEN22169 : _GEN22166;
wire  _GEN22171 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN22172 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN22173 = io_x[34] ? _GEN22172 : _GEN22171;
wire  _GEN22174 = io_x[39] ? _GEN21910 : _GEN22173;
wire  _GEN22175 = io_x[46] ? _GEN22174 : _GEN22170;
wire  _GEN22176 = io_x[18] ? _GEN22175 : _GEN22164;
wire  _GEN22177 = io_x[49] ? _GEN22176 : _GEN22144;
wire  _GEN22178 = io_x[24] ? _GEN22177 : _GEN22009;
wire  _GEN22179 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22180 = io_x[27] ? _GEN22179 : _GEN21750;
wire  _GEN22181 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22182 = io_x[27] ? _GEN22181 : _GEN21750;
wire  _GEN22183 = io_x[29] ? _GEN22182 : _GEN22180;
wire  _GEN22184 = io_x[75] ? _GEN21758 : _GEN22183;
wire  _GEN22185 = io_x[38] ? _GEN21833 : _GEN22184;
wire  _GEN22186 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN22187 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22188 = io_x[27] ? _GEN22187 : _GEN21750;
wire  _GEN22189 = io_x[29] ? _GEN22188 : _GEN21743;
wire  _GEN22190 = io_x[75] ? _GEN21758 : _GEN22189;
wire  _GEN22191 = io_x[38] ? _GEN22190 : _GEN22186;
wire  _GEN22192 = io_x[34] ? _GEN22191 : _GEN22185;
wire  _GEN22193 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN22194 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22195 = io_x[27] ? _GEN22194 : _GEN21750;
wire  _GEN22196 = io_x[29] ? _GEN22195 : _GEN22193;
wire  _GEN22197 = io_x[75] ? _GEN21772 : _GEN22196;
wire  _GEN22198 = io_x[38] ? _GEN22197 : _GEN21833;
wire  _GEN22199 = io_x[34] ? _GEN21927 : _GEN22198;
wire  _GEN22200 = io_x[39] ? _GEN22199 : _GEN22192;
wire  _GEN22201 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22202 = io_x[27] ? _GEN22201 : _GEN21739;
wire  _GEN22203 = io_x[29] ? _GEN22202 : _GEN21743;
wire  _GEN22204 = io_x[75] ? _GEN22203 : _GEN21758;
wire  _GEN22205 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22206 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22207 = io_x[27] ? _GEN22206 : _GEN22205;
wire  _GEN22208 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22209 = io_x[27] ? _GEN21739 : _GEN22208;
wire  _GEN22210 = io_x[29] ? _GEN22209 : _GEN22207;
wire  _GEN22211 = io_x[75] ? _GEN21772 : _GEN22210;
wire  _GEN22212 = io_x[38] ? _GEN22211 : _GEN22204;
wire  _GEN22213 = io_x[34] ? _GEN21766 : _GEN22212;
wire  _GEN22214 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22215 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22216 = io_x[27] ? _GEN22215 : _GEN22214;
wire  _GEN22217 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22218 = io_x[27] ? _GEN21739 : _GEN22217;
wire  _GEN22219 = io_x[29] ? _GEN22218 : _GEN22216;
wire  _GEN22220 = io_x[75] ? _GEN21758 : _GEN22219;
wire  _GEN22221 = io_x[38] ? _GEN21871 : _GEN22220;
wire  _GEN22222 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22223 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN22224 = io_x[38] ? _GEN22223 : _GEN22222;
wire  _GEN22225 = io_x[34] ? _GEN22224 : _GEN22221;
wire  _GEN22226 = io_x[39] ? _GEN22225 : _GEN22213;
wire  _GEN22227 = io_x[46] ? _GEN22226 : _GEN22200;
wire  _GEN22228 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22229 = io_x[27] ? _GEN21739 : _GEN22228;
wire  _GEN22230 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22231 = io_x[27] ? _GEN21750 : _GEN22230;
wire  _GEN22232 = io_x[29] ? _GEN22231 : _GEN22229;
wire  _GEN22233 = io_x[75] ? _GEN21772 : _GEN22232;
wire  _GEN22234 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22235 = io_x[27] ? _GEN21739 : _GEN22234;
wire  _GEN22236 = io_x[29] ? _GEN21743 : _GEN22235;
wire  _GEN22237 = io_x[75] ? _GEN21772 : _GEN22236;
wire  _GEN22238 = io_x[38] ? _GEN22237 : _GEN22233;
wire  _GEN22239 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22240 = io_x[27] ? _GEN21739 : _GEN22239;
wire  _GEN22241 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22242 = io_x[27] ? _GEN21750 : _GEN22241;
wire  _GEN22243 = io_x[29] ? _GEN22242 : _GEN22240;
wire  _GEN22244 = io_x[75] ? _GEN22243 : _GEN21772;
wire  _GEN22245 = io_x[38] ? _GEN21871 : _GEN22244;
wire  _GEN22246 = io_x[34] ? _GEN22245 : _GEN22238;
wire  _GEN22247 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22248 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN22249 = io_x[29] ? _GEN21744 : _GEN22248;
wire  _GEN22250 = io_x[75] ? _GEN21758 : _GEN22249;
wire  _GEN22251 = io_x[38] ? _GEN22250 : _GEN22247;
wire  _GEN22252 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN22253 = io_x[38] ? _GEN22252 : _GEN21871;
wire  _GEN22254 = io_x[34] ? _GEN22253 : _GEN22251;
wire  _GEN22255 = io_x[39] ? _GEN22254 : _GEN22246;
wire  _GEN22256 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22257 = io_x[27] ? _GEN21739 : _GEN22256;
wire  _GEN22258 = io_x[29] ? _GEN21743 : _GEN22257;
wire  _GEN22259 = io_x[75] ? _GEN22258 : _GEN21758;
wire  _GEN22260 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22261 = io_x[38] ? _GEN22260 : _GEN22259;
wire  _GEN22262 = io_x[34] ? _GEN21766 : _GEN22261;
wire  _GEN22263 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN22264 = io_x[34] ? _GEN22263 : _GEN21766;
wire  _GEN22265 = io_x[39] ? _GEN22264 : _GEN22262;
wire  _GEN22266 = io_x[46] ? _GEN22265 : _GEN22255;
wire  _GEN22267 = io_x[18] ? _GEN22266 : _GEN22227;
wire  _GEN22268 = 1'b0;
wire  _GEN22269 = io_x[49] ? _GEN22268 : _GEN22267;
wire  _GEN22270 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN22271 = io_x[38] ? _GEN21833 : _GEN22270;
wire  _GEN22272 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN22273 = io_x[34] ? _GEN22272 : _GEN22271;
wire  _GEN22274 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22275 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN22276 = io_x[38] ? _GEN22275 : _GEN22274;
wire  _GEN22277 = io_x[34] ? _GEN21927 : _GEN22276;
wire  _GEN22278 = io_x[39] ? _GEN22277 : _GEN22273;
wire  _GEN22279 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN22280 = io_x[75] ? _GEN22279 : _GEN21758;
wire  _GEN22281 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22282 = io_x[38] ? _GEN22281 : _GEN22280;
wire  _GEN22283 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22284 = io_x[27] ? _GEN22283 : _GEN21739;
wire  _GEN22285 = io_x[29] ? _GEN22284 : _GEN21744;
wire  _GEN22286 = io_x[75] ? _GEN21758 : _GEN22285;
wire  _GEN22287 = io_x[38] ? _GEN22286 : _GEN21871;
wire  _GEN22288 = io_x[34] ? _GEN22287 : _GEN22282;
wire  _GEN22289 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22290 = io_x[27] ? _GEN21750 : _GEN22289;
wire  _GEN22291 = io_x[29] ? _GEN21744 : _GEN22290;
wire  _GEN22292 = io_x[75] ? _GEN21772 : _GEN22291;
wire  _GEN22293 = io_x[38] ? _GEN21871 : _GEN22292;
wire  _GEN22294 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22295 = io_x[27] ? _GEN21739 : _GEN22294;
wire  _GEN22296 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN22297 = io_x[29] ? _GEN22296 : _GEN22295;
wire  _GEN22298 = io_x[75] ? _GEN21772 : _GEN22297;
wire  _GEN22299 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22300 = io_x[27] ? _GEN22299 : _GEN21750;
wire  _GEN22301 = io_x[29] ? _GEN22300 : _GEN21744;
wire  _GEN22302 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN22303 = io_x[75] ? _GEN22302 : _GEN22301;
wire  _GEN22304 = io_x[38] ? _GEN22303 : _GEN22298;
wire  _GEN22305 = io_x[34] ? _GEN22304 : _GEN22293;
wire  _GEN22306 = io_x[39] ? _GEN22305 : _GEN22288;
wire  _GEN22307 = io_x[46] ? _GEN22306 : _GEN22278;
wire  _GEN22308 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22309 = io_x[38] ? _GEN22308 : _GEN21833;
wire  _GEN22310 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN22311 = io_x[34] ? _GEN22310 : _GEN22309;
wire  _GEN22312 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN22313 = io_x[34] ? _GEN21766 : _GEN22312;
wire  _GEN22314 = io_x[39] ? _GEN22313 : _GEN22311;
wire  _GEN22315 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN22316 = io_x[29] ? _GEN21743 : _GEN22315;
wire  _GEN22317 = io_x[75] ? _GEN21758 : _GEN22316;
wire  _GEN22318 = io_x[38] ? _GEN22317 : _GEN21871;
wire  _GEN22319 = io_x[34] ? _GEN21766 : _GEN22318;
wire  _GEN22320 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN22321 = io_x[75] ? _GEN21758 : _GEN22320;
wire  _GEN22322 = io_x[38] ? _GEN22321 : _GEN21833;
wire  _GEN22323 = io_x[34] ? _GEN21766 : _GEN22322;
wire  _GEN22324 = io_x[39] ? _GEN22323 : _GEN22319;
wire  _GEN22325 = io_x[46] ? _GEN22324 : _GEN22314;
wire  _GEN22326 = io_x[18] ? _GEN22325 : _GEN22307;
wire  _GEN22327 = 1'b0;
wire  _GEN22328 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN22329 = io_x[46] ? _GEN22145 : _GEN22328;
wire  _GEN22330 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22331 = io_x[27] ? _GEN21739 : _GEN22330;
wire  _GEN22332 = io_x[29] ? _GEN22331 : _GEN21743;
wire  _GEN22333 = io_x[75] ? _GEN22332 : _GEN21758;
wire  _GEN22334 = io_x[38] ? _GEN22333 : _GEN21833;
wire  _GEN22335 = io_x[34] ? _GEN21927 : _GEN22334;
wire  _GEN22336 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN22337 = io_x[39] ? _GEN22336 : _GEN22335;
wire  _GEN22338 = io_x[46] ? _GEN22145 : _GEN22337;
wire  _GEN22339 = io_x[18] ? _GEN22338 : _GEN22329;
wire  _GEN22340 = io_x[49] ? _GEN22339 : _GEN22326;
wire  _GEN22341 = io_x[24] ? _GEN22340 : _GEN22269;
wire  _GEN22342 = io_x[80] ? _GEN22341 : _GEN22178;
wire  _GEN22343 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22344 = io_x[27] ? _GEN21739 : _GEN22343;
wire  _GEN22345 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22346 = io_x[27] ? _GEN22345 : _GEN21739;
wire  _GEN22347 = io_x[29] ? _GEN22346 : _GEN22344;
wire  _GEN22348 = io_x[75] ? _GEN21758 : _GEN22347;
wire  _GEN22349 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22350 = io_x[27] ? _GEN21739 : _GEN22349;
wire  _GEN22351 = io_x[29] ? _GEN21744 : _GEN22350;
wire  _GEN22352 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22353 = io_x[27] ? _GEN21739 : _GEN22352;
wire  _GEN22354 = io_x[29] ? _GEN21743 : _GEN22353;
wire  _GEN22355 = io_x[75] ? _GEN22354 : _GEN22351;
wire  _GEN22356 = io_x[38] ? _GEN22355 : _GEN22348;
wire  _GEN22357 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22358 = io_x[27] ? _GEN22357 : _GEN21739;
wire  _GEN22359 = io_x[29] ? _GEN22358 : _GEN21743;
wire  _GEN22360 = io_x[75] ? _GEN21758 : _GEN22359;
wire  _GEN22361 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22362 = io_x[27] ? _GEN21739 : _GEN22361;
wire  _GEN22363 = io_x[29] ? _GEN21744 : _GEN22362;
wire  _GEN22364 = io_x[75] ? _GEN21758 : _GEN22363;
wire  _GEN22365 = io_x[38] ? _GEN22364 : _GEN22360;
wire  _GEN22366 = io_x[34] ? _GEN22365 : _GEN22356;
wire  _GEN22367 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22368 = io_x[27] ? _GEN21750 : _GEN22367;
wire  _GEN22369 = io_x[29] ? _GEN21744 : _GEN22368;
wire  _GEN22370 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22371 = io_x[27] ? _GEN21739 : _GEN22370;
wire  _GEN22372 = io_x[29] ? _GEN21743 : _GEN22371;
wire  _GEN22373 = io_x[75] ? _GEN22372 : _GEN22369;
wire  _GEN22374 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22375 = io_x[27] ? _GEN21739 : _GEN22374;
wire  _GEN22376 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22377 = io_x[27] ? _GEN21750 : _GEN22376;
wire  _GEN22378 = io_x[29] ? _GEN22377 : _GEN22375;
wire  _GEN22379 = io_x[75] ? _GEN21772 : _GEN22378;
wire  _GEN22380 = io_x[38] ? _GEN22379 : _GEN22373;
wire  _GEN22381 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22382 = io_x[27] ? _GEN21739 : _GEN22381;
wire  _GEN22383 = io_x[29] ? _GEN21743 : _GEN22382;
wire  _GEN22384 = io_x[75] ? _GEN22383 : _GEN21758;
wire  _GEN22385 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22386 = io_x[27] ? _GEN21739 : _GEN22385;
wire  _GEN22387 = io_x[29] ? _GEN21743 : _GEN22386;
wire  _GEN22388 = io_x[75] ? _GEN22387 : _GEN21758;
wire  _GEN22389 = io_x[38] ? _GEN22388 : _GEN22384;
wire  _GEN22390 = io_x[34] ? _GEN22389 : _GEN22380;
wire  _GEN22391 = io_x[39] ? _GEN22390 : _GEN22366;
wire  _GEN22392 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22393 = io_x[27] ? _GEN21739 : _GEN22392;
wire  _GEN22394 = io_x[29] ? _GEN21743 : _GEN22393;
wire  _GEN22395 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22396 = io_x[27] ? _GEN21739 : _GEN22395;
wire  _GEN22397 = io_x[29] ? _GEN21743 : _GEN22396;
wire  _GEN22398 = io_x[75] ? _GEN22397 : _GEN22394;
wire  _GEN22399 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22400 = io_x[27] ? _GEN22399 : _GEN21739;
wire  _GEN22401 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22402 = io_x[27] ? _GEN21739 : _GEN22401;
wire  _GEN22403 = io_x[29] ? _GEN22402 : _GEN22400;
wire  _GEN22404 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22405 = io_x[27] ? _GEN21739 : _GEN22404;
wire  _GEN22406 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22407 = io_x[27] ? _GEN21739 : _GEN22406;
wire  _GEN22408 = io_x[29] ? _GEN22407 : _GEN22405;
wire  _GEN22409 = io_x[75] ? _GEN22408 : _GEN22403;
wire  _GEN22410 = io_x[38] ? _GEN22409 : _GEN22398;
wire  _GEN22411 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22412 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22413 = io_x[27] ? _GEN22412 : _GEN22411;
wire  _GEN22414 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22415 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22416 = io_x[27] ? _GEN22415 : _GEN22414;
wire  _GEN22417 = io_x[29] ? _GEN22416 : _GEN22413;
wire  _GEN22418 = io_x[75] ? _GEN21758 : _GEN22417;
wire  _GEN22419 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22420 = io_x[38] ? _GEN22419 : _GEN22418;
wire  _GEN22421 = io_x[34] ? _GEN22420 : _GEN22410;
wire  _GEN22422 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22423 = io_x[27] ? _GEN21739 : _GEN22422;
wire  _GEN22424 = io_x[29] ? _GEN21744 : _GEN22423;
wire  _GEN22425 = io_x[75] ? _GEN22424 : _GEN21758;
wire  _GEN22426 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22427 = io_x[27] ? _GEN21739 : _GEN22426;
wire  _GEN22428 = io_x[29] ? _GEN21744 : _GEN22427;
wire  _GEN22429 = io_x[75] ? _GEN22428 : _GEN21758;
wire  _GEN22430 = io_x[38] ? _GEN22429 : _GEN22425;
wire  _GEN22431 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22432 = io_x[27] ? _GEN21739 : _GEN22431;
wire  _GEN22433 = io_x[29] ? _GEN21743 : _GEN22432;
wire  _GEN22434 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22435 = io_x[27] ? _GEN21739 : _GEN22434;
wire  _GEN22436 = io_x[29] ? _GEN21743 : _GEN22435;
wire  _GEN22437 = io_x[75] ? _GEN22436 : _GEN22433;
wire  _GEN22438 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22439 = io_x[27] ? _GEN21739 : _GEN22438;
wire  _GEN22440 = io_x[29] ? _GEN21743 : _GEN22439;
wire  _GEN22441 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22442 = io_x[27] ? _GEN21739 : _GEN22441;
wire  _GEN22443 = io_x[29] ? _GEN22442 : _GEN21744;
wire  _GEN22444 = io_x[75] ? _GEN22443 : _GEN22440;
wire  _GEN22445 = io_x[38] ? _GEN22444 : _GEN22437;
wire  _GEN22446 = io_x[34] ? _GEN22445 : _GEN22430;
wire  _GEN22447 = io_x[39] ? _GEN22446 : _GEN22421;
wire  _GEN22448 = io_x[46] ? _GEN22447 : _GEN22391;
wire  _GEN22449 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22450 = io_x[27] ? _GEN21739 : _GEN22449;
wire  _GEN22451 = io_x[29] ? _GEN21743 : _GEN22450;
wire  _GEN22452 = io_x[75] ? _GEN22451 : _GEN21758;
wire  _GEN22453 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22454 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22455 = io_x[27] ? _GEN22454 : _GEN22453;
wire  _GEN22456 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22457 = io_x[27] ? _GEN21739 : _GEN22456;
wire  _GEN22458 = io_x[29] ? _GEN22457 : _GEN22455;
wire  _GEN22459 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22460 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22461 = io_x[27] ? _GEN22460 : _GEN22459;
wire  _GEN22462 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22463 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22464 = io_x[27] ? _GEN22463 : _GEN22462;
wire  _GEN22465 = io_x[29] ? _GEN22464 : _GEN22461;
wire  _GEN22466 = io_x[75] ? _GEN22465 : _GEN22458;
wire  _GEN22467 = io_x[38] ? _GEN22466 : _GEN22452;
wire  _GEN22468 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22469 = io_x[27] ? _GEN22468 : _GEN21739;
wire  _GEN22470 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22471 = io_x[27] ? _GEN22470 : _GEN21750;
wire  _GEN22472 = io_x[29] ? _GEN22471 : _GEN22469;
wire  _GEN22473 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22474 = io_x[27] ? _GEN21739 : _GEN22473;
wire  _GEN22475 = io_x[29] ? _GEN21743 : _GEN22474;
wire  _GEN22476 = io_x[75] ? _GEN22475 : _GEN22472;
wire  _GEN22477 = io_x[38] ? _GEN22476 : _GEN21833;
wire  _GEN22478 = io_x[34] ? _GEN22477 : _GEN22467;
wire  _GEN22479 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22480 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22481 = io_x[27] ? _GEN22480 : _GEN22479;
wire  _GEN22482 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22483 = io_x[27] ? _GEN21750 : _GEN22482;
wire  _GEN22484 = io_x[29] ? _GEN22483 : _GEN22481;
wire  _GEN22485 = io_x[75] ? _GEN21772 : _GEN22484;
wire  _GEN22486 = io_x[38] ? _GEN22485 : _GEN21871;
wire  _GEN22487 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22488 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22489 = io_x[27] ? _GEN22488 : _GEN22487;
wire  _GEN22490 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22491 = io_x[27] ? _GEN21739 : _GEN22490;
wire  _GEN22492 = io_x[29] ? _GEN22491 : _GEN22489;
wire  _GEN22493 = io_x[75] ? _GEN21758 : _GEN22492;
wire  _GEN22494 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22495 = io_x[27] ? _GEN21739 : _GEN22494;
wire  _GEN22496 = io_x[29] ? _GEN21744 : _GEN22495;
wire  _GEN22497 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22498 = io_x[27] ? _GEN21739 : _GEN22497;
wire  _GEN22499 = io_x[29] ? _GEN21743 : _GEN22498;
wire  _GEN22500 = io_x[75] ? _GEN22499 : _GEN22496;
wire  _GEN22501 = io_x[38] ? _GEN22500 : _GEN22493;
wire  _GEN22502 = io_x[34] ? _GEN22501 : _GEN22486;
wire  _GEN22503 = io_x[39] ? _GEN22502 : _GEN22478;
wire  _GEN22504 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22505 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22506 = io_x[27] ? _GEN22505 : _GEN22504;
wire  _GEN22507 = io_x[29] ? _GEN21744 : _GEN22506;
wire  _GEN22508 = io_x[75] ? _GEN22507 : _GEN21758;
wire  _GEN22509 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22510 = io_x[27] ? _GEN22509 : _GEN21739;
wire  _GEN22511 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22512 = io_x[27] ? _GEN21739 : _GEN22511;
wire  _GEN22513 = io_x[29] ? _GEN22512 : _GEN22510;
wire  _GEN22514 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22515 = io_x[27] ? _GEN21739 : _GEN22514;
wire  _GEN22516 = io_x[29] ? _GEN21744 : _GEN22515;
wire  _GEN22517 = io_x[75] ? _GEN22516 : _GEN22513;
wire  _GEN22518 = io_x[38] ? _GEN22517 : _GEN22508;
wire  _GEN22519 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22520 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22521 = io_x[27] ? _GEN22520 : _GEN22519;
wire  _GEN22522 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22523 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22524 = io_x[27] ? _GEN22523 : _GEN22522;
wire  _GEN22525 = io_x[29] ? _GEN22524 : _GEN22521;
wire  _GEN22526 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN22527 = io_x[29] ? _GEN22526 : _GEN21743;
wire  _GEN22528 = io_x[75] ? _GEN22527 : _GEN22525;
wire  _GEN22529 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22530 = io_x[27] ? _GEN21739 : _GEN22529;
wire  _GEN22531 = io_x[29] ? _GEN21743 : _GEN22530;
wire  _GEN22532 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22533 = io_x[27] ? _GEN21739 : _GEN22532;
wire  _GEN22534 = io_x[29] ? _GEN21743 : _GEN22533;
wire  _GEN22535 = io_x[75] ? _GEN22534 : _GEN22531;
wire  _GEN22536 = io_x[38] ? _GEN22535 : _GEN22528;
wire  _GEN22537 = io_x[34] ? _GEN22536 : _GEN22518;
wire  _GEN22538 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN22539 = io_x[29] ? _GEN21743 : _GEN22538;
wire  _GEN22540 = io_x[75] ? _GEN22539 : _GEN21758;
wire  _GEN22541 = io_x[38] ? _GEN21833 : _GEN22540;
wire  _GEN22542 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22543 = io_x[27] ? _GEN22542 : _GEN21739;
wire  _GEN22544 = io_x[29] ? _GEN22543 : _GEN21743;
wire  _GEN22545 = io_x[75] ? _GEN21772 : _GEN22544;
wire  _GEN22546 = io_x[38] ? _GEN22545 : _GEN21833;
wire  _GEN22547 = io_x[34] ? _GEN22546 : _GEN22541;
wire  _GEN22548 = io_x[39] ? _GEN22547 : _GEN22537;
wire  _GEN22549 = io_x[46] ? _GEN22548 : _GEN22503;
wire  _GEN22550 = io_x[18] ? _GEN22549 : _GEN22448;
wire  _GEN22551 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22552 = io_x[27] ? _GEN21739 : _GEN22551;
wire  _GEN22553 = io_x[29] ? _GEN21743 : _GEN22552;
wire  _GEN22554 = io_x[75] ? _GEN22553 : _GEN21758;
wire  _GEN22555 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22556 = io_x[27] ? _GEN21739 : _GEN22555;
wire  _GEN22557 = io_x[29] ? _GEN21744 : _GEN22556;
wire  _GEN22558 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22559 = io_x[27] ? _GEN21739 : _GEN22558;
wire  _GEN22560 = io_x[29] ? _GEN21743 : _GEN22559;
wire  _GEN22561 = io_x[75] ? _GEN22560 : _GEN22557;
wire  _GEN22562 = io_x[38] ? _GEN22561 : _GEN22554;
wire  _GEN22563 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22564 = io_x[27] ? _GEN21739 : _GEN22563;
wire  _GEN22565 = io_x[29] ? _GEN21743 : _GEN22564;
wire  _GEN22566 = io_x[75] ? _GEN21758 : _GEN22565;
wire  _GEN22567 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22568 = io_x[27] ? _GEN22567 : _GEN21739;
wire  _GEN22569 = io_x[29] ? _GEN22568 : _GEN21744;
wire  _GEN22570 = io_x[75] ? _GEN21772 : _GEN22569;
wire  _GEN22571 = io_x[38] ? _GEN22570 : _GEN22566;
wire  _GEN22572 = io_x[34] ? _GEN22571 : _GEN22562;
wire  _GEN22573 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN22574 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22575 = io_x[27] ? _GEN21739 : _GEN22574;
wire  _GEN22576 = io_x[29] ? _GEN21743 : _GEN22575;
wire  _GEN22577 = io_x[75] ? _GEN22576 : _GEN21772;
wire  _GEN22578 = io_x[38] ? _GEN21871 : _GEN22577;
wire  _GEN22579 = io_x[34] ? _GEN22578 : _GEN22573;
wire  _GEN22580 = io_x[39] ? _GEN22579 : _GEN22572;
wire  _GEN22581 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22582 = io_x[27] ? _GEN21739 : _GEN22581;
wire  _GEN22583 = io_x[29] ? _GEN21744 : _GEN22582;
wire  _GEN22584 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22585 = io_x[27] ? _GEN21739 : _GEN22584;
wire  _GEN22586 = io_x[29] ? _GEN21744 : _GEN22585;
wire  _GEN22587 = io_x[75] ? _GEN22586 : _GEN22583;
wire  _GEN22588 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22589 = io_x[27] ? _GEN21739 : _GEN22588;
wire  _GEN22590 = io_x[29] ? _GEN21744 : _GEN22589;
wire  _GEN22591 = io_x[75] ? _GEN22590 : _GEN21758;
wire  _GEN22592 = io_x[38] ? _GEN22591 : _GEN22587;
wire  _GEN22593 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22594 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22595 = io_x[27] ? _GEN21739 : _GEN22594;
wire  _GEN22596 = io_x[29] ? _GEN21743 : _GEN22595;
wire  _GEN22597 = io_x[75] ? _GEN21772 : _GEN22596;
wire  _GEN22598 = io_x[38] ? _GEN22597 : _GEN22593;
wire  _GEN22599 = io_x[34] ? _GEN22598 : _GEN22592;
wire  _GEN22600 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22601 = io_x[27] ? _GEN21739 : _GEN22600;
wire  _GEN22602 = io_x[29] ? _GEN22601 : _GEN21744;
wire  _GEN22603 = io_x[75] ? _GEN22602 : _GEN21772;
wire  _GEN22604 = io_x[38] ? _GEN22603 : _GEN21833;
wire  _GEN22605 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22606 = io_x[27] ? _GEN21739 : _GEN22605;
wire  _GEN22607 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22608 = io_x[27] ? _GEN21750 : _GEN22607;
wire  _GEN22609 = io_x[29] ? _GEN22608 : _GEN22606;
wire  _GEN22610 = io_x[75] ? _GEN22609 : _GEN21758;
wire  _GEN22611 = io_x[38] ? _GEN21833 : _GEN22610;
wire  _GEN22612 = io_x[34] ? _GEN22611 : _GEN22604;
wire  _GEN22613 = io_x[39] ? _GEN22612 : _GEN22599;
wire  _GEN22614 = io_x[46] ? _GEN22613 : _GEN22580;
wire  _GEN22615 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22616 = io_x[27] ? _GEN21739 : _GEN22615;
wire  _GEN22617 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN22618 = io_x[29] ? _GEN22617 : _GEN22616;
wire  _GEN22619 = io_x[75] ? _GEN21758 : _GEN22618;
wire  _GEN22620 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22621 = io_x[27] ? _GEN21739 : _GEN22620;
wire  _GEN22622 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22623 = io_x[27] ? _GEN22622 : _GEN21739;
wire  _GEN22624 = io_x[29] ? _GEN22623 : _GEN22621;
wire  _GEN22625 = io_x[75] ? _GEN22624 : _GEN21772;
wire  _GEN22626 = io_x[38] ? _GEN22625 : _GEN22619;
wire  _GEN22627 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN22628 = io_x[75] ? _GEN21772 : _GEN22627;
wire  _GEN22629 = io_x[38] ? _GEN22628 : _GEN21871;
wire  _GEN22630 = io_x[34] ? _GEN22629 : _GEN22626;
wire  _GEN22631 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22632 = io_x[27] ? _GEN21739 : _GEN22631;
wire  _GEN22633 = io_x[29] ? _GEN21743 : _GEN22632;
wire  _GEN22634 = io_x[75] ? _GEN21758 : _GEN22633;
wire  _GEN22635 = io_x[38] ? _GEN21833 : _GEN22634;
wire  _GEN22636 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22637 = io_x[27] ? _GEN21739 : _GEN22636;
wire  _GEN22638 = io_x[29] ? _GEN21743 : _GEN22637;
wire  _GEN22639 = io_x[75] ? _GEN22638 : _GEN21758;
wire  _GEN22640 = io_x[38] ? _GEN21833 : _GEN22639;
wire  _GEN22641 = io_x[34] ? _GEN22640 : _GEN22635;
wire  _GEN22642 = io_x[39] ? _GEN22641 : _GEN22630;
wire  _GEN22643 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22644 = io_x[27] ? _GEN21739 : _GEN22643;
wire  _GEN22645 = io_x[29] ? _GEN21743 : _GEN22644;
wire  _GEN22646 = io_x[75] ? _GEN22645 : _GEN21772;
wire  _GEN22647 = io_x[38] ? _GEN21833 : _GEN22646;
wire  _GEN22648 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22649 = io_x[27] ? _GEN21739 : _GEN22648;
wire  _GEN22650 = io_x[29] ? _GEN21743 : _GEN22649;
wire  _GEN22651 = io_x[75] ? _GEN21772 : _GEN22650;
wire  _GEN22652 = io_x[38] ? _GEN22651 : _GEN21833;
wire  _GEN22653 = io_x[34] ? _GEN22652 : _GEN22647;
wire  _GEN22654 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22655 = io_x[38] ? _GEN22654 : _GEN21833;
wire  _GEN22656 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22657 = io_x[38] ? _GEN21833 : _GEN22656;
wire  _GEN22658 = io_x[34] ? _GEN22657 : _GEN22655;
wire  _GEN22659 = io_x[39] ? _GEN22658 : _GEN22653;
wire  _GEN22660 = io_x[46] ? _GEN22659 : _GEN22642;
wire  _GEN22661 = io_x[18] ? _GEN22660 : _GEN22614;
wire  _GEN22662 = io_x[49] ? _GEN22661 : _GEN22550;
wire  _GEN22663 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22664 = io_x[27] ? _GEN21739 : _GEN22663;
wire  _GEN22665 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22666 = io_x[27] ? _GEN21739 : _GEN22665;
wire  _GEN22667 = io_x[29] ? _GEN22666 : _GEN22664;
wire  _GEN22668 = io_x[75] ? _GEN22667 : _GEN21758;
wire  _GEN22669 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22670 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22671 = io_x[27] ? _GEN22670 : _GEN22669;
wire  _GEN22672 = io_x[29] ? _GEN21743 : _GEN22671;
wire  _GEN22673 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22674 = io_x[27] ? _GEN21739 : _GEN22673;
wire  _GEN22675 = io_x[29] ? _GEN21743 : _GEN22674;
wire  _GEN22676 = io_x[75] ? _GEN22675 : _GEN22672;
wire  _GEN22677 = io_x[38] ? _GEN22676 : _GEN22668;
wire  _GEN22678 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22679 = io_x[27] ? _GEN21750 : _GEN22678;
wire  _GEN22680 = io_x[29] ? _GEN21744 : _GEN22679;
wire  _GEN22681 = io_x[75] ? _GEN21758 : _GEN22680;
wire  _GEN22682 = io_x[38] ? _GEN22681 : _GEN21871;
wire  _GEN22683 = io_x[34] ? _GEN22682 : _GEN22677;
wire  _GEN22684 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN22685 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22686 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22687 = io_x[27] ? _GEN22686 : _GEN22685;
wire  _GEN22688 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22689 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22690 = io_x[27] ? _GEN22689 : _GEN22688;
wire  _GEN22691 = io_x[29] ? _GEN22690 : _GEN22687;
wire  _GEN22692 = io_x[75] ? _GEN21772 : _GEN22691;
wire  _GEN22693 = io_x[38] ? _GEN22692 : _GEN22684;
wire  _GEN22694 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN22695 = io_x[29] ? _GEN22694 : _GEN21743;
wire  _GEN22696 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN22697 = io_x[75] ? _GEN22696 : _GEN22695;
wire  _GEN22698 = io_x[38] ? _GEN21871 : _GEN22697;
wire  _GEN22699 = io_x[34] ? _GEN22698 : _GEN22693;
wire  _GEN22700 = io_x[39] ? _GEN22699 : _GEN22683;
wire  _GEN22701 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22702 = io_x[27] ? _GEN21739 : _GEN22701;
wire  _GEN22703 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22704 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22705 = io_x[27] ? _GEN22704 : _GEN22703;
wire  _GEN22706 = io_x[29] ? _GEN22705 : _GEN22702;
wire  _GEN22707 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22708 = io_x[27] ? _GEN22707 : _GEN21739;
wire  _GEN22709 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN22710 = io_x[29] ? _GEN22709 : _GEN22708;
wire  _GEN22711 = io_x[75] ? _GEN22710 : _GEN22706;
wire  _GEN22712 = io_x[38] ? _GEN22711 : _GEN21833;
wire  _GEN22713 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22714 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22715 = io_x[27] ? _GEN22714 : _GEN22713;
wire  _GEN22716 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22717 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22718 = io_x[27] ? _GEN22717 : _GEN22716;
wire  _GEN22719 = io_x[29] ? _GEN22718 : _GEN22715;
wire  _GEN22720 = io_x[75] ? _GEN21772 : _GEN22719;
wire  _GEN22721 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22722 = io_x[38] ? _GEN22721 : _GEN22720;
wire  _GEN22723 = io_x[34] ? _GEN22722 : _GEN22712;
wire  _GEN22724 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22725 = io_x[27] ? _GEN21739 : _GEN22724;
wire  _GEN22726 = io_x[29] ? _GEN22725 : _GEN21743;
wire  _GEN22727 = io_x[75] ? _GEN21758 : _GEN22726;
wire  _GEN22728 = io_x[38] ? _GEN22727 : _GEN21871;
wire  _GEN22729 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN22730 = io_x[29] ? _GEN22729 : _GEN21744;
wire  _GEN22731 = io_x[75] ? _GEN22730 : _GEN21758;
wire  _GEN22732 = io_x[38] ? _GEN22731 : _GEN21833;
wire  _GEN22733 = io_x[34] ? _GEN22732 : _GEN22728;
wire  _GEN22734 = io_x[39] ? _GEN22733 : _GEN22723;
wire  _GEN22735 = io_x[46] ? _GEN22734 : _GEN22700;
wire  _GEN22736 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22737 = io_x[27] ? _GEN22736 : _GEN21739;
wire  _GEN22738 = io_x[29] ? _GEN22737 : _GEN21743;
wire  _GEN22739 = io_x[75] ? _GEN21772 : _GEN22738;
wire  _GEN22740 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22741 = io_x[27] ? _GEN21750 : _GEN22740;
wire  _GEN22742 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22743 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22744 = io_x[27] ? _GEN22743 : _GEN22742;
wire  _GEN22745 = io_x[29] ? _GEN22744 : _GEN22741;
wire  _GEN22746 = io_x[75] ? _GEN21758 : _GEN22745;
wire  _GEN22747 = io_x[38] ? _GEN22746 : _GEN22739;
wire  _GEN22748 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22749 = io_x[27] ? _GEN22748 : _GEN21750;
wire  _GEN22750 = io_x[29] ? _GEN22749 : _GEN21743;
wire  _GEN22751 = io_x[75] ? _GEN21758 : _GEN22750;
wire  _GEN22752 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22753 = io_x[27] ? _GEN22752 : _GEN21739;
wire  _GEN22754 = io_x[29] ? _GEN22753 : _GEN21743;
wire  _GEN22755 = io_x[75] ? _GEN21758 : _GEN22754;
wire  _GEN22756 = io_x[38] ? _GEN22755 : _GEN22751;
wire  _GEN22757 = io_x[34] ? _GEN22756 : _GEN22747;
wire  _GEN22758 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN22759 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22760 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22761 = io_x[27] ? _GEN22760 : _GEN22759;
wire  _GEN22762 = io_x[29] ? _GEN22761 : _GEN22758;
wire  _GEN22763 = io_x[75] ? _GEN21758 : _GEN22762;
wire  _GEN22764 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22765 = io_x[27] ? _GEN21739 : _GEN22764;
wire  _GEN22766 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22767 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22768 = io_x[27] ? _GEN22767 : _GEN22766;
wire  _GEN22769 = io_x[29] ? _GEN22768 : _GEN22765;
wire  _GEN22770 = io_x[75] ? _GEN21772 : _GEN22769;
wire  _GEN22771 = io_x[38] ? _GEN22770 : _GEN22763;
wire  _GEN22772 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22773 = io_x[27] ? _GEN22772 : _GEN21739;
wire  _GEN22774 = io_x[29] ? _GEN22773 : _GEN21743;
wire  _GEN22775 = io_x[75] ? _GEN21772 : _GEN22774;
wire  _GEN22776 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN22777 = io_x[75] ? _GEN21758 : _GEN22776;
wire  _GEN22778 = io_x[38] ? _GEN22777 : _GEN22775;
wire  _GEN22779 = io_x[34] ? _GEN22778 : _GEN22771;
wire  _GEN22780 = io_x[39] ? _GEN22779 : _GEN22757;
wire  _GEN22781 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22782 = io_x[27] ? _GEN21739 : _GEN22781;
wire  _GEN22783 = io_x[29] ? _GEN22782 : _GEN21743;
wire  _GEN22784 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN22785 = io_x[29] ? _GEN21744 : _GEN22784;
wire  _GEN22786 = io_x[75] ? _GEN22785 : _GEN22783;
wire  _GEN22787 = io_x[38] ? _GEN22786 : _GEN21833;
wire  _GEN22788 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22789 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22790 = io_x[27] ? _GEN22789 : _GEN22788;
wire  _GEN22791 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22792 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22793 = io_x[27] ? _GEN22792 : _GEN22791;
wire  _GEN22794 = io_x[29] ? _GEN22793 : _GEN22790;
wire  _GEN22795 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22796 = io_x[27] ? _GEN21739 : _GEN22795;
wire  _GEN22797 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22798 = io_x[27] ? _GEN22797 : _GEN21739;
wire  _GEN22799 = io_x[29] ? _GEN22798 : _GEN22796;
wire  _GEN22800 = io_x[75] ? _GEN22799 : _GEN22794;
wire  _GEN22801 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22802 = io_x[27] ? _GEN22801 : _GEN21739;
wire  _GEN22803 = io_x[29] ? _GEN22802 : _GEN21744;
wire  _GEN22804 = io_x[75] ? _GEN22803 : _GEN21758;
wire  _GEN22805 = io_x[38] ? _GEN22804 : _GEN22800;
wire  _GEN22806 = io_x[34] ? _GEN22805 : _GEN22787;
wire  _GEN22807 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN22808 = io_x[29] ? _GEN22807 : _GEN21743;
wire  _GEN22809 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22810 = io_x[27] ? _GEN21739 : _GEN22809;
wire  _GEN22811 = io_x[29] ? _GEN22810 : _GEN21744;
wire  _GEN22812 = io_x[75] ? _GEN22811 : _GEN22808;
wire  _GEN22813 = io_x[38] ? _GEN22812 : _GEN21833;
wire  _GEN22814 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN22815 = io_x[29] ? _GEN21743 : _GEN22814;
wire  _GEN22816 = io_x[75] ? _GEN21772 : _GEN22815;
wire  _GEN22817 = io_x[38] ? _GEN22816 : _GEN21833;
wire  _GEN22818 = io_x[34] ? _GEN22817 : _GEN22813;
wire  _GEN22819 = io_x[39] ? _GEN22818 : _GEN22806;
wire  _GEN22820 = io_x[46] ? _GEN22819 : _GEN22780;
wire  _GEN22821 = io_x[18] ? _GEN22820 : _GEN22735;
wire  _GEN22822 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22823 = io_x[27] ? _GEN22822 : _GEN21739;
wire  _GEN22824 = io_x[29] ? _GEN22823 : _GEN21744;
wire  _GEN22825 = io_x[75] ? _GEN21758 : _GEN22824;
wire  _GEN22826 = io_x[38] ? _GEN22825 : _GEN21833;
wire  _GEN22827 = io_x[34] ? _GEN22826 : _GEN21766;
wire  _GEN22828 = io_x[39] ? _GEN21910 : _GEN22827;
wire  _GEN22829 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22830 = io_x[27] ? _GEN22829 : _GEN21739;
wire  _GEN22831 = io_x[29] ? _GEN22830 : _GEN21743;
wire  _GEN22832 = io_x[75] ? _GEN21772 : _GEN22831;
wire  _GEN22833 = io_x[38] ? _GEN22832 : _GEN21833;
wire  _GEN22834 = io_x[34] ? _GEN22833 : _GEN21766;
wire  _GEN22835 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22836 = io_x[27] ? _GEN22835 : _GEN21750;
wire  _GEN22837 = io_x[29] ? _GEN22836 : _GEN21744;
wire  _GEN22838 = io_x[75] ? _GEN22837 : _GEN21758;
wire  _GEN22839 = io_x[38] ? _GEN22838 : _GEN21833;
wire  _GEN22840 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22841 = io_x[27] ? _GEN22840 : _GEN21750;
wire  _GEN22842 = io_x[29] ? _GEN22841 : _GEN21744;
wire  _GEN22843 = io_x[75] ? _GEN22842 : _GEN21758;
wire  _GEN22844 = io_x[38] ? _GEN21833 : _GEN22843;
wire  _GEN22845 = io_x[34] ? _GEN22844 : _GEN22839;
wire  _GEN22846 = io_x[39] ? _GEN22845 : _GEN22834;
wire  _GEN22847 = io_x[46] ? _GEN22846 : _GEN22828;
wire  _GEN22848 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN22849 = io_x[75] ? _GEN21758 : _GEN22848;
wire  _GEN22850 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22851 = io_x[27] ? _GEN21750 : _GEN22850;
wire  _GEN22852 = io_x[29] ? _GEN21743 : _GEN22851;
wire  _GEN22853 = io_x[75] ? _GEN21758 : _GEN22852;
wire  _GEN22854 = io_x[38] ? _GEN22853 : _GEN22849;
wire  _GEN22855 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN22856 = io_x[29] ? _GEN22855 : _GEN21743;
wire  _GEN22857 = io_x[75] ? _GEN22856 : _GEN21758;
wire  _GEN22858 = io_x[38] ? _GEN21871 : _GEN22857;
wire  _GEN22859 = io_x[34] ? _GEN22858 : _GEN22854;
wire  _GEN22860 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN22861 = io_x[38] ? _GEN21833 : _GEN22860;
wire  _GEN22862 = io_x[34] ? _GEN21927 : _GEN22861;
wire  _GEN22863 = io_x[39] ? _GEN22862 : _GEN22859;
wire  _GEN22864 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22865 = io_x[27] ? _GEN22864 : _GEN21739;
wire  _GEN22866 = io_x[29] ? _GEN21743 : _GEN22865;
wire  _GEN22867 = io_x[75] ? _GEN21758 : _GEN22866;
wire  _GEN22868 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22869 = io_x[27] ? _GEN21739 : _GEN22868;
wire  _GEN22870 = io_x[29] ? _GEN21743 : _GEN22869;
wire  _GEN22871 = io_x[75] ? _GEN21772 : _GEN22870;
wire  _GEN22872 = io_x[38] ? _GEN22871 : _GEN22867;
wire  _GEN22873 = io_x[34] ? _GEN22872 : _GEN21766;
wire  _GEN22874 = io_x[39] ? _GEN21910 : _GEN22873;
wire  _GEN22875 = io_x[46] ? _GEN22874 : _GEN22863;
wire  _GEN22876 = io_x[18] ? _GEN22875 : _GEN22847;
wire  _GEN22877 = io_x[49] ? _GEN22876 : _GEN22821;
wire  _GEN22878 = io_x[24] ? _GEN22877 : _GEN22662;
wire  _GEN22879 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN22880 = io_x[29] ? _GEN21743 : _GEN22879;
wire  _GEN22881 = io_x[75] ? _GEN21758 : _GEN22880;
wire  _GEN22882 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22883 = io_x[27] ? _GEN21739 : _GEN22882;
wire  _GEN22884 = io_x[29] ? _GEN21743 : _GEN22883;
wire  _GEN22885 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22886 = io_x[27] ? _GEN21739 : _GEN22885;
wire  _GEN22887 = io_x[29] ? _GEN21743 : _GEN22886;
wire  _GEN22888 = io_x[75] ? _GEN22887 : _GEN22884;
wire  _GEN22889 = io_x[38] ? _GEN22888 : _GEN22881;
wire  _GEN22890 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN22891 = io_x[34] ? _GEN22890 : _GEN22889;
wire  _GEN22892 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22893 = io_x[27] ? _GEN21739 : _GEN22892;
wire  _GEN22894 = io_x[29] ? _GEN21744 : _GEN22893;
wire  _GEN22895 = io_x[75] ? _GEN21758 : _GEN22894;
wire  _GEN22896 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22897 = io_x[27] ? _GEN21739 : _GEN22896;
wire  _GEN22898 = io_x[29] ? _GEN21744 : _GEN22897;
wire  _GEN22899 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN22900 = io_x[75] ? _GEN22899 : _GEN22898;
wire  _GEN22901 = io_x[38] ? _GEN22900 : _GEN22895;
wire  _GEN22902 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22903 = io_x[27] ? _GEN21739 : _GEN22902;
wire  _GEN22904 = io_x[29] ? _GEN21743 : _GEN22903;
wire  _GEN22905 = io_x[75] ? _GEN21758 : _GEN22904;
wire  _GEN22906 = io_x[38] ? _GEN22905 : _GEN21871;
wire  _GEN22907 = io_x[34] ? _GEN22906 : _GEN22901;
wire  _GEN22908 = io_x[39] ? _GEN22907 : _GEN22891;
wire  _GEN22909 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22910 = io_x[27] ? _GEN21739 : _GEN22909;
wire  _GEN22911 = io_x[29] ? _GEN21744 : _GEN22910;
wire  _GEN22912 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22913 = io_x[27] ? _GEN21739 : _GEN22912;
wire  _GEN22914 = io_x[29] ? _GEN21743 : _GEN22913;
wire  _GEN22915 = io_x[75] ? _GEN22914 : _GEN22911;
wire  _GEN22916 = io_x[38] ? _GEN22915 : _GEN21833;
wire  _GEN22917 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN22918 = io_x[38] ? _GEN22917 : _GEN21833;
wire  _GEN22919 = io_x[34] ? _GEN22918 : _GEN22916;
wire  _GEN22920 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22921 = io_x[27] ? _GEN21750 : _GEN22920;
wire  _GEN22922 = io_x[29] ? _GEN21744 : _GEN22921;
wire  _GEN22923 = io_x[75] ? _GEN21772 : _GEN22922;
wire  _GEN22924 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22925 = io_x[27] ? _GEN21750 : _GEN22924;
wire  _GEN22926 = io_x[29] ? _GEN21744 : _GEN22925;
wire  _GEN22927 = io_x[75] ? _GEN21758 : _GEN22926;
wire  _GEN22928 = io_x[38] ? _GEN22927 : _GEN22923;
wire  _GEN22929 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22930 = io_x[27] ? _GEN21739 : _GEN22929;
wire  _GEN22931 = io_x[29] ? _GEN21743 : _GEN22930;
wire  _GEN22932 = io_x[75] ? _GEN22931 : _GEN21758;
wire  _GEN22933 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22934 = io_x[27] ? _GEN21739 : _GEN22933;
wire  _GEN22935 = io_x[29] ? _GEN21744 : _GEN22934;
wire  _GEN22936 = io_x[75] ? _GEN22935 : _GEN21772;
wire  _GEN22937 = io_x[38] ? _GEN22936 : _GEN22932;
wire  _GEN22938 = io_x[34] ? _GEN22937 : _GEN22928;
wire  _GEN22939 = io_x[39] ? _GEN22938 : _GEN22919;
wire  _GEN22940 = io_x[46] ? _GEN22939 : _GEN22908;
wire  _GEN22941 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN22942 = io_x[29] ? _GEN22941 : _GEN21744;
wire  _GEN22943 = io_x[75] ? _GEN21758 : _GEN22942;
wire  _GEN22944 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22945 = io_x[27] ? _GEN21739 : _GEN22944;
wire  _GEN22946 = io_x[29] ? _GEN21744 : _GEN22945;
wire  _GEN22947 = io_x[75] ? _GEN21758 : _GEN22946;
wire  _GEN22948 = io_x[38] ? _GEN22947 : _GEN22943;
wire  _GEN22949 = io_x[34] ? _GEN21766 : _GEN22948;
wire  _GEN22950 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22951 = io_x[27] ? _GEN21739 : _GEN22950;
wire  _GEN22952 = io_x[29] ? _GEN21743 : _GEN22951;
wire  _GEN22953 = io_x[75] ? _GEN21758 : _GEN22952;
wire  _GEN22954 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22955 = io_x[27] ? _GEN21739 : _GEN22954;
wire  _GEN22956 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22957 = io_x[27] ? _GEN21739 : _GEN22956;
wire  _GEN22958 = io_x[29] ? _GEN22957 : _GEN22955;
wire  _GEN22959 = io_x[75] ? _GEN21758 : _GEN22958;
wire  _GEN22960 = io_x[38] ? _GEN22959 : _GEN22953;
wire  _GEN22961 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN22962 = io_x[38] ? _GEN21833 : _GEN22961;
wire  _GEN22963 = io_x[34] ? _GEN22962 : _GEN22960;
wire  _GEN22964 = io_x[39] ? _GEN22963 : _GEN22949;
wire  _GEN22965 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22966 = io_x[27] ? _GEN21739 : _GEN22965;
wire  _GEN22967 = io_x[29] ? _GEN21743 : _GEN22966;
wire  _GEN22968 = io_x[75] ? _GEN21772 : _GEN22967;
wire  _GEN22969 = io_x[38] ? _GEN22968 : _GEN21871;
wire  _GEN22970 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22971 = io_x[27] ? _GEN21739 : _GEN22970;
wire  _GEN22972 = io_x[29] ? _GEN21744 : _GEN22971;
wire  _GEN22973 = io_x[75] ? _GEN21758 : _GEN22972;
wire  _GEN22974 = io_x[38] ? _GEN21871 : _GEN22973;
wire  _GEN22975 = io_x[34] ? _GEN22974 : _GEN22969;
wire  _GEN22976 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22977 = io_x[27] ? _GEN21739 : _GEN22976;
wire  _GEN22978 = io_x[29] ? _GEN21743 : _GEN22977;
wire  _GEN22979 = io_x[75] ? _GEN21772 : _GEN22978;
wire  _GEN22980 = io_x[38] ? _GEN21871 : _GEN22979;
wire  _GEN22981 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22982 = io_x[27] ? _GEN21739 : _GEN22981;
wire  _GEN22983 = io_x[29] ? _GEN21744 : _GEN22982;
wire  _GEN22984 = io_x[75] ? _GEN21758 : _GEN22983;
wire  _GEN22985 = io_x[38] ? _GEN21871 : _GEN22984;
wire  _GEN22986 = io_x[34] ? _GEN22985 : _GEN22980;
wire  _GEN22987 = io_x[39] ? _GEN22986 : _GEN22975;
wire  _GEN22988 = io_x[46] ? _GEN22987 : _GEN22964;
wire  _GEN22989 = io_x[18] ? _GEN22988 : _GEN22940;
wire  _GEN22990 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22991 = io_x[27] ? _GEN21739 : _GEN22990;
wire  _GEN22992 = io_x[29] ? _GEN21743 : _GEN22991;
wire  _GEN22993 = io_x[75] ? _GEN22992 : _GEN21758;
wire  _GEN22994 = io_x[38] ? _GEN21833 : _GEN22993;
wire  _GEN22995 = io_x[34] ? _GEN21927 : _GEN22994;
wire  _GEN22996 = io_x[39] ? _GEN21910 : _GEN22995;
wire  _GEN22997 = io_x[46] ? _GEN22145 : _GEN22996;
wire  _GEN22998 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN22999 = io_x[27] ? _GEN21739 : _GEN22998;
wire  _GEN23000 = io_x[29] ? _GEN21743 : _GEN22999;
wire  _GEN23001 = io_x[75] ? _GEN23000 : _GEN21758;
wire  _GEN23002 = io_x[38] ? _GEN23001 : _GEN21833;
wire  _GEN23003 = io_x[34] ? _GEN21927 : _GEN23002;
wire  _GEN23004 = io_x[39] ? _GEN21910 : _GEN23003;
wire  _GEN23005 = io_x[46] ? _GEN22145 : _GEN23004;
wire  _GEN23006 = io_x[18] ? _GEN23005 : _GEN22997;
wire  _GEN23007 = io_x[49] ? _GEN23006 : _GEN22989;
wire  _GEN23008 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23009 = io_x[27] ? _GEN23008 : _GEN21739;
wire  _GEN23010 = io_x[29] ? _GEN21743 : _GEN23009;
wire  _GEN23011 = io_x[75] ? _GEN23010 : _GEN21758;
wire  _GEN23012 = io_x[38] ? _GEN21871 : _GEN23011;
wire  _GEN23013 = io_x[34] ? _GEN21927 : _GEN23012;
wire  _GEN23014 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23015 = io_x[27] ? _GEN23014 : _GEN21739;
wire  _GEN23016 = io_x[29] ? _GEN23015 : _GEN21744;
wire  _GEN23017 = io_x[75] ? _GEN21758 : _GEN23016;
wire  _GEN23018 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23019 = io_x[27] ? _GEN23018 : _GEN21739;
wire  _GEN23020 = io_x[29] ? _GEN21744 : _GEN23019;
wire  _GEN23021 = io_x[75] ? _GEN21758 : _GEN23020;
wire  _GEN23022 = io_x[38] ? _GEN23021 : _GEN23017;
wire  _GEN23023 = io_x[34] ? _GEN21927 : _GEN23022;
wire  _GEN23024 = io_x[39] ? _GEN23023 : _GEN23013;
wire  _GEN23025 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN23026 = io_x[38] ? _GEN21871 : _GEN23025;
wire  _GEN23027 = io_x[34] ? _GEN23026 : _GEN21766;
wire  _GEN23028 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN23029 = io_x[75] ? _GEN21758 : _GEN23028;
wire  _GEN23030 = io_x[38] ? _GEN21871 : _GEN23029;
wire  _GEN23031 = io_x[34] ? _GEN23030 : _GEN21766;
wire  _GEN23032 = io_x[39] ? _GEN23031 : _GEN23027;
wire  _GEN23033 = io_x[46] ? _GEN23032 : _GEN23024;
wire  _GEN23034 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN23035 = io_x[38] ? _GEN21833 : _GEN23034;
wire  _GEN23036 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23037 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23038 = io_x[27] ? _GEN23037 : _GEN23036;
wire  _GEN23039 = io_x[29] ? _GEN23038 : _GEN21743;
wire  _GEN23040 = io_x[75] ? _GEN23039 : _GEN21772;
wire  _GEN23041 = io_x[38] ? _GEN21833 : _GEN23040;
wire  _GEN23042 = io_x[34] ? _GEN23041 : _GEN23035;
wire  _GEN23043 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23044 = io_x[27] ? _GEN23043 : _GEN21739;
wire  _GEN23045 = io_x[29] ? _GEN23044 : _GEN21743;
wire  _GEN23046 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN23047 = io_x[29] ? _GEN23046 : _GEN21744;
wire  _GEN23048 = io_x[75] ? _GEN23047 : _GEN23045;
wire  _GEN23049 = io_x[38] ? _GEN23048 : _GEN21833;
wire  _GEN23050 = io_x[34] ? _GEN21927 : _GEN23049;
wire  _GEN23051 = io_x[39] ? _GEN23050 : _GEN23042;
wire  _GEN23052 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN23053 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23054 = io_x[27] ? _GEN23053 : _GEN21739;
wire  _GEN23055 = io_x[29] ? _GEN23054 : _GEN21743;
wire  _GEN23056 = io_x[75] ? _GEN23055 : _GEN23052;
wire  _GEN23057 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN23058 = io_x[29] ? _GEN23057 : _GEN21744;
wire  _GEN23059 = io_x[75] ? _GEN23058 : _GEN21772;
wire  _GEN23060 = io_x[38] ? _GEN23059 : _GEN23056;
wire  _GEN23061 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN23062 = io_x[29] ? _GEN23061 : _GEN21744;
wire  _GEN23063 = io_x[75] ? _GEN21758 : _GEN23062;
wire  _GEN23064 = io_x[38] ? _GEN21871 : _GEN23063;
wire  _GEN23065 = io_x[34] ? _GEN23064 : _GEN23060;
wire  _GEN23066 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN23067 = io_x[38] ? _GEN23066 : _GEN21871;
wire  _GEN23068 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23069 = io_x[27] ? _GEN21739 : _GEN23068;
wire  _GEN23070 = io_x[29] ? _GEN21744 : _GEN23069;
wire  _GEN23071 = io_x[75] ? _GEN21758 : _GEN23070;
wire  _GEN23072 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN23073 = io_x[29] ? _GEN23072 : _GEN21743;
wire  _GEN23074 = io_x[75] ? _GEN23073 : _GEN21772;
wire  _GEN23075 = io_x[38] ? _GEN23074 : _GEN23071;
wire  _GEN23076 = io_x[34] ? _GEN23075 : _GEN23067;
wire  _GEN23077 = io_x[39] ? _GEN23076 : _GEN23065;
wire  _GEN23078 = io_x[46] ? _GEN23077 : _GEN23051;
wire  _GEN23079 = io_x[18] ? _GEN23078 : _GEN23033;
wire  _GEN23080 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN23081 = io_x[34] ? _GEN23080 : _GEN21766;
wire  _GEN23082 = io_x[39] ? _GEN22327 : _GEN23081;
wire  _GEN23083 = io_x[46] ? _GEN22145 : _GEN23082;
wire  _GEN23084 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23085 = io_x[27] ? _GEN23084 : _GEN21739;
wire  _GEN23086 = io_x[29] ? _GEN23085 : _GEN21743;
wire  _GEN23087 = io_x[75] ? _GEN23086 : _GEN21758;
wire  _GEN23088 = io_x[38] ? _GEN23087 : _GEN21833;
wire  _GEN23089 = io_x[34] ? _GEN21766 : _GEN23088;
wire  _GEN23090 = io_x[39] ? _GEN22327 : _GEN23089;
wire  _GEN23091 = io_x[46] ? _GEN22145 : _GEN23090;
wire  _GEN23092 = io_x[18] ? _GEN23091 : _GEN23083;
wire  _GEN23093 = io_x[49] ? _GEN23092 : _GEN23079;
wire  _GEN23094 = io_x[24] ? _GEN23093 : _GEN23007;
wire  _GEN23095 = io_x[80] ? _GEN23094 : _GEN22878;
wire  _GEN23096 = io_x[16] ? _GEN23095 : _GEN22342;
wire  _GEN23097 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN23098 = io_x[29] ? _GEN23097 : _GEN21744;
wire  _GEN23099 = io_x[75] ? _GEN21758 : _GEN23098;
wire  _GEN23100 = io_x[38] ? _GEN23099 : _GEN21833;
wire  _GEN23101 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN23102 = io_x[38] ? _GEN23101 : _GEN21833;
wire  _GEN23103 = io_x[34] ? _GEN23102 : _GEN23100;
wire  _GEN23104 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN23105 = io_x[75] ? _GEN21772 : _GEN23104;
wire  _GEN23106 = io_x[38] ? _GEN21871 : _GEN23105;
wire  _GEN23107 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23108 = io_x[27] ? _GEN21739 : _GEN23107;
wire  _GEN23109 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23110 = io_x[27] ? _GEN23109 : _GEN21739;
wire  _GEN23111 = io_x[29] ? _GEN23110 : _GEN23108;
wire  _GEN23112 = io_x[75] ? _GEN21772 : _GEN23111;
wire  _GEN23113 = io_x[38] ? _GEN21833 : _GEN23112;
wire  _GEN23114 = io_x[34] ? _GEN23113 : _GEN23106;
wire  _GEN23115 = io_x[39] ? _GEN23114 : _GEN23103;
wire  _GEN23116 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23117 = io_x[27] ? _GEN21739 : _GEN23116;
wire  _GEN23118 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23119 = io_x[27] ? _GEN23118 : _GEN21739;
wire  _GEN23120 = io_x[29] ? _GEN23119 : _GEN23117;
wire  _GEN23121 = io_x[75] ? _GEN21772 : _GEN23120;
wire  _GEN23122 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23123 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23124 = io_x[27] ? _GEN23123 : _GEN23122;
wire  _GEN23125 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23126 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23127 = io_x[27] ? _GEN23126 : _GEN23125;
wire  _GEN23128 = io_x[29] ? _GEN23127 : _GEN23124;
wire  _GEN23129 = io_x[75] ? _GEN21772 : _GEN23128;
wire  _GEN23130 = io_x[38] ? _GEN23129 : _GEN23121;
wire  _GEN23131 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23132 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23133 = io_x[27] ? _GEN23132 : _GEN23131;
wire  _GEN23134 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23135 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23136 = io_x[27] ? _GEN23135 : _GEN23134;
wire  _GEN23137 = io_x[29] ? _GEN23136 : _GEN23133;
wire  _GEN23138 = io_x[75] ? _GEN21758 : _GEN23137;
wire  _GEN23139 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23140 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23141 = io_x[27] ? _GEN23140 : _GEN23139;
wire  _GEN23142 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23143 = io_x[27] ? _GEN21739 : _GEN23142;
wire  _GEN23144 = io_x[29] ? _GEN23143 : _GEN23141;
wire  _GEN23145 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN23146 = io_x[75] ? _GEN23145 : _GEN23144;
wire  _GEN23147 = io_x[38] ? _GEN23146 : _GEN23138;
wire  _GEN23148 = io_x[34] ? _GEN23147 : _GEN23130;
wire  _GEN23149 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23150 = io_x[27] ? _GEN23149 : _GEN21739;
wire  _GEN23151 = io_x[29] ? _GEN23150 : _GEN21743;
wire  _GEN23152 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN23153 = io_x[75] ? _GEN23152 : _GEN23151;
wire  _GEN23154 = io_x[38] ? _GEN23153 : _GEN21871;
wire  _GEN23155 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23156 = io_x[38] ? _GEN23155 : _GEN21833;
wire  _GEN23157 = io_x[34] ? _GEN23156 : _GEN23154;
wire  _GEN23158 = io_x[39] ? _GEN23157 : _GEN23148;
wire  _GEN23159 = io_x[46] ? _GEN23158 : _GEN23115;
wire  _GEN23160 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23161 = io_x[38] ? _GEN23160 : _GEN21833;
wire  _GEN23162 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN23163 = io_x[34] ? _GEN23162 : _GEN23161;
wire  _GEN23164 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23165 = io_x[27] ? _GEN23164 : _GEN21739;
wire  _GEN23166 = io_x[29] ? _GEN23165 : _GEN21743;
wire  _GEN23167 = io_x[75] ? _GEN21772 : _GEN23166;
wire  _GEN23168 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23169 = io_x[27] ? _GEN23168 : _GEN21739;
wire  _GEN23170 = io_x[29] ? _GEN23169 : _GEN21744;
wire  _GEN23171 = io_x[75] ? _GEN21758 : _GEN23170;
wire  _GEN23172 = io_x[38] ? _GEN23171 : _GEN23167;
wire  _GEN23173 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN23174 = io_x[34] ? _GEN23173 : _GEN23172;
wire  _GEN23175 = io_x[39] ? _GEN23174 : _GEN23163;
wire  _GEN23176 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23177 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23178 = io_x[27] ? _GEN23177 : _GEN23176;
wire  _GEN23179 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23180 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23181 = io_x[27] ? _GEN23180 : _GEN23179;
wire  _GEN23182 = io_x[29] ? _GEN23181 : _GEN23178;
wire  _GEN23183 = io_x[75] ? _GEN21758 : _GEN23182;
wire  _GEN23184 = io_x[38] ? _GEN23183 : _GEN21833;
wire  _GEN23185 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23186 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23187 = io_x[27] ? _GEN23186 : _GEN23185;
wire  _GEN23188 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23189 = io_x[27] ? _GEN21739 : _GEN23188;
wire  _GEN23190 = io_x[29] ? _GEN23189 : _GEN23187;
wire  _GEN23191 = io_x[75] ? _GEN21758 : _GEN23190;
wire  _GEN23192 = io_x[38] ? _GEN21833 : _GEN23191;
wire  _GEN23193 = io_x[34] ? _GEN23192 : _GEN23184;
wire  _GEN23194 = io_x[39] ? _GEN21910 : _GEN23193;
wire  _GEN23195 = io_x[46] ? _GEN23194 : _GEN23175;
wire  _GEN23196 = io_x[18] ? _GEN23195 : _GEN23159;
wire  _GEN23197 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN23198 = io_x[29] ? _GEN21743 : _GEN23197;
wire  _GEN23199 = io_x[75] ? _GEN21758 : _GEN23198;
wire  _GEN23200 = io_x[38] ? _GEN23199 : _GEN21833;
wire  _GEN23201 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23202 = io_x[38] ? _GEN21833 : _GEN23201;
wire  _GEN23203 = io_x[34] ? _GEN23202 : _GEN23200;
wire  _GEN23204 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN23205 = io_x[38] ? _GEN23204 : _GEN21871;
wire  _GEN23206 = io_x[34] ? _GEN21766 : _GEN23205;
wire  _GEN23207 = io_x[39] ? _GEN23206 : _GEN23203;
wire  _GEN23208 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23209 = io_x[27] ? _GEN21739 : _GEN23208;
wire  _GEN23210 = io_x[29] ? _GEN23209 : _GEN21743;
wire  _GEN23211 = io_x[75] ? _GEN21772 : _GEN23210;
wire  _GEN23212 = io_x[38] ? _GEN21871 : _GEN23211;
wire  _GEN23213 = io_x[34] ? _GEN21927 : _GEN23212;
wire  _GEN23214 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23215 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23216 = io_x[27] ? _GEN23215 : _GEN23214;
wire  _GEN23217 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23218 = io_x[27] ? _GEN21739 : _GEN23217;
wire  _GEN23219 = io_x[29] ? _GEN23218 : _GEN23216;
wire  _GEN23220 = io_x[75] ? _GEN23219 : _GEN21758;
wire  _GEN23221 = io_x[38] ? _GEN21833 : _GEN23220;
wire  _GEN23222 = io_x[34] ? _GEN23221 : _GEN21927;
wire  _GEN23223 = io_x[39] ? _GEN23222 : _GEN23213;
wire  _GEN23224 = io_x[46] ? _GEN23223 : _GEN23207;
wire  _GEN23225 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN23226 = io_x[34] ? _GEN23225 : _GEN21927;
wire  _GEN23227 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN23228 = io_x[38] ? _GEN23227 : _GEN21833;
wire  _GEN23229 = io_x[34] ? _GEN21766 : _GEN23228;
wire  _GEN23230 = io_x[39] ? _GEN23229 : _GEN23226;
wire  _GEN23231 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN23232 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23233 = io_x[38] ? _GEN23232 : _GEN21833;
wire  _GEN23234 = io_x[34] ? _GEN23233 : _GEN23231;
wire  _GEN23235 = io_x[39] ? _GEN21910 : _GEN23234;
wire  _GEN23236 = io_x[46] ? _GEN23235 : _GEN23230;
wire  _GEN23237 = io_x[18] ? _GEN23236 : _GEN23224;
wire  _GEN23238 = io_x[49] ? _GEN23237 : _GEN23196;
wire  _GEN23239 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23240 = io_x[27] ? _GEN21739 : _GEN23239;
wire  _GEN23241 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23242 = io_x[27] ? _GEN23241 : _GEN21739;
wire  _GEN23243 = io_x[29] ? _GEN23242 : _GEN23240;
wire  _GEN23244 = io_x[75] ? _GEN21758 : _GEN23243;
wire  _GEN23245 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN23246 = io_x[75] ? _GEN21758 : _GEN23245;
wire  _GEN23247 = io_x[38] ? _GEN23246 : _GEN23244;
wire  _GEN23248 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23249 = io_x[27] ? _GEN21750 : _GEN23248;
wire  _GEN23250 = io_x[29] ? _GEN23249 : _GEN21744;
wire  _GEN23251 = io_x[75] ? _GEN21758 : _GEN23250;
wire  _GEN23252 = io_x[38] ? _GEN23251 : _GEN21833;
wire  _GEN23253 = io_x[34] ? _GEN23252 : _GEN23247;
wire  _GEN23254 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23255 = io_x[27] ? _GEN23254 : _GEN21750;
wire  _GEN23256 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23257 = io_x[27] ? _GEN23256 : _GEN21750;
wire  _GEN23258 = io_x[29] ? _GEN23257 : _GEN23255;
wire  _GEN23259 = io_x[75] ? _GEN21772 : _GEN23258;
wire  _GEN23260 = io_x[38] ? _GEN21871 : _GEN23259;
wire  _GEN23261 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23262 = io_x[27] ? _GEN21739 : _GEN23261;
wire  _GEN23263 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23264 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23265 = io_x[27] ? _GEN23264 : _GEN23263;
wire  _GEN23266 = io_x[29] ? _GEN23265 : _GEN23262;
wire  _GEN23267 = io_x[75] ? _GEN21758 : _GEN23266;
wire  _GEN23268 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23269 = io_x[27] ? _GEN23268 : _GEN21739;
wire  _GEN23270 = io_x[29] ? _GEN23269 : _GEN21743;
wire  _GEN23271 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23272 = io_x[27] ? _GEN21739 : _GEN23271;
wire  _GEN23273 = io_x[29] ? _GEN21743 : _GEN23272;
wire  _GEN23274 = io_x[75] ? _GEN23273 : _GEN23270;
wire  _GEN23275 = io_x[38] ? _GEN23274 : _GEN23267;
wire  _GEN23276 = io_x[34] ? _GEN23275 : _GEN23260;
wire  _GEN23277 = io_x[39] ? _GEN23276 : _GEN23253;
wire  _GEN23278 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23279 = io_x[27] ? _GEN21739 : _GEN23278;
wire  _GEN23280 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23281 = io_x[27] ? _GEN21739 : _GEN23280;
wire  _GEN23282 = io_x[29] ? _GEN23281 : _GEN23279;
wire  _GEN23283 = io_x[75] ? _GEN21758 : _GEN23282;
wire  _GEN23284 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23285 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23286 = io_x[27] ? _GEN23285 : _GEN23284;
wire  _GEN23287 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23288 = io_x[27] ? _GEN21750 : _GEN23287;
wire  _GEN23289 = io_x[29] ? _GEN23288 : _GEN23286;
wire  _GEN23290 = io_x[75] ? _GEN21758 : _GEN23289;
wire  _GEN23291 = io_x[38] ? _GEN23290 : _GEN23283;
wire  _GEN23292 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23293 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23294 = io_x[27] ? _GEN23293 : _GEN23292;
wire  _GEN23295 = io_x[29] ? _GEN21744 : _GEN23294;
wire  _GEN23296 = io_x[75] ? _GEN21758 : _GEN23295;
wire  _GEN23297 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23298 = io_x[27] ? _GEN21750 : _GEN23297;
wire  _GEN23299 = io_x[29] ? _GEN23298 : _GEN21743;
wire  _GEN23300 = io_x[75] ? _GEN21758 : _GEN23299;
wire  _GEN23301 = io_x[38] ? _GEN23300 : _GEN23296;
wire  _GEN23302 = io_x[34] ? _GEN23301 : _GEN23291;
wire  _GEN23303 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN23304 = io_x[29] ? _GEN23303 : _GEN21744;
wire  _GEN23305 = io_x[75] ? _GEN21758 : _GEN23304;
wire  _GEN23306 = io_x[38] ? _GEN21833 : _GEN23305;
wire  _GEN23307 = io_x[34] ? _GEN21927 : _GEN23306;
wire  _GEN23308 = io_x[39] ? _GEN23307 : _GEN23302;
wire  _GEN23309 = io_x[46] ? _GEN23308 : _GEN23277;
wire  _GEN23310 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23311 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN23312 = io_x[29] ? _GEN21744 : _GEN23311;
wire  _GEN23313 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23314 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23315 = io_x[27] ? _GEN23314 : _GEN23313;
wire  _GEN23316 = io_x[29] ? _GEN23315 : _GEN21743;
wire  _GEN23317 = io_x[75] ? _GEN23316 : _GEN23312;
wire  _GEN23318 = io_x[38] ? _GEN23317 : _GEN23310;
wire  _GEN23319 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23320 = io_x[27] ? _GEN23319 : _GEN21739;
wire  _GEN23321 = io_x[29] ? _GEN21743 : _GEN23320;
wire  _GEN23322 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23323 = io_x[27] ? _GEN23322 : _GEN21739;
wire  _GEN23324 = io_x[29] ? _GEN23323 : _GEN21743;
wire  _GEN23325 = io_x[75] ? _GEN23324 : _GEN23321;
wire  _GEN23326 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN23327 = io_x[38] ? _GEN23326 : _GEN23325;
wire  _GEN23328 = io_x[34] ? _GEN23327 : _GEN23318;
wire  _GEN23329 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23330 = io_x[27] ? _GEN23329 : _GEN21739;
wire  _GEN23331 = io_x[29] ? _GEN23330 : _GEN21743;
wire  _GEN23332 = io_x[75] ? _GEN21758 : _GEN23331;
wire  _GEN23333 = io_x[38] ? _GEN21871 : _GEN23332;
wire  _GEN23334 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23335 = io_x[27] ? _GEN23334 : _GEN21739;
wire  _GEN23336 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23337 = io_x[27] ? _GEN23336 : _GEN21739;
wire  _GEN23338 = io_x[29] ? _GEN23337 : _GEN23335;
wire  _GEN23339 = io_x[75] ? _GEN21772 : _GEN23338;
wire  _GEN23340 = io_x[38] ? _GEN21833 : _GEN23339;
wire  _GEN23341 = io_x[34] ? _GEN23340 : _GEN23333;
wire  _GEN23342 = io_x[39] ? _GEN23341 : _GEN23328;
wire  _GEN23343 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23344 = io_x[27] ? _GEN23343 : _GEN21739;
wire  _GEN23345 = io_x[29] ? _GEN23344 : _GEN21743;
wire  _GEN23346 = io_x[75] ? _GEN23345 : _GEN21758;
wire  _GEN23347 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23348 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23349 = io_x[27] ? _GEN23348 : _GEN23347;
wire  _GEN23350 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23351 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23352 = io_x[27] ? _GEN23351 : _GEN23350;
wire  _GEN23353 = io_x[29] ? _GEN23352 : _GEN23349;
wire  _GEN23354 = io_x[75] ? _GEN21772 : _GEN23353;
wire  _GEN23355 = io_x[38] ? _GEN23354 : _GEN23346;
wire  _GEN23356 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23357 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23358 = io_x[27] ? _GEN23357 : _GEN23356;
wire  _GEN23359 = io_x[29] ? _GEN21743 : _GEN23358;
wire  _GEN23360 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23361 = io_x[27] ? _GEN23360 : _GEN21739;
wire  _GEN23362 = io_x[29] ? _GEN23361 : _GEN21743;
wire  _GEN23363 = io_x[75] ? _GEN23362 : _GEN23359;
wire  _GEN23364 = io_x[38] ? _GEN21833 : _GEN23363;
wire  _GEN23365 = io_x[34] ? _GEN23364 : _GEN23355;
wire  _GEN23366 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN23367 = io_x[75] ? _GEN23366 : _GEN21758;
wire  _GEN23368 = io_x[38] ? _GEN21833 : _GEN23367;
wire  _GEN23369 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23370 = io_x[38] ? _GEN23369 : _GEN21833;
wire  _GEN23371 = io_x[34] ? _GEN23370 : _GEN23368;
wire  _GEN23372 = io_x[39] ? _GEN23371 : _GEN23365;
wire  _GEN23373 = io_x[46] ? _GEN23372 : _GEN23342;
wire  _GEN23374 = io_x[18] ? _GEN23373 : _GEN23309;
wire  _GEN23375 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN23376 = io_x[29] ? _GEN23375 : _GEN21743;
wire  _GEN23377 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23378 = io_x[27] ? _GEN23377 : _GEN21739;
wire  _GEN23379 = io_x[29] ? _GEN23378 : _GEN21743;
wire  _GEN23380 = io_x[75] ? _GEN23379 : _GEN23376;
wire  _GEN23381 = io_x[38] ? _GEN23380 : _GEN21871;
wire  _GEN23382 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23383 = io_x[38] ? _GEN23382 : _GEN21871;
wire  _GEN23384 = io_x[34] ? _GEN23383 : _GEN23381;
wire  _GEN23385 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23386 = io_x[27] ? _GEN23385 : _GEN21739;
wire  _GEN23387 = io_x[29] ? _GEN23386 : _GEN21743;
wire  _GEN23388 = io_x[75] ? _GEN23387 : _GEN21772;
wire  _GEN23389 = io_x[38] ? _GEN21833 : _GEN23388;
wire  _GEN23390 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN23391 = io_x[38] ? _GEN21833 : _GEN23390;
wire  _GEN23392 = io_x[34] ? _GEN23391 : _GEN23389;
wire  _GEN23393 = io_x[39] ? _GEN23392 : _GEN23384;
wire  _GEN23394 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23395 = io_x[27] ? _GEN23394 : _GEN21739;
wire  _GEN23396 = io_x[29] ? _GEN21743 : _GEN23395;
wire  _GEN23397 = io_x[75] ? _GEN21758 : _GEN23396;
wire  _GEN23398 = io_x[38] ? _GEN21833 : _GEN23397;
wire  _GEN23399 = io_x[34] ? _GEN21927 : _GEN23398;
wire  _GEN23400 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23401 = io_x[27] ? _GEN23400 : _GEN21739;
wire  _GEN23402 = io_x[29] ? _GEN23401 : _GEN21743;
wire  _GEN23403 = io_x[75] ? _GEN23402 : _GEN21758;
wire  _GEN23404 = io_x[38] ? _GEN21833 : _GEN23403;
wire  _GEN23405 = io_x[34] ? _GEN23404 : _GEN21927;
wire  _GEN23406 = io_x[39] ? _GEN23405 : _GEN23399;
wire  _GEN23407 = io_x[46] ? _GEN23406 : _GEN23393;
wire  _GEN23408 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN23409 = io_x[75] ? _GEN21758 : _GEN23408;
wire  _GEN23410 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN23411 = io_x[38] ? _GEN23410 : _GEN23409;
wire  _GEN23412 = io_x[34] ? _GEN23411 : _GEN21927;
wire  _GEN23413 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23414 = io_x[27] ? _GEN23413 : _GEN21739;
wire  _GEN23415 = io_x[29] ? _GEN23414 : _GEN21743;
wire  _GEN23416 = io_x[75] ? _GEN23415 : _GEN21772;
wire  _GEN23417 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN23418 = io_x[38] ? _GEN23417 : _GEN23416;
wire  _GEN23419 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23420 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23421 = io_x[27] ? _GEN23420 : _GEN23419;
wire  _GEN23422 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23423 = io_x[27] ? _GEN23422 : _GEN21750;
wire  _GEN23424 = io_x[29] ? _GEN23423 : _GEN23421;
wire  _GEN23425 = io_x[75] ? _GEN23424 : _GEN21772;
wire  _GEN23426 = io_x[38] ? _GEN21833 : _GEN23425;
wire  _GEN23427 = io_x[34] ? _GEN23426 : _GEN23418;
wire  _GEN23428 = io_x[39] ? _GEN23427 : _GEN23412;
wire  _GEN23429 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN23430 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23431 = io_x[38] ? _GEN23430 : _GEN21833;
wire  _GEN23432 = io_x[34] ? _GEN23431 : _GEN23429;
wire  _GEN23433 = io_x[39] ? _GEN21910 : _GEN23432;
wire  _GEN23434 = io_x[46] ? _GEN23433 : _GEN23428;
wire  _GEN23435 = io_x[18] ? _GEN23434 : _GEN23407;
wire  _GEN23436 = io_x[49] ? _GEN23435 : _GEN23374;
wire  _GEN23437 = io_x[24] ? _GEN23436 : _GEN23238;
wire  _GEN23438 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN23439 = io_x[38] ? _GEN21833 : _GEN23438;
wire  _GEN23440 = io_x[34] ? _GEN21927 : _GEN23439;
wire  _GEN23441 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23442 = io_x[27] ? _GEN23441 : _GEN21750;
wire  _GEN23443 = io_x[29] ? _GEN21744 : _GEN23442;
wire  _GEN23444 = io_x[75] ? _GEN23443 : _GEN21758;
wire  _GEN23445 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23446 = io_x[38] ? _GEN23445 : _GEN23444;
wire  _GEN23447 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN23448 = io_x[29] ? _GEN21743 : _GEN23447;
wire  _GEN23449 = io_x[75] ? _GEN23448 : _GEN21758;
wire  _GEN23450 = io_x[38] ? _GEN21871 : _GEN23449;
wire  _GEN23451 = io_x[34] ? _GEN23450 : _GEN23446;
wire  _GEN23452 = io_x[39] ? _GEN23451 : _GEN23440;
wire  _GEN23453 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23454 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23455 = io_x[27] ? _GEN23454 : _GEN23453;
wire  _GEN23456 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23457 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23458 = io_x[27] ? _GEN23457 : _GEN23456;
wire  _GEN23459 = io_x[29] ? _GEN23458 : _GEN23455;
wire  _GEN23460 = io_x[75] ? _GEN21758 : _GEN23459;
wire  _GEN23461 = io_x[38] ? _GEN23460 : _GEN21833;
wire  _GEN23462 = io_x[34] ? _GEN21766 : _GEN23461;
wire  _GEN23463 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23464 = io_x[27] ? _GEN23463 : _GEN21739;
wire  _GEN23465 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23466 = io_x[27] ? _GEN23465 : _GEN21739;
wire  _GEN23467 = io_x[29] ? _GEN23466 : _GEN23464;
wire  _GEN23468 = io_x[75] ? _GEN21758 : _GEN23467;
wire  _GEN23469 = io_x[38] ? _GEN21871 : _GEN23468;
wire  _GEN23470 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23471 = io_x[27] ? _GEN23470 : _GEN21739;
wire  _GEN23472 = io_x[29] ? _GEN21743 : _GEN23471;
wire  _GEN23473 = io_x[75] ? _GEN21772 : _GEN23472;
wire  _GEN23474 = io_x[38] ? _GEN21871 : _GEN23473;
wire  _GEN23475 = io_x[34] ? _GEN23474 : _GEN23469;
wire  _GEN23476 = io_x[39] ? _GEN23475 : _GEN23462;
wire  _GEN23477 = io_x[46] ? _GEN23476 : _GEN23452;
wire  _GEN23478 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23479 = io_x[27] ? _GEN21739 : _GEN23478;
wire  _GEN23480 = io_x[29] ? _GEN23479 : _GEN21743;
wire  _GEN23481 = io_x[75] ? _GEN21772 : _GEN23480;
wire  _GEN23482 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN23483 = io_x[29] ? _GEN21743 : _GEN23482;
wire  _GEN23484 = io_x[75] ? _GEN21772 : _GEN23483;
wire  _GEN23485 = io_x[38] ? _GEN23484 : _GEN23481;
wire  _GEN23486 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN23487 = io_x[29] ? _GEN21744 : _GEN23486;
wire  _GEN23488 = io_x[75] ? _GEN21758 : _GEN23487;
wire  _GEN23489 = io_x[38] ? _GEN21833 : _GEN23488;
wire  _GEN23490 = io_x[34] ? _GEN23489 : _GEN23485;
wire  _GEN23491 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23492 = io_x[38] ? _GEN21833 : _GEN23491;
wire  _GEN23493 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN23494 = io_x[34] ? _GEN23493 : _GEN23492;
wire  _GEN23495 = io_x[39] ? _GEN23494 : _GEN23490;
wire  _GEN23496 = io_x[34] ? _GEN21766 : _GEN21927;
wire  _GEN23497 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN23498 = io_x[39] ? _GEN23497 : _GEN23496;
wire  _GEN23499 = io_x[46] ? _GEN23498 : _GEN23495;
wire  _GEN23500 = io_x[18] ? _GEN23499 : _GEN23477;
wire  _GEN23501 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN23502 = io_x[46] ? _GEN22145 : _GEN23501;
wire  _GEN23503 = 1'b0;
wire  _GEN23504 = io_x[18] ? _GEN23503 : _GEN23502;
wire  _GEN23505 = io_x[49] ? _GEN23504 : _GEN23500;
wire  _GEN23506 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN23507 = io_x[38] ? _GEN23506 : _GEN21833;
wire  _GEN23508 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23509 = io_x[27] ? _GEN23508 : _GEN21739;
wire  _GEN23510 = io_x[29] ? _GEN23509 : _GEN21743;
wire  _GEN23511 = io_x[75] ? _GEN23510 : _GEN21758;
wire  _GEN23512 = io_x[38] ? _GEN23511 : _GEN21833;
wire  _GEN23513 = io_x[34] ? _GEN23512 : _GEN23507;
wire  _GEN23514 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN23515 = io_x[75] ? _GEN23514 : _GEN21772;
wire  _GEN23516 = io_x[38] ? _GEN23515 : _GEN21833;
wire  _GEN23517 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN23518 = io_x[75] ? _GEN21758 : _GEN23517;
wire  _GEN23519 = io_x[38] ? _GEN21833 : _GEN23518;
wire  _GEN23520 = io_x[34] ? _GEN23519 : _GEN23516;
wire  _GEN23521 = io_x[39] ? _GEN23520 : _GEN23513;
wire  _GEN23522 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23523 = io_x[27] ? _GEN23522 : _GEN21739;
wire  _GEN23524 = io_x[29] ? _GEN23523 : _GEN21743;
wire  _GEN23525 = io_x[75] ? _GEN21772 : _GEN23524;
wire  _GEN23526 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23527 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23528 = io_x[27] ? _GEN23527 : _GEN23526;
wire  _GEN23529 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23530 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23531 = io_x[27] ? _GEN23530 : _GEN23529;
wire  _GEN23532 = io_x[29] ? _GEN23531 : _GEN23528;
wire  _GEN23533 = io_x[75] ? _GEN21758 : _GEN23532;
wire  _GEN23534 = io_x[38] ? _GEN23533 : _GEN23525;
wire  _GEN23535 = io_x[34] ? _GEN21766 : _GEN23534;
wire  _GEN23536 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23537 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23538 = io_x[27] ? _GEN23537 : _GEN23536;
wire  _GEN23539 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23540 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23541 = io_x[27] ? _GEN23540 : _GEN23539;
wire  _GEN23542 = io_x[29] ? _GEN23541 : _GEN23538;
wire  _GEN23543 = io_x[75] ? _GEN21758 : _GEN23542;
wire  _GEN23544 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23545 = io_x[27] ? _GEN23544 : _GEN21750;
wire  _GEN23546 = io_x[29] ? _GEN21743 : _GEN23545;
wire  _GEN23547 = io_x[75] ? _GEN21758 : _GEN23546;
wire  _GEN23548 = io_x[38] ? _GEN23547 : _GEN23543;
wire  _GEN23549 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23550 = io_x[27] ? _GEN23549 : _GEN21739;
wire  _GEN23551 = io_x[29] ? _GEN21743 : _GEN23550;
wire  _GEN23552 = io_x[75] ? _GEN21758 : _GEN23551;
wire  _GEN23553 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23554 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23555 = io_x[27] ? _GEN23554 : _GEN23553;
wire  _GEN23556 = io_x[29] ? _GEN23555 : _GEN21744;
wire  _GEN23557 = io_x[75] ? _GEN21772 : _GEN23556;
wire  _GEN23558 = io_x[38] ? _GEN23557 : _GEN23552;
wire  _GEN23559 = io_x[34] ? _GEN23558 : _GEN23548;
wire  _GEN23560 = io_x[39] ? _GEN23559 : _GEN23535;
wire  _GEN23561 = io_x[46] ? _GEN23560 : _GEN23521;
wire  _GEN23562 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23563 = io_x[27] ? _GEN23562 : _GEN21739;
wire  _GEN23564 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23565 = io_x[27] ? _GEN23564 : _GEN21739;
wire  _GEN23566 = io_x[29] ? _GEN23565 : _GEN23563;
wire  _GEN23567 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN23568 = io_x[29] ? _GEN21744 : _GEN23567;
wire  _GEN23569 = io_x[75] ? _GEN23568 : _GEN23566;
wire  _GEN23570 = io_x[38] ? _GEN21833 : _GEN23569;
wire  _GEN23571 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23572 = io_x[27] ? _GEN23571 : _GEN21739;
wire  _GEN23573 = io_x[29] ? _GEN23572 : _GEN21743;
wire  _GEN23574 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23575 = io_x[27] ? _GEN23574 : _GEN21739;
wire  _GEN23576 = io_x[29] ? _GEN21744 : _GEN23575;
wire  _GEN23577 = io_x[75] ? _GEN23576 : _GEN23573;
wire  _GEN23578 = io_x[38] ? _GEN21833 : _GEN23577;
wire  _GEN23579 = io_x[34] ? _GEN23578 : _GEN23570;
wire  _GEN23580 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN23581 = io_x[75] ? _GEN21772 : _GEN23580;
wire  _GEN23582 = io_x[38] ? _GEN21833 : _GEN23581;
wire  _GEN23583 = io_x[34] ? _GEN21927 : _GEN23582;
wire  _GEN23584 = io_x[39] ? _GEN23583 : _GEN23579;
wire  _GEN23585 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN23586 = io_x[75] ? _GEN23585 : _GEN21758;
wire  _GEN23587 = io_x[38] ? _GEN21833 : _GEN23586;
wire  _GEN23588 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN23589 = io_x[75] ? _GEN21758 : _GEN23588;
wire  _GEN23590 = io_x[38] ? _GEN21833 : _GEN23589;
wire  _GEN23591 = io_x[34] ? _GEN23590 : _GEN23587;
wire  _GEN23592 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23593 = io_x[38] ? _GEN23592 : _GEN21833;
wire  _GEN23594 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23595 = io_x[38] ? _GEN23594 : _GEN21833;
wire  _GEN23596 = io_x[34] ? _GEN23595 : _GEN23593;
wire  _GEN23597 = io_x[39] ? _GEN23596 : _GEN23591;
wire  _GEN23598 = io_x[46] ? _GEN23597 : _GEN23584;
wire  _GEN23599 = io_x[18] ? _GEN23598 : _GEN23561;
wire  _GEN23600 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN23601 = io_x[46] ? _GEN22145 : _GEN23600;
wire  _GEN23602 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN23603 = io_x[75] ? _GEN23602 : _GEN21758;
wire  _GEN23604 = io_x[38] ? _GEN23603 : _GEN21833;
wire  _GEN23605 = io_x[34] ? _GEN21927 : _GEN23604;
wire  _GEN23606 = io_x[39] ? _GEN23605 : _GEN21910;
wire  _GEN23607 = io_x[46] ? _GEN22145 : _GEN23606;
wire  _GEN23608 = io_x[18] ? _GEN23607 : _GEN23601;
wire  _GEN23609 = io_x[49] ? _GEN23608 : _GEN23599;
wire  _GEN23610 = io_x[24] ? _GEN23609 : _GEN23505;
wire  _GEN23611 = io_x[80] ? _GEN23610 : _GEN23437;
wire  _GEN23612 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23613 = io_x[27] ? _GEN23612 : _GEN21739;
wire  _GEN23614 = io_x[29] ? _GEN23613 : _GEN21743;
wire  _GEN23615 = io_x[75] ? _GEN21758 : _GEN23614;
wire  _GEN23616 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23617 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23618 = io_x[27] ? _GEN23617 : _GEN23616;
wire  _GEN23619 = io_x[29] ? _GEN23618 : _GEN21744;
wire  _GEN23620 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23621 = io_x[27] ? _GEN21739 : _GEN23620;
wire  _GEN23622 = io_x[29] ? _GEN21743 : _GEN23621;
wire  _GEN23623 = io_x[75] ? _GEN23622 : _GEN23619;
wire  _GEN23624 = io_x[38] ? _GEN23623 : _GEN23615;
wire  _GEN23625 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN23626 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23627 = io_x[27] ? _GEN23626 : _GEN21739;
wire  _GEN23628 = io_x[29] ? _GEN23627 : _GEN23625;
wire  _GEN23629 = io_x[75] ? _GEN21758 : _GEN23628;
wire  _GEN23630 = io_x[38] ? _GEN23629 : _GEN21833;
wire  _GEN23631 = io_x[34] ? _GEN23630 : _GEN23624;
wire  _GEN23632 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23633 = io_x[27] ? _GEN23632 : _GEN21739;
wire  _GEN23634 = io_x[29] ? _GEN23633 : _GEN21743;
wire  _GEN23635 = io_x[75] ? _GEN23634 : _GEN21772;
wire  _GEN23636 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23637 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23638 = io_x[27] ? _GEN23637 : _GEN23636;
wire  _GEN23639 = io_x[29] ? _GEN23638 : _GEN21744;
wire  _GEN23640 = io_x[75] ? _GEN21772 : _GEN23639;
wire  _GEN23641 = io_x[38] ? _GEN23640 : _GEN23635;
wire  _GEN23642 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23643 = io_x[27] ? _GEN23642 : _GEN21739;
wire  _GEN23644 = io_x[29] ? _GEN21743 : _GEN23643;
wire  _GEN23645 = io_x[75] ? _GEN21772 : _GEN23644;
wire  _GEN23646 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23647 = io_x[27] ? _GEN23646 : _GEN21739;
wire  _GEN23648 = io_x[29] ? _GEN23647 : _GEN21744;
wire  _GEN23649 = io_x[75] ? _GEN21758 : _GEN23648;
wire  _GEN23650 = io_x[38] ? _GEN23649 : _GEN23645;
wire  _GEN23651 = io_x[34] ? _GEN23650 : _GEN23641;
wire  _GEN23652 = io_x[39] ? _GEN23651 : _GEN23631;
wire  _GEN23653 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23654 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23655 = io_x[27] ? _GEN21739 : _GEN23654;
wire  _GEN23656 = io_x[29] ? _GEN21743 : _GEN23655;
wire  _GEN23657 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23658 = io_x[27] ? _GEN23657 : _GEN21739;
wire  _GEN23659 = io_x[29] ? _GEN23658 : _GEN21744;
wire  _GEN23660 = io_x[75] ? _GEN23659 : _GEN23656;
wire  _GEN23661 = io_x[38] ? _GEN23660 : _GEN23653;
wire  _GEN23662 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23663 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23664 = io_x[27] ? _GEN23663 : _GEN23662;
wire  _GEN23665 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23666 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23667 = io_x[27] ? _GEN23666 : _GEN23665;
wire  _GEN23668 = io_x[29] ? _GEN23667 : _GEN23664;
wire  _GEN23669 = io_x[75] ? _GEN21758 : _GEN23668;
wire  _GEN23670 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23671 = io_x[38] ? _GEN23670 : _GEN23669;
wire  _GEN23672 = io_x[34] ? _GEN23671 : _GEN23661;
wire  _GEN23673 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23674 = io_x[27] ? _GEN23673 : _GEN21739;
wire  _GEN23675 = io_x[29] ? _GEN23674 : _GEN21743;
wire  _GEN23676 = io_x[75] ? _GEN23675 : _GEN21758;
wire  _GEN23677 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23678 = io_x[27] ? _GEN23677 : _GEN21750;
wire  _GEN23679 = io_x[29] ? _GEN21743 : _GEN23678;
wire  _GEN23680 = io_x[75] ? _GEN23679 : _GEN21758;
wire  _GEN23681 = io_x[38] ? _GEN23680 : _GEN23676;
wire  _GEN23682 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN23683 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN23684 = io_x[75] ? _GEN23683 : _GEN23682;
wire  _GEN23685 = io_x[38] ? _GEN23684 : _GEN21833;
wire  _GEN23686 = io_x[34] ? _GEN23685 : _GEN23681;
wire  _GEN23687 = io_x[39] ? _GEN23686 : _GEN23672;
wire  _GEN23688 = io_x[46] ? _GEN23687 : _GEN23652;
wire  _GEN23689 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23690 = io_x[27] ? _GEN21739 : _GEN23689;
wire  _GEN23691 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23692 = io_x[27] ? _GEN23691 : _GEN21739;
wire  _GEN23693 = io_x[29] ? _GEN23692 : _GEN23690;
wire  _GEN23694 = io_x[75] ? _GEN21772 : _GEN23693;
wire  _GEN23695 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23696 = io_x[27] ? _GEN23695 : _GEN21739;
wire  _GEN23697 = io_x[29] ? _GEN23696 : _GEN21744;
wire  _GEN23698 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23699 = io_x[27] ? _GEN23698 : _GEN21739;
wire  _GEN23700 = io_x[29] ? _GEN23699 : _GEN21743;
wire  _GEN23701 = io_x[75] ? _GEN23700 : _GEN23697;
wire  _GEN23702 = io_x[38] ? _GEN23701 : _GEN23694;
wire  _GEN23703 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23704 = io_x[27] ? _GEN23703 : _GEN21739;
wire  _GEN23705 = io_x[29] ? _GEN23704 : _GEN21743;
wire  _GEN23706 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23707 = io_x[27] ? _GEN21739 : _GEN23706;
wire  _GEN23708 = io_x[29] ? _GEN21743 : _GEN23707;
wire  _GEN23709 = io_x[75] ? _GEN23708 : _GEN23705;
wire  _GEN23710 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23711 = io_x[27] ? _GEN23710 : _GEN21739;
wire  _GEN23712 = io_x[29] ? _GEN23711 : _GEN21743;
wire  _GEN23713 = io_x[75] ? _GEN21758 : _GEN23712;
wire  _GEN23714 = io_x[38] ? _GEN23713 : _GEN23709;
wire  _GEN23715 = io_x[34] ? _GEN23714 : _GEN23702;
wire  _GEN23716 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23717 = io_x[27] ? _GEN21739 : _GEN23716;
wire  _GEN23718 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23719 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23720 = io_x[27] ? _GEN23719 : _GEN23718;
wire  _GEN23721 = io_x[29] ? _GEN23720 : _GEN23717;
wire  _GEN23722 = io_x[75] ? _GEN21772 : _GEN23721;
wire  _GEN23723 = io_x[38] ? _GEN23722 : _GEN21871;
wire  _GEN23724 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23725 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23726 = io_x[27] ? _GEN23725 : _GEN23724;
wire  _GEN23727 = io_x[29] ? _GEN23726 : _GEN21743;
wire  _GEN23728 = io_x[75] ? _GEN21772 : _GEN23727;
wire  _GEN23729 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN23730 = io_x[75] ? _GEN21758 : _GEN23729;
wire  _GEN23731 = io_x[38] ? _GEN23730 : _GEN23728;
wire  _GEN23732 = io_x[34] ? _GEN23731 : _GEN23723;
wire  _GEN23733 = io_x[39] ? _GEN23732 : _GEN23715;
wire  _GEN23734 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23735 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23736 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23737 = io_x[27] ? _GEN23736 : _GEN23735;
wire  _GEN23738 = io_x[29] ? _GEN21743 : _GEN23737;
wire  _GEN23739 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23740 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23741 = io_x[27] ? _GEN23740 : _GEN23739;
wire  _GEN23742 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23743 = io_x[27] ? _GEN23742 : _GEN21739;
wire  _GEN23744 = io_x[29] ? _GEN23743 : _GEN23741;
wire  _GEN23745 = io_x[75] ? _GEN23744 : _GEN23738;
wire  _GEN23746 = io_x[38] ? _GEN23745 : _GEN23734;
wire  _GEN23747 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23748 = io_x[27] ? _GEN21750 : _GEN23747;
wire  _GEN23749 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23750 = io_x[27] ? _GEN21739 : _GEN23749;
wire  _GEN23751 = io_x[29] ? _GEN23750 : _GEN23748;
wire  _GEN23752 = io_x[75] ? _GEN21758 : _GEN23751;
wire  _GEN23753 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23754 = io_x[38] ? _GEN23753 : _GEN23752;
wire  _GEN23755 = io_x[34] ? _GEN23754 : _GEN23746;
wire  _GEN23756 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23757 = io_x[27] ? _GEN23756 : _GEN21739;
wire  _GEN23758 = io_x[29] ? _GEN21743 : _GEN23757;
wire  _GEN23759 = io_x[75] ? _GEN21758 : _GEN23758;
wire  _GEN23760 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23761 = io_x[38] ? _GEN23760 : _GEN23759;
wire  _GEN23762 = io_x[34] ? _GEN23761 : _GEN21927;
wire  _GEN23763 = io_x[39] ? _GEN23762 : _GEN23755;
wire  _GEN23764 = io_x[46] ? _GEN23763 : _GEN23733;
wire  _GEN23765 = io_x[18] ? _GEN23764 : _GEN23688;
wire  _GEN23766 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN23767 = io_x[34] ? _GEN21766 : _GEN23766;
wire  _GEN23768 = io_x[39] ? _GEN21910 : _GEN23767;
wire  _GEN23769 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23770 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23771 = io_x[38] ? _GEN23770 : _GEN23769;
wire  _GEN23772 = io_x[34] ? _GEN23771 : _GEN21766;
wire  _GEN23773 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN23774 = io_x[75] ? _GEN23773 : _GEN21758;
wire  _GEN23775 = io_x[38] ? _GEN21833 : _GEN23774;
wire  _GEN23776 = io_x[34] ? _GEN23775 : _GEN21766;
wire  _GEN23777 = io_x[39] ? _GEN23776 : _GEN23772;
wire  _GEN23778 = io_x[46] ? _GEN23777 : _GEN23768;
wire  _GEN23779 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23780 = io_x[27] ? _GEN23779 : _GEN21739;
wire  _GEN23781 = io_x[29] ? _GEN23780 : _GEN21743;
wire  _GEN23782 = io_x[75] ? _GEN21758 : _GEN23781;
wire  _GEN23783 = io_x[38] ? _GEN23782 : _GEN21871;
wire  _GEN23784 = io_x[34] ? _GEN23783 : _GEN21766;
wire  _GEN23785 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN23786 = io_x[39] ? _GEN23785 : _GEN23784;
wire  _GEN23787 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23788 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23789 = io_x[38] ? _GEN23788 : _GEN23787;
wire  _GEN23790 = io_x[34] ? _GEN23789 : _GEN21927;
wire  _GEN23791 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23792 = io_x[27] ? _GEN21739 : _GEN23791;
wire  _GEN23793 = io_x[29] ? _GEN21743 : _GEN23792;
wire  _GEN23794 = io_x[75] ? _GEN23793 : _GEN21758;
wire  _GEN23795 = io_x[38] ? _GEN23794 : _GEN21833;
wire  _GEN23796 = io_x[34] ? _GEN23795 : _GEN21927;
wire  _GEN23797 = io_x[39] ? _GEN23796 : _GEN23790;
wire  _GEN23798 = io_x[46] ? _GEN23797 : _GEN23786;
wire  _GEN23799 = io_x[18] ? _GEN23798 : _GEN23778;
wire  _GEN23800 = io_x[49] ? _GEN23799 : _GEN23765;
wire  _GEN23801 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23802 = io_x[27] ? _GEN23801 : _GEN21739;
wire  _GEN23803 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23804 = io_x[27] ? _GEN23803 : _GEN21750;
wire  _GEN23805 = io_x[29] ? _GEN23804 : _GEN23802;
wire  _GEN23806 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23807 = io_x[27] ? _GEN23806 : _GEN21739;
wire  _GEN23808 = io_x[29] ? _GEN21743 : _GEN23807;
wire  _GEN23809 = io_x[75] ? _GEN23808 : _GEN23805;
wire  _GEN23810 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23811 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23812 = io_x[27] ? _GEN23811 : _GEN23810;
wire  _GEN23813 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23814 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23815 = io_x[27] ? _GEN23814 : _GEN23813;
wire  _GEN23816 = io_x[29] ? _GEN23815 : _GEN23812;
wire  _GEN23817 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23818 = io_x[27] ? _GEN23817 : _GEN21739;
wire  _GEN23819 = io_x[29] ? _GEN23818 : _GEN21743;
wire  _GEN23820 = io_x[75] ? _GEN23819 : _GEN23816;
wire  _GEN23821 = io_x[38] ? _GEN23820 : _GEN23809;
wire  _GEN23822 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23823 = io_x[27] ? _GEN21739 : _GEN23822;
wire  _GEN23824 = io_x[29] ? _GEN21744 : _GEN23823;
wire  _GEN23825 = io_x[75] ? _GEN21758 : _GEN23824;
wire  _GEN23826 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23827 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23828 = io_x[27] ? _GEN23827 : _GEN23826;
wire  _GEN23829 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23830 = io_x[27] ? _GEN23829 : _GEN21739;
wire  _GEN23831 = io_x[29] ? _GEN23830 : _GEN23828;
wire  _GEN23832 = io_x[75] ? _GEN21758 : _GEN23831;
wire  _GEN23833 = io_x[38] ? _GEN23832 : _GEN23825;
wire  _GEN23834 = io_x[34] ? _GEN23833 : _GEN23821;
wire  _GEN23835 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN23836 = io_x[29] ? _GEN23835 : _GEN21743;
wire  _GEN23837 = io_x[75] ? _GEN23836 : _GEN21772;
wire  _GEN23838 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23839 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23840 = io_x[27] ? _GEN23839 : _GEN23838;
wire  _GEN23841 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23842 = io_x[27] ? _GEN23841 : _GEN21750;
wire  _GEN23843 = io_x[29] ? _GEN23842 : _GEN23840;
wire  _GEN23844 = io_x[75] ? _GEN21772 : _GEN23843;
wire  _GEN23845 = io_x[38] ? _GEN23844 : _GEN23837;
wire  _GEN23846 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23847 = io_x[27] ? _GEN23846 : _GEN21739;
wire  _GEN23848 = io_x[29] ? _GEN23847 : _GEN21743;
wire  _GEN23849 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23850 = io_x[27] ? _GEN23849 : _GEN21739;
wire  _GEN23851 = io_x[29] ? _GEN23850 : _GEN21743;
wire  _GEN23852 = io_x[75] ? _GEN23851 : _GEN23848;
wire  _GEN23853 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23854 = io_x[27] ? _GEN23853 : _GEN21739;
wire  _GEN23855 = io_x[29] ? _GEN23854 : _GEN21744;
wire  _GEN23856 = io_x[75] ? _GEN21758 : _GEN23855;
wire  _GEN23857 = io_x[38] ? _GEN23856 : _GEN23852;
wire  _GEN23858 = io_x[34] ? _GEN23857 : _GEN23845;
wire  _GEN23859 = io_x[39] ? _GEN23858 : _GEN23834;
wire  _GEN23860 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN23861 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23862 = io_x[27] ? _GEN21739 : _GEN23861;
wire  _GEN23863 = io_x[29] ? _GEN21743 : _GEN23862;
wire  _GEN23864 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23865 = io_x[27] ? _GEN23864 : _GEN21750;
wire  _GEN23866 = io_x[29] ? _GEN23865 : _GEN21744;
wire  _GEN23867 = io_x[75] ? _GEN23866 : _GEN23863;
wire  _GEN23868 = io_x[38] ? _GEN23867 : _GEN23860;
wire  _GEN23869 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23870 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23871 = io_x[27] ? _GEN23870 : _GEN23869;
wire  _GEN23872 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23873 = io_x[27] ? _GEN21739 : _GEN23872;
wire  _GEN23874 = io_x[29] ? _GEN23873 : _GEN23871;
wire  _GEN23875 = io_x[75] ? _GEN21758 : _GEN23874;
wire  _GEN23876 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN23877 = io_x[29] ? _GEN23876 : _GEN21743;
wire  _GEN23878 = io_x[75] ? _GEN21772 : _GEN23877;
wire  _GEN23879 = io_x[38] ? _GEN23878 : _GEN23875;
wire  _GEN23880 = io_x[34] ? _GEN23879 : _GEN23868;
wire  _GEN23881 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN23882 = io_x[75] ? _GEN21758 : _GEN23881;
wire  _GEN23883 = io_x[38] ? _GEN23882 : _GEN21871;
wire  _GEN23884 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN23885 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23886 = io_x[27] ? _GEN21750 : _GEN23885;
wire  _GEN23887 = io_x[29] ? _GEN23886 : _GEN21743;
wire  _GEN23888 = io_x[75] ? _GEN23887 : _GEN23884;
wire  _GEN23889 = io_x[38] ? _GEN23888 : _GEN21833;
wire  _GEN23890 = io_x[34] ? _GEN23889 : _GEN23883;
wire  _GEN23891 = io_x[39] ? _GEN23890 : _GEN23880;
wire  _GEN23892 = io_x[46] ? _GEN23891 : _GEN23859;
wire  _GEN23893 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23894 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23895 = io_x[27] ? _GEN23894 : _GEN23893;
wire  _GEN23896 = io_x[29] ? _GEN23895 : _GEN21743;
wire  _GEN23897 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23898 = io_x[27] ? _GEN23897 : _GEN21750;
wire  _GEN23899 = io_x[29] ? _GEN23898 : _GEN21744;
wire  _GEN23900 = io_x[75] ? _GEN23899 : _GEN23896;
wire  _GEN23901 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23902 = io_x[27] ? _GEN23901 : _GEN21739;
wire  _GEN23903 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23904 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23905 = io_x[27] ? _GEN23904 : _GEN23903;
wire  _GEN23906 = io_x[29] ? _GEN23905 : _GEN23902;
wire  _GEN23907 = io_x[75] ? _GEN21758 : _GEN23906;
wire  _GEN23908 = io_x[38] ? _GEN23907 : _GEN23900;
wire  _GEN23909 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23910 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23911 = io_x[27] ? _GEN23910 : _GEN23909;
wire  _GEN23912 = io_x[29] ? _GEN23911 : _GEN21744;
wire  _GEN23913 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN23914 = io_x[29] ? _GEN23913 : _GEN21743;
wire  _GEN23915 = io_x[75] ? _GEN23914 : _GEN23912;
wire  _GEN23916 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23917 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23918 = io_x[27] ? _GEN23917 : _GEN23916;
wire  _GEN23919 = io_x[29] ? _GEN23918 : _GEN21743;
wire  _GEN23920 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23921 = io_x[27] ? _GEN23920 : _GEN21739;
wire  _GEN23922 = io_x[29] ? _GEN23921 : _GEN21743;
wire  _GEN23923 = io_x[75] ? _GEN23922 : _GEN23919;
wire  _GEN23924 = io_x[38] ? _GEN23923 : _GEN23915;
wire  _GEN23925 = io_x[34] ? _GEN23924 : _GEN23908;
wire  _GEN23926 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23927 = io_x[27] ? _GEN23926 : _GEN21739;
wire  _GEN23928 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23929 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23930 = io_x[27] ? _GEN23929 : _GEN23928;
wire  _GEN23931 = io_x[29] ? _GEN23930 : _GEN23927;
wire  _GEN23932 = io_x[75] ? _GEN21772 : _GEN23931;
wire  _GEN23933 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23934 = io_x[27] ? _GEN23933 : _GEN21750;
wire  _GEN23935 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23936 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23937 = io_x[27] ? _GEN23936 : _GEN23935;
wire  _GEN23938 = io_x[29] ? _GEN23937 : _GEN23934;
wire  _GEN23939 = io_x[75] ? _GEN21772 : _GEN23938;
wire  _GEN23940 = io_x[38] ? _GEN23939 : _GEN23932;
wire  _GEN23941 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23942 = io_x[27] ? _GEN23941 : _GEN21750;
wire  _GEN23943 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23944 = io_x[27] ? _GEN23943 : _GEN21739;
wire  _GEN23945 = io_x[29] ? _GEN23944 : _GEN23942;
wire  _GEN23946 = io_x[75] ? _GEN21772 : _GEN23945;
wire  _GEN23947 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23948 = io_x[27] ? _GEN23947 : _GEN21750;
wire  _GEN23949 = io_x[29] ? _GEN23948 : _GEN21743;
wire  _GEN23950 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23951 = io_x[27] ? _GEN23950 : _GEN21739;
wire  _GEN23952 = io_x[29] ? _GEN23951 : _GEN21743;
wire  _GEN23953 = io_x[75] ? _GEN23952 : _GEN23949;
wire  _GEN23954 = io_x[38] ? _GEN23953 : _GEN23946;
wire  _GEN23955 = io_x[34] ? _GEN23954 : _GEN23940;
wire  _GEN23956 = io_x[39] ? _GEN23955 : _GEN23925;
wire  _GEN23957 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23958 = io_x[27] ? _GEN23957 : _GEN21739;
wire  _GEN23959 = io_x[29] ? _GEN21743 : _GEN23958;
wire  _GEN23960 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN23961 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23962 = io_x[27] ? _GEN23961 : _GEN21750;
wire  _GEN23963 = io_x[29] ? _GEN23962 : _GEN23960;
wire  _GEN23964 = io_x[75] ? _GEN23963 : _GEN23959;
wire  _GEN23965 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23966 = io_x[27] ? _GEN23965 : _GEN21739;
wire  _GEN23967 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23968 = io_x[27] ? _GEN21739 : _GEN23967;
wire  _GEN23969 = io_x[29] ? _GEN23968 : _GEN23966;
wire  _GEN23970 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23971 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23972 = io_x[27] ? _GEN23971 : _GEN23970;
wire  _GEN23973 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23974 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23975 = io_x[27] ? _GEN23974 : _GEN23973;
wire  _GEN23976 = io_x[29] ? _GEN23975 : _GEN23972;
wire  _GEN23977 = io_x[75] ? _GEN23976 : _GEN23969;
wire  _GEN23978 = io_x[38] ? _GEN23977 : _GEN23964;
wire  _GEN23979 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23980 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23981 = io_x[27] ? _GEN23980 : _GEN23979;
wire  _GEN23982 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23983 = io_x[27] ? _GEN23982 : _GEN21750;
wire  _GEN23984 = io_x[29] ? _GEN23983 : _GEN23981;
wire  _GEN23985 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23986 = io_x[27] ? _GEN23985 : _GEN21739;
wire  _GEN23987 = io_x[29] ? _GEN23986 : _GEN21743;
wire  _GEN23988 = io_x[75] ? _GEN23987 : _GEN23984;
wire  _GEN23989 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23990 = io_x[27] ? _GEN21750 : _GEN23989;
wire  _GEN23991 = io_x[29] ? _GEN21744 : _GEN23990;
wire  _GEN23992 = io_x[75] ? _GEN23991 : _GEN21758;
wire  _GEN23993 = io_x[38] ? _GEN23992 : _GEN23988;
wire  _GEN23994 = io_x[34] ? _GEN23993 : _GEN23978;
wire  _GEN23995 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN23996 = io_x[27] ? _GEN23995 : _GEN21739;
wire  _GEN23997 = io_x[29] ? _GEN23996 : _GEN21743;
wire  _GEN23998 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN23999 = io_x[29] ? _GEN21744 : _GEN23998;
wire  _GEN24000 = io_x[75] ? _GEN23999 : _GEN23997;
wire  _GEN24001 = io_x[38] ? _GEN24000 : _GEN21833;
wire  _GEN24002 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24003 = io_x[27] ? _GEN21739 : _GEN24002;
wire  _GEN24004 = io_x[29] ? _GEN24003 : _GEN21743;
wire  _GEN24005 = io_x[75] ? _GEN21772 : _GEN24004;
wire  _GEN24006 = io_x[38] ? _GEN24005 : _GEN21833;
wire  _GEN24007 = io_x[34] ? _GEN24006 : _GEN24001;
wire  _GEN24008 = io_x[39] ? _GEN24007 : _GEN23994;
wire  _GEN24009 = io_x[46] ? _GEN24008 : _GEN23956;
wire  _GEN24010 = io_x[18] ? _GEN24009 : _GEN23892;
wire  _GEN24011 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN24012 = io_x[75] ? _GEN21758 : _GEN24011;
wire  _GEN24013 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24014 = io_x[27] ? _GEN24013 : _GEN21750;
wire  _GEN24015 = io_x[29] ? _GEN24014 : _GEN21743;
wire  _GEN24016 = io_x[75] ? _GEN21772 : _GEN24015;
wire  _GEN24017 = io_x[38] ? _GEN24016 : _GEN24012;
wire  _GEN24018 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24019 = io_x[29] ? _GEN24018 : _GEN21744;
wire  _GEN24020 = io_x[75] ? _GEN21772 : _GEN24019;
wire  _GEN24021 = io_x[38] ? _GEN24020 : _GEN21833;
wire  _GEN24022 = io_x[34] ? _GEN24021 : _GEN24017;
wire  _GEN24023 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24024 = io_x[27] ? _GEN24023 : _GEN21739;
wire  _GEN24025 = io_x[29] ? _GEN24024 : _GEN21743;
wire  _GEN24026 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24027 = io_x[29] ? _GEN24026 : _GEN21743;
wire  _GEN24028 = io_x[75] ? _GEN24027 : _GEN24025;
wire  _GEN24029 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24030 = io_x[38] ? _GEN24029 : _GEN24028;
wire  _GEN24031 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24032 = io_x[27] ? _GEN21739 : _GEN24031;
wire  _GEN24033 = io_x[29] ? _GEN21743 : _GEN24032;
wire  _GEN24034 = io_x[75] ? _GEN21758 : _GEN24033;
wire  _GEN24035 = io_x[38] ? _GEN21833 : _GEN24034;
wire  _GEN24036 = io_x[34] ? _GEN24035 : _GEN24030;
wire  _GEN24037 = io_x[39] ? _GEN24036 : _GEN24022;
wire  _GEN24038 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24039 = io_x[27] ? _GEN21739 : _GEN24038;
wire  _GEN24040 = io_x[29] ? _GEN21744 : _GEN24039;
wire  _GEN24041 = io_x[75] ? _GEN24040 : _GEN21772;
wire  _GEN24042 = io_x[38] ? _GEN21871 : _GEN24041;
wire  _GEN24043 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24044 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24045 = io_x[27] ? _GEN21739 : _GEN24044;
wire  _GEN24046 = io_x[29] ? _GEN21744 : _GEN24045;
wire  _GEN24047 = io_x[75] ? _GEN24046 : _GEN21758;
wire  _GEN24048 = io_x[38] ? _GEN24047 : _GEN24043;
wire  _GEN24049 = io_x[34] ? _GEN24048 : _GEN24042;
wire  _GEN24050 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24051 = io_x[38] ? _GEN21833 : _GEN24050;
wire  _GEN24052 = io_x[34] ? _GEN24051 : _GEN21927;
wire  _GEN24053 = io_x[39] ? _GEN24052 : _GEN24049;
wire  _GEN24054 = io_x[46] ? _GEN24053 : _GEN24037;
wire  _GEN24055 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24056 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24057 = io_x[27] ? _GEN24056 : _GEN21739;
wire  _GEN24058 = io_x[29] ? _GEN24057 : _GEN24055;
wire  _GEN24059 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24060 = io_x[29] ? _GEN21743 : _GEN24059;
wire  _GEN24061 = io_x[75] ? _GEN24060 : _GEN24058;
wire  _GEN24062 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24063 = io_x[27] ? _GEN21750 : _GEN24062;
wire  _GEN24064 = io_x[29] ? _GEN24063 : _GEN21743;
wire  _GEN24065 = io_x[75] ? _GEN24064 : _GEN21772;
wire  _GEN24066 = io_x[38] ? _GEN24065 : _GEN24061;
wire  _GEN24067 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24068 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24069 = io_x[27] ? _GEN24068 : _GEN24067;
wire  _GEN24070 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24071 = io_x[27] ? _GEN24070 : _GEN21739;
wire  _GEN24072 = io_x[29] ? _GEN24071 : _GEN24069;
wire  _GEN24073 = io_x[75] ? _GEN24072 : _GEN21772;
wire  _GEN24074 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24075 = io_x[27] ? _GEN24074 : _GEN21739;
wire  _GEN24076 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24077 = io_x[27] ? _GEN24076 : _GEN21739;
wire  _GEN24078 = io_x[29] ? _GEN24077 : _GEN24075;
wire  _GEN24079 = io_x[75] ? _GEN21772 : _GEN24078;
wire  _GEN24080 = io_x[38] ? _GEN24079 : _GEN24073;
wire  _GEN24081 = io_x[34] ? _GEN24080 : _GEN24066;
wire  _GEN24082 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24083 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24084 = io_x[27] ? _GEN24083 : _GEN21739;
wire  _GEN24085 = io_x[29] ? _GEN24084 : _GEN21744;
wire  _GEN24086 = io_x[75] ? _GEN21758 : _GEN24085;
wire  _GEN24087 = io_x[38] ? _GEN24086 : _GEN24082;
wire  _GEN24088 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24089 = io_x[27] ? _GEN24088 : _GEN21739;
wire  _GEN24090 = io_x[29] ? _GEN21743 : _GEN24089;
wire  _GEN24091 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24092 = io_x[27] ? _GEN24091 : _GEN21739;
wire  _GEN24093 = io_x[29] ? _GEN24092 : _GEN21743;
wire  _GEN24094 = io_x[75] ? _GEN24093 : _GEN24090;
wire  _GEN24095 = io_x[38] ? _GEN21833 : _GEN24094;
wire  _GEN24096 = io_x[34] ? _GEN24095 : _GEN24087;
wire  _GEN24097 = io_x[39] ? _GEN24096 : _GEN24081;
wire  _GEN24098 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24099 = io_x[27] ? _GEN21739 : _GEN24098;
wire  _GEN24100 = io_x[29] ? _GEN24099 : _GEN21743;
wire  _GEN24101 = io_x[75] ? _GEN24100 : _GEN21772;
wire  _GEN24102 = io_x[38] ? _GEN21871 : _GEN24101;
wire  _GEN24103 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24104 = io_x[27] ? _GEN21739 : _GEN24103;
wire  _GEN24105 = io_x[29] ? _GEN21743 : _GEN24104;
wire  _GEN24106 = io_x[75] ? _GEN21772 : _GEN24105;
wire  _GEN24107 = io_x[38] ? _GEN24106 : _GEN21833;
wire  _GEN24108 = io_x[34] ? _GEN24107 : _GEN24102;
wire  _GEN24109 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24110 = io_x[27] ? _GEN24109 : _GEN21750;
wire  _GEN24111 = io_x[29] ? _GEN24110 : _GEN21744;
wire  _GEN24112 = io_x[75] ? _GEN24111 : _GEN21758;
wire  _GEN24113 = io_x[38] ? _GEN24112 : _GEN21833;
wire  _GEN24114 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24115 = io_x[75] ? _GEN24114 : _GEN21758;
wire  _GEN24116 = io_x[38] ? _GEN21833 : _GEN24115;
wire  _GEN24117 = io_x[34] ? _GEN24116 : _GEN24113;
wire  _GEN24118 = io_x[39] ? _GEN24117 : _GEN24108;
wire  _GEN24119 = io_x[46] ? _GEN24118 : _GEN24097;
wire  _GEN24120 = io_x[18] ? _GEN24119 : _GEN24054;
wire  _GEN24121 = io_x[49] ? _GEN24120 : _GEN24010;
wire  _GEN24122 = io_x[24] ? _GEN24121 : _GEN23800;
wire  _GEN24123 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24124 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24125 = io_x[27] ? _GEN24124 : _GEN24123;
wire  _GEN24126 = io_x[29] ? _GEN21743 : _GEN24125;
wire  _GEN24127 = io_x[75] ? _GEN24126 : _GEN21758;
wire  _GEN24128 = io_x[38] ? _GEN21871 : _GEN24127;
wire  _GEN24129 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24130 = io_x[27] ? _GEN21739 : _GEN24129;
wire  _GEN24131 = io_x[29] ? _GEN24130 : _GEN21743;
wire  _GEN24132 = io_x[75] ? _GEN24131 : _GEN21758;
wire  _GEN24133 = io_x[38] ? _GEN21833 : _GEN24132;
wire  _GEN24134 = io_x[34] ? _GEN24133 : _GEN24128;
wire  _GEN24135 = io_x[39] ? _GEN21910 : _GEN24134;
wire  _GEN24136 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN24137 = io_x[34] ? _GEN21766 : _GEN24136;
wire  _GEN24138 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN24139 = io_x[38] ? _GEN21871 : _GEN24138;
wire  _GEN24140 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24141 = io_x[27] ? _GEN24140 : _GEN21739;
wire  _GEN24142 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24143 = io_x[27] ? _GEN21739 : _GEN24142;
wire  _GEN24144 = io_x[29] ? _GEN24143 : _GEN24141;
wire  _GEN24145 = io_x[75] ? _GEN21758 : _GEN24144;
wire  _GEN24146 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24147 = io_x[27] ? _GEN24146 : _GEN21739;
wire  _GEN24148 = io_x[29] ? _GEN21743 : _GEN24147;
wire  _GEN24149 = io_x[75] ? _GEN24148 : _GEN21772;
wire  _GEN24150 = io_x[38] ? _GEN24149 : _GEN24145;
wire  _GEN24151 = io_x[34] ? _GEN24150 : _GEN24139;
wire  _GEN24152 = io_x[39] ? _GEN24151 : _GEN24137;
wire  _GEN24153 = io_x[46] ? _GEN24152 : _GEN24135;
wire  _GEN24154 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24155 = io_x[27] ? _GEN21750 : _GEN24154;
wire  _GEN24156 = io_x[29] ? _GEN24155 : _GEN21744;
wire  _GEN24157 = io_x[75] ? _GEN21758 : _GEN24156;
wire  _GEN24158 = io_x[38] ? _GEN21871 : _GEN24157;
wire  _GEN24159 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24160 = io_x[29] ? _GEN24159 : _GEN21743;
wire  _GEN24161 = io_x[75] ? _GEN24160 : _GEN21772;
wire  _GEN24162 = io_x[38] ? _GEN21833 : _GEN24161;
wire  _GEN24163 = io_x[34] ? _GEN24162 : _GEN24158;
wire  _GEN24164 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24165 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24166 = io_x[27] ? _GEN24165 : _GEN24164;
wire  _GEN24167 = io_x[29] ? _GEN24166 : _GEN21743;
wire  _GEN24168 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24169 = io_x[27] ? _GEN21739 : _GEN24168;
wire  _GEN24170 = io_x[29] ? _GEN24169 : _GEN21743;
wire  _GEN24171 = io_x[75] ? _GEN24170 : _GEN24167;
wire  _GEN24172 = io_x[38] ? _GEN24171 : _GEN21833;
wire  _GEN24173 = io_x[34] ? _GEN21927 : _GEN24172;
wire  _GEN24174 = io_x[39] ? _GEN24173 : _GEN24163;
wire  _GEN24175 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN24176 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24177 = io_x[38] ? _GEN24176 : _GEN24175;
wire  _GEN24178 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN24179 = io_x[38] ? _GEN21871 : _GEN24178;
wire  _GEN24180 = io_x[34] ? _GEN24179 : _GEN24177;
wire  _GEN24181 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN24182 = io_x[34] ? _GEN24181 : _GEN21766;
wire  _GEN24183 = io_x[39] ? _GEN24182 : _GEN24180;
wire  _GEN24184 = io_x[46] ? _GEN24183 : _GEN24174;
wire  _GEN24185 = io_x[18] ? _GEN24184 : _GEN24153;
wire  _GEN24186 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN24187 = io_x[34] ? _GEN21927 : _GEN24186;
wire  _GEN24188 = io_x[39] ? _GEN22327 : _GEN24187;
wire  _GEN24189 = io_x[46] ? _GEN22145 : _GEN24188;
wire  _GEN24190 = 1'b1;
wire  _GEN24191 = io_x[18] ? _GEN24190 : _GEN24189;
wire  _GEN24192 = io_x[49] ? _GEN24191 : _GEN24185;
wire  _GEN24193 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN24194 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24195 = io_x[27] ? _GEN21739 : _GEN24194;
wire  _GEN24196 = io_x[29] ? _GEN24195 : _GEN21743;
wire  _GEN24197 = io_x[75] ? _GEN24196 : _GEN21758;
wire  _GEN24198 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN24199 = io_x[38] ? _GEN24198 : _GEN24197;
wire  _GEN24200 = io_x[34] ? _GEN24199 : _GEN24193;
wire  _GEN24201 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24202 = io_x[75] ? _GEN21758 : _GEN24201;
wire  _GEN24203 = io_x[38] ? _GEN24202 : _GEN21833;
wire  _GEN24204 = io_x[34] ? _GEN21766 : _GEN24203;
wire  _GEN24205 = io_x[39] ? _GEN24204 : _GEN24200;
wire  _GEN24206 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24207 = io_x[27] ? _GEN21750 : _GEN24206;
wire  _GEN24208 = io_x[29] ? _GEN21743 : _GEN24207;
wire  _GEN24209 = io_x[75] ? _GEN24208 : _GEN21758;
wire  _GEN24210 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24211 = io_x[27] ? _GEN24210 : _GEN21739;
wire  _GEN24212 = io_x[29] ? _GEN24211 : _GEN21743;
wire  _GEN24213 = io_x[75] ? _GEN21772 : _GEN24212;
wire  _GEN24214 = io_x[38] ? _GEN24213 : _GEN24209;
wire  _GEN24215 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN24216 = io_x[38] ? _GEN21871 : _GEN24215;
wire  _GEN24217 = io_x[34] ? _GEN24216 : _GEN24214;
wire  _GEN24218 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN24219 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24220 = io_x[27] ? _GEN21750 : _GEN24219;
wire  _GEN24221 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24222 = io_x[27] ? _GEN24221 : _GEN21739;
wire  _GEN24223 = io_x[29] ? _GEN24222 : _GEN24220;
wire  _GEN24224 = io_x[75] ? _GEN24223 : _GEN21772;
wire  _GEN24225 = io_x[38] ? _GEN24224 : _GEN24218;
wire  _GEN24226 = io_x[34] ? _GEN24225 : _GEN21766;
wire  _GEN24227 = io_x[39] ? _GEN24226 : _GEN24217;
wire  _GEN24228 = io_x[46] ? _GEN24227 : _GEN24205;
wire  _GEN24229 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24230 = io_x[27] ? _GEN24229 : _GEN21739;
wire  _GEN24231 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24232 = io_x[27] ? _GEN21739 : _GEN24231;
wire  _GEN24233 = io_x[29] ? _GEN24232 : _GEN24230;
wire  _GEN24234 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24235 = io_x[27] ? _GEN24234 : _GEN21739;
wire  _GEN24236 = io_x[29] ? _GEN24235 : _GEN21743;
wire  _GEN24237 = io_x[75] ? _GEN24236 : _GEN24233;
wire  _GEN24238 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24239 = io_x[27] ? _GEN24238 : _GEN21750;
wire  _GEN24240 = io_x[29] ? _GEN24239 : _GEN21743;
wire  _GEN24241 = io_x[75] ? _GEN21772 : _GEN24240;
wire  _GEN24242 = io_x[38] ? _GEN24241 : _GEN24237;
wire  _GEN24243 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24244 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24245 = io_x[29] ? _GEN24244 : _GEN24243;
wire  _GEN24246 = io_x[75] ? _GEN24245 : _GEN21772;
wire  _GEN24247 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24248 = io_x[27] ? _GEN24247 : _GEN21739;
wire  _GEN24249 = io_x[29] ? _GEN24248 : _GEN21744;
wire  _GEN24250 = io_x[75] ? _GEN21758 : _GEN24249;
wire  _GEN24251 = io_x[38] ? _GEN24250 : _GEN24246;
wire  _GEN24252 = io_x[34] ? _GEN24251 : _GEN24242;
wire  _GEN24253 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24254 = io_x[29] ? _GEN24253 : _GEN21743;
wire  _GEN24255 = io_x[75] ? _GEN21772 : _GEN24254;
wire  _GEN24256 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24257 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24258 = io_x[27] ? _GEN24257 : _GEN24256;
wire  _GEN24259 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24260 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24261 = io_x[27] ? _GEN24260 : _GEN24259;
wire  _GEN24262 = io_x[29] ? _GEN24261 : _GEN24258;
wire  _GEN24263 = io_x[75] ? _GEN21772 : _GEN24262;
wire  _GEN24264 = io_x[38] ? _GEN24263 : _GEN24255;
wire  _GEN24265 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24266 = io_x[29] ? _GEN24265 : _GEN21743;
wire  _GEN24267 = io_x[75] ? _GEN21758 : _GEN24266;
wire  _GEN24268 = io_x[38] ? _GEN21833 : _GEN24267;
wire  _GEN24269 = io_x[34] ? _GEN24268 : _GEN24264;
wire  _GEN24270 = io_x[39] ? _GEN24269 : _GEN24252;
wire  _GEN24271 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24272 = io_x[29] ? _GEN24271 : _GEN21743;
wire  _GEN24273 = io_x[75] ? _GEN24272 : _GEN21758;
wire  _GEN24274 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24275 = io_x[38] ? _GEN24274 : _GEN24273;
wire  _GEN24276 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24277 = io_x[75] ? _GEN21758 : _GEN24276;
wire  _GEN24278 = io_x[38] ? _GEN21871 : _GEN24277;
wire  _GEN24279 = io_x[34] ? _GEN24278 : _GEN24275;
wire  _GEN24280 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24281 = io_x[27] ? _GEN24280 : _GEN21750;
wire  _GEN24282 = io_x[29] ? _GEN21744 : _GEN24281;
wire  _GEN24283 = io_x[75] ? _GEN21758 : _GEN24282;
wire  _GEN24284 = io_x[38] ? _GEN24283 : _GEN21871;
wire  _GEN24285 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN24286 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24287 = io_x[29] ? _GEN21743 : _GEN24286;
wire  _GEN24288 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24289 = io_x[27] ? _GEN24288 : _GEN21739;
wire  _GEN24290 = io_x[29] ? _GEN24289 : _GEN21743;
wire  _GEN24291 = io_x[75] ? _GEN24290 : _GEN24287;
wire  _GEN24292 = io_x[38] ? _GEN24291 : _GEN24285;
wire  _GEN24293 = io_x[34] ? _GEN24292 : _GEN24284;
wire  _GEN24294 = io_x[39] ? _GEN24293 : _GEN24279;
wire  _GEN24295 = io_x[46] ? _GEN24294 : _GEN24270;
wire  _GEN24296 = io_x[18] ? _GEN24295 : _GEN24228;
wire  _GEN24297 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24298 = io_x[38] ? _GEN21833 : _GEN24297;
wire  _GEN24299 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN24300 = io_x[75] ? _GEN24299 : _GEN21758;
wire  _GEN24301 = io_x[38] ? _GEN24300 : _GEN21833;
wire  _GEN24302 = io_x[34] ? _GEN24301 : _GEN24298;
wire  _GEN24303 = io_x[39] ? _GEN22327 : _GEN24302;
wire  _GEN24304 = io_x[46] ? _GEN22145 : _GEN24303;
wire  _GEN24305 = io_x[39] ? _GEN22327 : _GEN21910;
wire  _GEN24306 = io_x[46] ? _GEN22145 : _GEN24305;
wire  _GEN24307 = io_x[18] ? _GEN24306 : _GEN24304;
wire  _GEN24308 = io_x[49] ? _GEN24307 : _GEN24296;
wire  _GEN24309 = io_x[24] ? _GEN24308 : _GEN24192;
wire  _GEN24310 = io_x[80] ? _GEN24309 : _GEN24122;
wire  _GEN24311 = io_x[16] ? _GEN24310 : _GEN23611;
wire  _GEN24312 = io_x[22] ? _GEN24311 : _GEN23096;
wire  _GEN24313 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24314 = io_x[27] ? _GEN21739 : _GEN24313;
wire  _GEN24315 = io_x[29] ? _GEN21743 : _GEN24314;
wire  _GEN24316 = io_x[75] ? _GEN21758 : _GEN24315;
wire  _GEN24317 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24318 = io_x[27] ? _GEN24317 : _GEN21739;
wire  _GEN24319 = io_x[29] ? _GEN24318 : _GEN21744;
wire  _GEN24320 = io_x[75] ? _GEN21772 : _GEN24319;
wire  _GEN24321 = io_x[38] ? _GEN24320 : _GEN24316;
wire  _GEN24322 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24323 = io_x[27] ? _GEN21739 : _GEN24322;
wire  _GEN24324 = io_x[29] ? _GEN21743 : _GEN24323;
wire  _GEN24325 = io_x[75] ? _GEN24324 : _GEN21772;
wire  _GEN24326 = io_x[38] ? _GEN24325 : _GEN21833;
wire  _GEN24327 = io_x[34] ? _GEN24326 : _GEN24321;
wire  _GEN24328 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24329 = io_x[27] ? _GEN21750 : _GEN24328;
wire  _GEN24330 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24331 = io_x[27] ? _GEN24330 : _GEN21750;
wire  _GEN24332 = io_x[29] ? _GEN24331 : _GEN24329;
wire  _GEN24333 = io_x[75] ? _GEN21758 : _GEN24332;
wire  _GEN24334 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24335 = io_x[75] ? _GEN21758 : _GEN24334;
wire  _GEN24336 = io_x[38] ? _GEN24335 : _GEN24333;
wire  _GEN24337 = io_x[34] ? _GEN24336 : _GEN21766;
wire  _GEN24338 = io_x[39] ? _GEN24337 : _GEN24327;
wire  _GEN24339 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24340 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24341 = io_x[27] ? _GEN24340 : _GEN24339;
wire  _GEN24342 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24343 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24344 = io_x[27] ? _GEN24343 : _GEN24342;
wire  _GEN24345 = io_x[29] ? _GEN24344 : _GEN24341;
wire  _GEN24346 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24347 = io_x[27] ? _GEN21739 : _GEN24346;
wire  _GEN24348 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24349 = io_x[27] ? _GEN24348 : _GEN21739;
wire  _GEN24350 = io_x[29] ? _GEN24349 : _GEN24347;
wire  _GEN24351 = io_x[75] ? _GEN24350 : _GEN24345;
wire  _GEN24352 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24353 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24354 = io_x[27] ? _GEN24353 : _GEN24352;
wire  _GEN24355 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24356 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24357 = io_x[27] ? _GEN24356 : _GEN24355;
wire  _GEN24358 = io_x[29] ? _GEN24357 : _GEN24354;
wire  _GEN24359 = io_x[75] ? _GEN21758 : _GEN24358;
wire  _GEN24360 = io_x[38] ? _GEN24359 : _GEN24351;
wire  _GEN24361 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24362 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24363 = io_x[27] ? _GEN24362 : _GEN24361;
wire  _GEN24364 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24365 = io_x[27] ? _GEN21750 : _GEN24364;
wire  _GEN24366 = io_x[29] ? _GEN24365 : _GEN24363;
wire  _GEN24367 = io_x[75] ? _GEN21758 : _GEN24366;
wire  _GEN24368 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24369 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24370 = io_x[27] ? _GEN24369 : _GEN24368;
wire  _GEN24371 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24372 = io_x[27] ? _GEN21739 : _GEN24371;
wire  _GEN24373 = io_x[29] ? _GEN24372 : _GEN24370;
wire  _GEN24374 = io_x[75] ? _GEN21758 : _GEN24373;
wire  _GEN24375 = io_x[38] ? _GEN24374 : _GEN24367;
wire  _GEN24376 = io_x[34] ? _GEN24375 : _GEN24360;
wire  _GEN24377 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24378 = io_x[27] ? _GEN21750 : _GEN24377;
wire  _GEN24379 = io_x[29] ? _GEN24378 : _GEN21744;
wire  _GEN24380 = io_x[75] ? _GEN24379 : _GEN21758;
wire  _GEN24381 = io_x[38] ? _GEN24380 : _GEN21833;
wire  _GEN24382 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24383 = io_x[38] ? _GEN24382 : _GEN21833;
wire  _GEN24384 = io_x[34] ? _GEN24383 : _GEN24381;
wire  _GEN24385 = io_x[39] ? _GEN24384 : _GEN24376;
wire  _GEN24386 = io_x[46] ? _GEN24385 : _GEN24338;
wire  _GEN24387 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24388 = io_x[27] ? _GEN21739 : _GEN24387;
wire  _GEN24389 = io_x[29] ? _GEN21743 : _GEN24388;
wire  _GEN24390 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24391 = io_x[29] ? _GEN21743 : _GEN24390;
wire  _GEN24392 = io_x[75] ? _GEN24391 : _GEN24389;
wire  _GEN24393 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24394 = io_x[27] ? _GEN21739 : _GEN24393;
wire  _GEN24395 = io_x[29] ? _GEN21743 : _GEN24394;
wire  _GEN24396 = io_x[75] ? _GEN21758 : _GEN24395;
wire  _GEN24397 = io_x[38] ? _GEN24396 : _GEN24392;
wire  _GEN24398 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24399 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24400 = io_x[27] ? _GEN24399 : _GEN21750;
wire  _GEN24401 = io_x[29] ? _GEN21744 : _GEN24400;
wire  _GEN24402 = io_x[75] ? _GEN21758 : _GEN24401;
wire  _GEN24403 = io_x[38] ? _GEN24402 : _GEN24398;
wire  _GEN24404 = io_x[34] ? _GEN24403 : _GEN24397;
wire  _GEN24405 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24406 = io_x[29] ? _GEN24405 : _GEN21744;
wire  _GEN24407 = io_x[75] ? _GEN21758 : _GEN24406;
wire  _GEN24408 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24409 = io_x[27] ? _GEN24408 : _GEN21739;
wire  _GEN24410 = io_x[29] ? _GEN24409 : _GEN21743;
wire  _GEN24411 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24412 = io_x[75] ? _GEN24411 : _GEN24410;
wire  _GEN24413 = io_x[38] ? _GEN24412 : _GEN24407;
wire  _GEN24414 = io_x[34] ? _GEN24413 : _GEN21766;
wire  _GEN24415 = io_x[39] ? _GEN24414 : _GEN24404;
wire  _GEN24416 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24417 = io_x[27] ? _GEN21739 : _GEN24416;
wire  _GEN24418 = io_x[29] ? _GEN21743 : _GEN24417;
wire  _GEN24419 = io_x[75] ? _GEN21758 : _GEN24418;
wire  _GEN24420 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24421 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24422 = io_x[27] ? _GEN24421 : _GEN24420;
wire  _GEN24423 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24424 = io_x[27] ? _GEN21750 : _GEN24423;
wire  _GEN24425 = io_x[29] ? _GEN24424 : _GEN24422;
wire  _GEN24426 = io_x[75] ? _GEN21758 : _GEN24425;
wire  _GEN24427 = io_x[38] ? _GEN24426 : _GEN24419;
wire  _GEN24428 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24429 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24430 = io_x[27] ? _GEN24429 : _GEN24428;
wire  _GEN24431 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24432 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24433 = io_x[27] ? _GEN24432 : _GEN24431;
wire  _GEN24434 = io_x[29] ? _GEN24433 : _GEN24430;
wire  _GEN24435 = io_x[75] ? _GEN21758 : _GEN24434;
wire  _GEN24436 = io_x[38] ? _GEN21833 : _GEN24435;
wire  _GEN24437 = io_x[34] ? _GEN24436 : _GEN24427;
wire  _GEN24438 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24439 = io_x[27] ? _GEN24438 : _GEN21739;
wire  _GEN24440 = io_x[29] ? _GEN21743 : _GEN24439;
wire  _GEN24441 = io_x[75] ? _GEN21758 : _GEN24440;
wire  _GEN24442 = io_x[38] ? _GEN24441 : _GEN21871;
wire  _GEN24443 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24444 = io_x[38] ? _GEN24443 : _GEN21833;
wire  _GEN24445 = io_x[34] ? _GEN24444 : _GEN24442;
wire  _GEN24446 = io_x[39] ? _GEN24445 : _GEN24437;
wire  _GEN24447 = io_x[46] ? _GEN24446 : _GEN24415;
wire  _GEN24448 = io_x[18] ? _GEN24447 : _GEN24386;
wire  _GEN24449 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24450 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24451 = io_x[27] ? _GEN24450 : _GEN21739;
wire  _GEN24452 = io_x[29] ? _GEN24451 : _GEN24449;
wire  _GEN24453 = io_x[75] ? _GEN21758 : _GEN24452;
wire  _GEN24454 = io_x[38] ? _GEN24453 : _GEN21833;
wire  _GEN24455 = io_x[34] ? _GEN21927 : _GEN24454;
wire  _GEN24456 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24457 = io_x[29] ? _GEN21743 : _GEN24456;
wire  _GEN24458 = io_x[75] ? _GEN21758 : _GEN24457;
wire  _GEN24459 = io_x[38] ? _GEN24458 : _GEN21833;
wire  _GEN24460 = io_x[34] ? _GEN21766 : _GEN24459;
wire  _GEN24461 = io_x[39] ? _GEN24460 : _GEN24455;
wire  _GEN24462 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24463 = io_x[27] ? _GEN21739 : _GEN24462;
wire  _GEN24464 = io_x[29] ? _GEN21743 : _GEN24463;
wire  _GEN24465 = io_x[75] ? _GEN21758 : _GEN24464;
wire  _GEN24466 = io_x[38] ? _GEN21871 : _GEN24465;
wire  _GEN24467 = io_x[34] ? _GEN21927 : _GEN24466;
wire  _GEN24468 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24469 = io_x[27] ? _GEN21739 : _GEN24468;
wire  _GEN24470 = io_x[29] ? _GEN21743 : _GEN24469;
wire  _GEN24471 = io_x[75] ? _GEN24470 : _GEN21758;
wire  _GEN24472 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24473 = io_x[27] ? _GEN21739 : _GEN24472;
wire  _GEN24474 = io_x[29] ? _GEN21743 : _GEN24473;
wire  _GEN24475 = io_x[75] ? _GEN24474 : _GEN21758;
wire  _GEN24476 = io_x[38] ? _GEN24475 : _GEN24471;
wire  _GEN24477 = io_x[34] ? _GEN24476 : _GEN21927;
wire  _GEN24478 = io_x[39] ? _GEN24477 : _GEN24467;
wire  _GEN24479 = io_x[46] ? _GEN24478 : _GEN24461;
wire  _GEN24480 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24481 = io_x[27] ? _GEN21739 : _GEN24480;
wire  _GEN24482 = io_x[29] ? _GEN21743 : _GEN24481;
wire  _GEN24483 = io_x[75] ? _GEN21758 : _GEN24482;
wire  _GEN24484 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24485 = io_x[27] ? _GEN21739 : _GEN24484;
wire  _GEN24486 = io_x[29] ? _GEN21743 : _GEN24485;
wire  _GEN24487 = io_x[75] ? _GEN21758 : _GEN24486;
wire  _GEN24488 = io_x[38] ? _GEN24487 : _GEN24483;
wire  _GEN24489 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24490 = io_x[75] ? _GEN21772 : _GEN24489;
wire  _GEN24491 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24492 = io_x[27] ? _GEN21739 : _GEN24491;
wire  _GEN24493 = io_x[29] ? _GEN21743 : _GEN24492;
wire  _GEN24494 = io_x[75] ? _GEN21772 : _GEN24493;
wire  _GEN24495 = io_x[38] ? _GEN24494 : _GEN24490;
wire  _GEN24496 = io_x[34] ? _GEN24495 : _GEN24488;
wire  _GEN24497 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24498 = io_x[27] ? _GEN21739 : _GEN24497;
wire  _GEN24499 = io_x[29] ? _GEN21744 : _GEN24498;
wire  _GEN24500 = io_x[75] ? _GEN24499 : _GEN21758;
wire  _GEN24501 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN24502 = io_x[38] ? _GEN24501 : _GEN24500;
wire  _GEN24503 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN24504 = io_x[34] ? _GEN24503 : _GEN24502;
wire  _GEN24505 = io_x[39] ? _GEN24504 : _GEN24496;
wire  _GEN24506 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24507 = io_x[38] ? _GEN21871 : _GEN24506;
wire  _GEN24508 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24509 = io_x[27] ? _GEN21739 : _GEN24508;
wire  _GEN24510 = io_x[29] ? _GEN21743 : _GEN24509;
wire  _GEN24511 = io_x[75] ? _GEN24510 : _GEN21758;
wire  _GEN24512 = io_x[38] ? _GEN21833 : _GEN24511;
wire  _GEN24513 = io_x[34] ? _GEN24512 : _GEN24507;
wire  _GEN24514 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24515 = io_x[27] ? _GEN21739 : _GEN24514;
wire  _GEN24516 = io_x[29] ? _GEN21743 : _GEN24515;
wire  _GEN24517 = io_x[75] ? _GEN24516 : _GEN21758;
wire  _GEN24518 = io_x[38] ? _GEN24517 : _GEN21833;
wire  _GEN24519 = io_x[34] ? _GEN24518 : _GEN21927;
wire  _GEN24520 = io_x[39] ? _GEN24519 : _GEN24513;
wire  _GEN24521 = io_x[46] ? _GEN24520 : _GEN24505;
wire  _GEN24522 = io_x[18] ? _GEN24521 : _GEN24479;
wire  _GEN24523 = io_x[49] ? _GEN24522 : _GEN24448;
wire  _GEN24524 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24525 = io_x[27] ? _GEN21739 : _GEN24524;
wire  _GEN24526 = io_x[29] ? _GEN24525 : _GEN21743;
wire  _GEN24527 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN24528 = io_x[75] ? _GEN24527 : _GEN24526;
wire  _GEN24529 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24530 = io_x[29] ? _GEN24529 : _GEN21743;
wire  _GEN24531 = io_x[75] ? _GEN21772 : _GEN24530;
wire  _GEN24532 = io_x[38] ? _GEN24531 : _GEN24528;
wire  _GEN24533 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24534 = io_x[27] ? _GEN21750 : _GEN24533;
wire  _GEN24535 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24536 = io_x[27] ? _GEN24535 : _GEN21750;
wire  _GEN24537 = io_x[29] ? _GEN24536 : _GEN24534;
wire  _GEN24538 = io_x[75] ? _GEN21758 : _GEN24537;
wire  _GEN24539 = io_x[38] ? _GEN24538 : _GEN21833;
wire  _GEN24540 = io_x[34] ? _GEN24539 : _GEN24532;
wire  _GEN24541 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24542 = io_x[29] ? _GEN24541 : _GEN21743;
wire  _GEN24543 = io_x[75] ? _GEN21772 : _GEN24542;
wire  _GEN24544 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24545 = io_x[75] ? _GEN21758 : _GEN24544;
wire  _GEN24546 = io_x[38] ? _GEN24545 : _GEN24543;
wire  _GEN24547 = io_x[34] ? _GEN24546 : _GEN21766;
wire  _GEN24548 = io_x[39] ? _GEN24547 : _GEN24540;
wire  _GEN24549 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24550 = io_x[27] ? _GEN21739 : _GEN24549;
wire  _GEN24551 = io_x[29] ? _GEN24550 : _GEN21743;
wire  _GEN24552 = io_x[75] ? _GEN21758 : _GEN24551;
wire  _GEN24553 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24554 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24555 = io_x[27] ? _GEN24554 : _GEN24553;
wire  _GEN24556 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24557 = io_x[27] ? _GEN21739 : _GEN24556;
wire  _GEN24558 = io_x[29] ? _GEN24557 : _GEN24555;
wire  _GEN24559 = io_x[75] ? _GEN21758 : _GEN24558;
wire  _GEN24560 = io_x[38] ? _GEN24559 : _GEN24552;
wire  _GEN24561 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24562 = io_x[27] ? _GEN21750 : _GEN24561;
wire  _GEN24563 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24564 = io_x[27] ? _GEN21739 : _GEN24563;
wire  _GEN24565 = io_x[29] ? _GEN24564 : _GEN24562;
wire  _GEN24566 = io_x[75] ? _GEN21758 : _GEN24565;
wire  _GEN24567 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24568 = io_x[29] ? _GEN24567 : _GEN21743;
wire  _GEN24569 = io_x[75] ? _GEN21758 : _GEN24568;
wire  _GEN24570 = io_x[38] ? _GEN24569 : _GEN24566;
wire  _GEN24571 = io_x[34] ? _GEN24570 : _GEN24560;
wire  _GEN24572 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24573 = io_x[38] ? _GEN24572 : _GEN21871;
wire  _GEN24574 = io_x[34] ? _GEN21927 : _GEN24573;
wire  _GEN24575 = io_x[39] ? _GEN24574 : _GEN24571;
wire  _GEN24576 = io_x[46] ? _GEN24575 : _GEN24548;
wire  _GEN24577 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24578 = io_x[27] ? _GEN24577 : _GEN21739;
wire  _GEN24579 = io_x[29] ? _GEN24578 : _GEN21743;
wire  _GEN24580 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24581 = io_x[29] ? _GEN24580 : _GEN21743;
wire  _GEN24582 = io_x[75] ? _GEN24581 : _GEN24579;
wire  _GEN24583 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24584 = io_x[27] ? _GEN24583 : _GEN21739;
wire  _GEN24585 = io_x[29] ? _GEN24584 : _GEN21744;
wire  _GEN24586 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24587 = io_x[27] ? _GEN21739 : _GEN24586;
wire  _GEN24588 = io_x[29] ? _GEN21743 : _GEN24587;
wire  _GEN24589 = io_x[75] ? _GEN24588 : _GEN24585;
wire  _GEN24590 = io_x[38] ? _GEN24589 : _GEN24582;
wire  _GEN24591 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24592 = io_x[29] ? _GEN24591 : _GEN21743;
wire  _GEN24593 = io_x[75] ? _GEN21758 : _GEN24592;
wire  _GEN24594 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24595 = io_x[27] ? _GEN24594 : _GEN21750;
wire  _GEN24596 = io_x[29] ? _GEN24595 : _GEN21743;
wire  _GEN24597 = io_x[75] ? _GEN21758 : _GEN24596;
wire  _GEN24598 = io_x[38] ? _GEN24597 : _GEN24593;
wire  _GEN24599 = io_x[34] ? _GEN24598 : _GEN24590;
wire  _GEN24600 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24601 = io_x[27] ? _GEN24600 : _GEN21739;
wire  _GEN24602 = io_x[29] ? _GEN24601 : _GEN21744;
wire  _GEN24603 = io_x[75] ? _GEN21772 : _GEN24602;
wire  _GEN24604 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24605 = io_x[75] ? _GEN21772 : _GEN24604;
wire  _GEN24606 = io_x[38] ? _GEN24605 : _GEN24603;
wire  _GEN24607 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24608 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24609 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24610 = io_x[27] ? _GEN24609 : _GEN24608;
wire  _GEN24611 = io_x[29] ? _GEN24610 : _GEN24607;
wire  _GEN24612 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24613 = io_x[27] ? _GEN24612 : _GEN21739;
wire  _GEN24614 = io_x[29] ? _GEN24613 : _GEN21744;
wire  _GEN24615 = io_x[75] ? _GEN24614 : _GEN24611;
wire  _GEN24616 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24617 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24618 = io_x[27] ? _GEN24617 : _GEN21739;
wire  _GEN24619 = io_x[29] ? _GEN24618 : _GEN24616;
wire  _GEN24620 = io_x[75] ? _GEN21758 : _GEN24619;
wire  _GEN24621 = io_x[38] ? _GEN24620 : _GEN24615;
wire  _GEN24622 = io_x[34] ? _GEN24621 : _GEN24606;
wire  _GEN24623 = io_x[39] ? _GEN24622 : _GEN24599;
wire  _GEN24624 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24625 = io_x[27] ? _GEN24624 : _GEN21739;
wire  _GEN24626 = io_x[29] ? _GEN24625 : _GEN21743;
wire  _GEN24627 = io_x[75] ? _GEN24626 : _GEN21758;
wire  _GEN24628 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24629 = io_x[27] ? _GEN21739 : _GEN24628;
wire  _GEN24630 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24631 = io_x[27] ? _GEN21739 : _GEN24630;
wire  _GEN24632 = io_x[29] ? _GEN24631 : _GEN24629;
wire  _GEN24633 = io_x[75] ? _GEN21758 : _GEN24632;
wire  _GEN24634 = io_x[38] ? _GEN24633 : _GEN24627;
wire  _GEN24635 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24636 = io_x[27] ? _GEN21739 : _GEN24635;
wire  _GEN24637 = io_x[29] ? _GEN21743 : _GEN24636;
wire  _GEN24638 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24639 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24640 = io_x[27] ? _GEN24639 : _GEN24638;
wire  _GEN24641 = io_x[29] ? _GEN24640 : _GEN21743;
wire  _GEN24642 = io_x[75] ? _GEN24641 : _GEN24637;
wire  _GEN24643 = io_x[38] ? _GEN21833 : _GEN24642;
wire  _GEN24644 = io_x[34] ? _GEN24643 : _GEN24634;
wire  _GEN24645 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24646 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24647 = io_x[75] ? _GEN21758 : _GEN24646;
wire  _GEN24648 = io_x[38] ? _GEN24647 : _GEN24645;
wire  _GEN24649 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24650 = io_x[29] ? _GEN24649 : _GEN21743;
wire  _GEN24651 = io_x[75] ? _GEN21772 : _GEN24650;
wire  _GEN24652 = io_x[38] ? _GEN24651 : _GEN21833;
wire  _GEN24653 = io_x[34] ? _GEN24652 : _GEN24648;
wire  _GEN24654 = io_x[39] ? _GEN24653 : _GEN24644;
wire  _GEN24655 = io_x[46] ? _GEN24654 : _GEN24623;
wire  _GEN24656 = io_x[18] ? _GEN24655 : _GEN24576;
wire  _GEN24657 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24658 = io_x[27] ? _GEN24657 : _GEN21739;
wire  _GEN24659 = io_x[29] ? _GEN24658 : _GEN21743;
wire  _GEN24660 = io_x[75] ? _GEN21758 : _GEN24659;
wire  _GEN24661 = io_x[38] ? _GEN24660 : _GEN21833;
wire  _GEN24662 = io_x[34] ? _GEN21927 : _GEN24661;
wire  _GEN24663 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24664 = io_x[27] ? _GEN24663 : _GEN21739;
wire  _GEN24665 = io_x[29] ? _GEN24664 : _GEN21743;
wire  _GEN24666 = io_x[75] ? _GEN21758 : _GEN24665;
wire  _GEN24667 = io_x[38] ? _GEN24666 : _GEN21833;
wire  _GEN24668 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24669 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24670 = io_x[27] ? _GEN24669 : _GEN24668;
wire  _GEN24671 = io_x[29] ? _GEN24670 : _GEN21743;
wire  _GEN24672 = io_x[75] ? _GEN24671 : _GEN21772;
wire  _GEN24673 = io_x[38] ? _GEN21833 : _GEN24672;
wire  _GEN24674 = io_x[34] ? _GEN24673 : _GEN24667;
wire  _GEN24675 = io_x[39] ? _GEN24674 : _GEN24662;
wire  _GEN24676 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24677 = io_x[27] ? _GEN21739 : _GEN24676;
wire  _GEN24678 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24679 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24680 = io_x[27] ? _GEN24679 : _GEN24678;
wire  _GEN24681 = io_x[29] ? _GEN24680 : _GEN24677;
wire  _GEN24682 = io_x[75] ? _GEN21758 : _GEN24681;
wire  _GEN24683 = io_x[38] ? _GEN21871 : _GEN24682;
wire  _GEN24684 = io_x[34] ? _GEN21927 : _GEN24683;
wire  _GEN24685 = io_x[39] ? _GEN21910 : _GEN24684;
wire  _GEN24686 = io_x[46] ? _GEN24685 : _GEN24675;
wire  _GEN24687 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24688 = io_x[27] ? _GEN24687 : _GEN21739;
wire  _GEN24689 = io_x[29] ? _GEN24688 : _GEN21743;
wire  _GEN24690 = io_x[75] ? _GEN21758 : _GEN24689;
wire  _GEN24691 = io_x[38] ? _GEN21833 : _GEN24690;
wire  _GEN24692 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24693 = io_x[29] ? _GEN24692 : _GEN21743;
wire  _GEN24694 = io_x[75] ? _GEN21758 : _GEN24693;
wire  _GEN24695 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24696 = io_x[27] ? _GEN21739 : _GEN24695;
wire  _GEN24697 = io_x[29] ? _GEN24696 : _GEN21743;
wire  _GEN24698 = io_x[75] ? _GEN21772 : _GEN24697;
wire  _GEN24699 = io_x[38] ? _GEN24698 : _GEN24694;
wire  _GEN24700 = io_x[34] ? _GEN24699 : _GEN24691;
wire  _GEN24701 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24702 = io_x[27] ? _GEN21739 : _GEN24701;
wire  _GEN24703 = io_x[29] ? _GEN24702 : _GEN21743;
wire  _GEN24704 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24705 = io_x[27] ? _GEN24704 : _GEN21739;
wire  _GEN24706 = io_x[29] ? _GEN24705 : _GEN21743;
wire  _GEN24707 = io_x[75] ? _GEN24706 : _GEN24703;
wire  _GEN24708 = io_x[38] ? _GEN24707 : _GEN21871;
wire  _GEN24709 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24710 = io_x[27] ? _GEN21750 : _GEN24709;
wire  _GEN24711 = io_x[29] ? _GEN24710 : _GEN21744;
wire  _GEN24712 = io_x[75] ? _GEN24711 : _GEN21772;
wire  _GEN24713 = io_x[38] ? _GEN21833 : _GEN24712;
wire  _GEN24714 = io_x[34] ? _GEN24713 : _GEN24708;
wire  _GEN24715 = io_x[39] ? _GEN24714 : _GEN24700;
wire  _GEN24716 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24717 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24718 = io_x[27] ? _GEN21739 : _GEN24717;
wire  _GEN24719 = io_x[29] ? _GEN24718 : _GEN24716;
wire  _GEN24720 = io_x[75] ? _GEN21772 : _GEN24719;
wire  _GEN24721 = io_x[38] ? _GEN21871 : _GEN24720;
wire  _GEN24722 = io_x[34] ? _GEN21927 : _GEN24721;
wire  _GEN24723 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24724 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24725 = io_x[27] ? _GEN24724 : _GEN21739;
wire  _GEN24726 = io_x[29] ? _GEN24725 : _GEN24723;
wire  _GEN24727 = io_x[75] ? _GEN24726 : _GEN21758;
wire  _GEN24728 = io_x[38] ? _GEN21833 : _GEN24727;
wire  _GEN24729 = io_x[34] ? _GEN24728 : _GEN21927;
wire  _GEN24730 = io_x[39] ? _GEN24729 : _GEN24722;
wire  _GEN24731 = io_x[46] ? _GEN24730 : _GEN24715;
wire  _GEN24732 = io_x[18] ? _GEN24731 : _GEN24686;
wire  _GEN24733 = io_x[49] ? _GEN24732 : _GEN24656;
wire  _GEN24734 = io_x[24] ? _GEN24733 : _GEN24523;
wire  _GEN24735 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24736 = io_x[29] ? _GEN24735 : _GEN21743;
wire  _GEN24737 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24738 = io_x[27] ? _GEN21739 : _GEN24737;
wire  _GEN24739 = io_x[29] ? _GEN21744 : _GEN24738;
wire  _GEN24740 = io_x[75] ? _GEN24739 : _GEN24736;
wire  _GEN24741 = io_x[38] ? _GEN21833 : _GEN24740;
wire  _GEN24742 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24743 = io_x[27] ? _GEN24742 : _GEN21739;
wire  _GEN24744 = io_x[29] ? _GEN21743 : _GEN24743;
wire  _GEN24745 = io_x[75] ? _GEN24744 : _GEN21758;
wire  _GEN24746 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24747 = io_x[75] ? _GEN21758 : _GEN24746;
wire  _GEN24748 = io_x[38] ? _GEN24747 : _GEN24745;
wire  _GEN24749 = io_x[34] ? _GEN24748 : _GEN24741;
wire  _GEN24750 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24751 = io_x[27] ? _GEN24750 : _GEN21750;
wire  _GEN24752 = io_x[29] ? _GEN21744 : _GEN24751;
wire  _GEN24753 = io_x[75] ? _GEN24752 : _GEN21758;
wire  _GEN24754 = io_x[38] ? _GEN21833 : _GEN24753;
wire  _GEN24755 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24756 = io_x[27] ? _GEN24755 : _GEN21739;
wire  _GEN24757 = io_x[29] ? _GEN21744 : _GEN24756;
wire  _GEN24758 = io_x[75] ? _GEN24757 : _GEN21758;
wire  _GEN24759 = io_x[38] ? _GEN21833 : _GEN24758;
wire  _GEN24760 = io_x[34] ? _GEN24759 : _GEN24754;
wire  _GEN24761 = io_x[39] ? _GEN24760 : _GEN24749;
wire  _GEN24762 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24763 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24764 = io_x[27] ? _GEN24763 : _GEN24762;
wire  _GEN24765 = io_x[29] ? _GEN21743 : _GEN24764;
wire  _GEN24766 = io_x[75] ? _GEN21772 : _GEN24765;
wire  _GEN24767 = io_x[38] ? _GEN24766 : _GEN21833;
wire  _GEN24768 = io_x[34] ? _GEN21766 : _GEN24767;
wire  _GEN24769 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24770 = io_x[27] ? _GEN24769 : _GEN21739;
wire  _GEN24771 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24772 = io_x[27] ? _GEN21739 : _GEN24771;
wire  _GEN24773 = io_x[29] ? _GEN24772 : _GEN24770;
wire  _GEN24774 = io_x[75] ? _GEN21772 : _GEN24773;
wire  _GEN24775 = io_x[38] ? _GEN21871 : _GEN24774;
wire  _GEN24776 = io_x[34] ? _GEN21927 : _GEN24775;
wire  _GEN24777 = io_x[39] ? _GEN24776 : _GEN24768;
wire  _GEN24778 = io_x[46] ? _GEN24777 : _GEN24761;
wire  _GEN24779 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24780 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24781 = io_x[27] ? _GEN24780 : _GEN24779;
wire  _GEN24782 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24783 = io_x[29] ? _GEN24782 : _GEN24781;
wire  _GEN24784 = io_x[75] ? _GEN21758 : _GEN24783;
wire  _GEN24785 = io_x[38] ? _GEN21833 : _GEN24784;
wire  _GEN24786 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN24787 = io_x[75] ? _GEN24786 : _GEN21772;
wire  _GEN24788 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24789 = io_x[27] ? _GEN21739 : _GEN24788;
wire  _GEN24790 = io_x[29] ? _GEN21743 : _GEN24789;
wire  _GEN24791 = io_x[75] ? _GEN24790 : _GEN21772;
wire  _GEN24792 = io_x[38] ? _GEN24791 : _GEN24787;
wire  _GEN24793 = io_x[34] ? _GEN24792 : _GEN24785;
wire  _GEN24794 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24795 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24796 = io_x[27] ? _GEN21739 : _GEN24795;
wire  _GEN24797 = io_x[29] ? _GEN21743 : _GEN24796;
wire  _GEN24798 = io_x[75] ? _GEN21758 : _GEN24797;
wire  _GEN24799 = io_x[38] ? _GEN24798 : _GEN24794;
wire  _GEN24800 = io_x[34] ? _GEN24799 : _GEN21766;
wire  _GEN24801 = io_x[39] ? _GEN24800 : _GEN24793;
wire  _GEN24802 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24803 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24804 = io_x[27] ? _GEN24803 : _GEN24802;
wire  _GEN24805 = io_x[29] ? _GEN21743 : _GEN24804;
wire  _GEN24806 = io_x[75] ? _GEN21758 : _GEN24805;
wire  _GEN24807 = io_x[38] ? _GEN24806 : _GEN21833;
wire  _GEN24808 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN24809 = io_x[34] ? _GEN24808 : _GEN24807;
wire  _GEN24810 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24811 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24812 = io_x[27] ? _GEN24811 : _GEN24810;
wire  _GEN24813 = io_x[29] ? _GEN21743 : _GEN24812;
wire  _GEN24814 = io_x[75] ? _GEN21758 : _GEN24813;
wire  _GEN24815 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24816 = io_x[75] ? _GEN21758 : _GEN24815;
wire  _GEN24817 = io_x[38] ? _GEN24816 : _GEN24814;
wire  _GEN24818 = io_x[34] ? _GEN24817 : _GEN21766;
wire  _GEN24819 = io_x[39] ? _GEN24818 : _GEN24809;
wire  _GEN24820 = io_x[46] ? _GEN24819 : _GEN24801;
wire  _GEN24821 = io_x[18] ? _GEN24820 : _GEN24778;
wire  _GEN24822 = io_x[18] ? _GEN24190 : _GEN23503;
wire  _GEN24823 = io_x[49] ? _GEN24822 : _GEN24821;
wire  _GEN24824 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24825 = io_x[75] ? _GEN24824 : _GEN21758;
wire  _GEN24826 = io_x[38] ? _GEN21833 : _GEN24825;
wire  _GEN24827 = io_x[34] ? _GEN21927 : _GEN24826;
wire  _GEN24828 = io_x[39] ? _GEN22327 : _GEN24827;
wire  _GEN24829 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24830 = io_x[27] ? _GEN24829 : _GEN21739;
wire  _GEN24831 = io_x[29] ? _GEN24830 : _GEN21743;
wire  _GEN24832 = io_x[75] ? _GEN21772 : _GEN24831;
wire  _GEN24833 = io_x[38] ? _GEN24832 : _GEN21833;
wire  _GEN24834 = io_x[34] ? _GEN21927 : _GEN24833;
wire  _GEN24835 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24836 = io_x[27] ? _GEN24835 : _GEN21739;
wire  _GEN24837 = io_x[29] ? _GEN24836 : _GEN21743;
wire  _GEN24838 = io_x[75] ? _GEN21772 : _GEN24837;
wire  _GEN24839 = io_x[38] ? _GEN21871 : _GEN24838;
wire  _GEN24840 = io_x[34] ? _GEN21927 : _GEN24839;
wire  _GEN24841 = io_x[39] ? _GEN24840 : _GEN24834;
wire  _GEN24842 = io_x[46] ? _GEN24841 : _GEN24828;
wire  _GEN24843 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24844 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24845 = io_x[27] ? _GEN24844 : _GEN24843;
wire  _GEN24846 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24847 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24848 = io_x[27] ? _GEN24847 : _GEN24846;
wire  _GEN24849 = io_x[29] ? _GEN24848 : _GEN24845;
wire  _GEN24850 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24851 = io_x[27] ? _GEN21750 : _GEN24850;
wire  _GEN24852 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24853 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24854 = io_x[27] ? _GEN24853 : _GEN24852;
wire  _GEN24855 = io_x[29] ? _GEN24854 : _GEN24851;
wire  _GEN24856 = io_x[75] ? _GEN24855 : _GEN24849;
wire  _GEN24857 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN24858 = io_x[38] ? _GEN24857 : _GEN24856;
wire  _GEN24859 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24860 = io_x[75] ? _GEN21758 : _GEN24859;
wire  _GEN24861 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24862 = io_x[27] ? _GEN24861 : _GEN21750;
wire  _GEN24863 = io_x[29] ? _GEN24862 : _GEN21744;
wire  _GEN24864 = io_x[75] ? _GEN21772 : _GEN24863;
wire  _GEN24865 = io_x[38] ? _GEN24864 : _GEN24860;
wire  _GEN24866 = io_x[34] ? _GEN24865 : _GEN24858;
wire  _GEN24867 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24868 = io_x[29] ? _GEN24867 : _GEN21744;
wire  _GEN24869 = io_x[75] ? _GEN24868 : _GEN21758;
wire  _GEN24870 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24871 = io_x[27] ? _GEN24870 : _GEN21739;
wire  _GEN24872 = io_x[29] ? _GEN24871 : _GEN21744;
wire  _GEN24873 = io_x[75] ? _GEN21758 : _GEN24872;
wire  _GEN24874 = io_x[38] ? _GEN24873 : _GEN24869;
wire  _GEN24875 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24876 = io_x[27] ? _GEN21750 : _GEN24875;
wire  _GEN24877 = io_x[29] ? _GEN24876 : _GEN21743;
wire  _GEN24878 = io_x[75] ? _GEN21758 : _GEN24877;
wire  _GEN24879 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24880 = io_x[27] ? _GEN24879 : _GEN21750;
wire  _GEN24881 = io_x[29] ? _GEN24880 : _GEN21743;
wire  _GEN24882 = io_x[75] ? _GEN21758 : _GEN24881;
wire  _GEN24883 = io_x[38] ? _GEN24882 : _GEN24878;
wire  _GEN24884 = io_x[34] ? _GEN24883 : _GEN24874;
wire  _GEN24885 = io_x[39] ? _GEN24884 : _GEN24866;
wire  _GEN24886 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24887 = io_x[27] ? _GEN21739 : _GEN24886;
wire  _GEN24888 = io_x[29] ? _GEN24887 : _GEN21743;
wire  _GEN24889 = io_x[75] ? _GEN24888 : _GEN21758;
wire  _GEN24890 = io_x[38] ? _GEN21833 : _GEN24889;
wire  _GEN24891 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24892 = io_x[27] ? _GEN21739 : _GEN24891;
wire  _GEN24893 = io_x[29] ? _GEN24892 : _GEN21743;
wire  _GEN24894 = io_x[75] ? _GEN21758 : _GEN24893;
wire  _GEN24895 = io_x[38] ? _GEN21833 : _GEN24894;
wire  _GEN24896 = io_x[34] ? _GEN24895 : _GEN24890;
wire  _GEN24897 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN24898 = io_x[29] ? _GEN24897 : _GEN21743;
wire  _GEN24899 = io_x[75] ? _GEN21772 : _GEN24898;
wire  _GEN24900 = io_x[38] ? _GEN21871 : _GEN24899;
wire  _GEN24901 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN24902 = io_x[29] ? _GEN24901 : _GEN21743;
wire  _GEN24903 = io_x[75] ? _GEN21772 : _GEN24902;
wire  _GEN24904 = io_x[38] ? _GEN24903 : _GEN21833;
wire  _GEN24905 = io_x[34] ? _GEN24904 : _GEN24900;
wire  _GEN24906 = io_x[39] ? _GEN24905 : _GEN24896;
wire  _GEN24907 = io_x[46] ? _GEN24906 : _GEN24885;
wire  _GEN24908 = io_x[18] ? _GEN24907 : _GEN24842;
wire  _GEN24909 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24910 = io_x[27] ? _GEN24909 : _GEN21739;
wire  _GEN24911 = io_x[29] ? _GEN24910 : _GEN21743;
wire  _GEN24912 = io_x[75] ? _GEN24911 : _GEN21758;
wire  _GEN24913 = io_x[38] ? _GEN24912 : _GEN21833;
wire  _GEN24914 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN24915 = io_x[34] ? _GEN24914 : _GEN24913;
wire  _GEN24916 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN24917 = io_x[34] ? _GEN21927 : _GEN24916;
wire  _GEN24918 = io_x[39] ? _GEN24917 : _GEN24915;
wire  _GEN24919 = io_x[46] ? _GEN22145 : _GEN24918;
wire  _GEN24920 = io_x[18] ? _GEN24919 : _GEN23503;
wire  _GEN24921 = io_x[49] ? _GEN24920 : _GEN24908;
wire  _GEN24922 = io_x[24] ? _GEN24921 : _GEN24823;
wire  _GEN24923 = io_x[80] ? _GEN24922 : _GEN24734;
wire  _GEN24924 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24925 = io_x[75] ? _GEN21758 : _GEN24924;
wire  _GEN24926 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24927 = io_x[27] ? _GEN21739 : _GEN24926;
wire  _GEN24928 = io_x[29] ? _GEN21743 : _GEN24927;
wire  _GEN24929 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24930 = io_x[27] ? _GEN21739 : _GEN24929;
wire  _GEN24931 = io_x[29] ? _GEN24930 : _GEN21743;
wire  _GEN24932 = io_x[75] ? _GEN24931 : _GEN24928;
wire  _GEN24933 = io_x[38] ? _GEN24932 : _GEN24925;
wire  _GEN24934 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24935 = io_x[27] ? _GEN21739 : _GEN24934;
wire  _GEN24936 = io_x[29] ? _GEN21744 : _GEN24935;
wire  _GEN24937 = io_x[75] ? _GEN21772 : _GEN24936;
wire  _GEN24938 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24939 = io_x[27] ? _GEN21739 : _GEN24938;
wire  _GEN24940 = io_x[29] ? _GEN21743 : _GEN24939;
wire  _GEN24941 = io_x[75] ? _GEN21758 : _GEN24940;
wire  _GEN24942 = io_x[38] ? _GEN24941 : _GEN24937;
wire  _GEN24943 = io_x[34] ? _GEN24942 : _GEN24933;
wire  _GEN24944 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24945 = io_x[27] ? _GEN24944 : _GEN21739;
wire  _GEN24946 = io_x[29] ? _GEN24945 : _GEN21744;
wire  _GEN24947 = io_x[75] ? _GEN21758 : _GEN24946;
wire  _GEN24948 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24949 = io_x[27] ? _GEN24948 : _GEN21739;
wire  _GEN24950 = io_x[29] ? _GEN24949 : _GEN21744;
wire  _GEN24951 = io_x[75] ? _GEN21758 : _GEN24950;
wire  _GEN24952 = io_x[38] ? _GEN24951 : _GEN24947;
wire  _GEN24953 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN24954 = io_x[75] ? _GEN24953 : _GEN21758;
wire  _GEN24955 = io_x[38] ? _GEN21871 : _GEN24954;
wire  _GEN24956 = io_x[34] ? _GEN24955 : _GEN24952;
wire  _GEN24957 = io_x[39] ? _GEN24956 : _GEN24943;
wire  _GEN24958 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24959 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24960 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24961 = io_x[27] ? _GEN24960 : _GEN24959;
wire  _GEN24962 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24963 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24964 = io_x[27] ? _GEN24963 : _GEN24962;
wire  _GEN24965 = io_x[29] ? _GEN24964 : _GEN24961;
wire  _GEN24966 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN24967 = io_x[75] ? _GEN24966 : _GEN24965;
wire  _GEN24968 = io_x[38] ? _GEN24967 : _GEN24958;
wire  _GEN24969 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24970 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24971 = io_x[27] ? _GEN24970 : _GEN24969;
wire  _GEN24972 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24973 = io_x[27] ? _GEN21739 : _GEN24972;
wire  _GEN24974 = io_x[29] ? _GEN24973 : _GEN24971;
wire  _GEN24975 = io_x[75] ? _GEN21772 : _GEN24974;
wire  _GEN24976 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24977 = io_x[27] ? _GEN24976 : _GEN21739;
wire  _GEN24978 = io_x[29] ? _GEN24977 : _GEN21743;
wire  _GEN24979 = io_x[75] ? _GEN24978 : _GEN21758;
wire  _GEN24980 = io_x[38] ? _GEN24979 : _GEN24975;
wire  _GEN24981 = io_x[34] ? _GEN24980 : _GEN24968;
wire  _GEN24982 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24983 = io_x[27] ? _GEN21739 : _GEN24982;
wire  _GEN24984 = io_x[29] ? _GEN21743 : _GEN24983;
wire  _GEN24985 = io_x[75] ? _GEN24984 : _GEN21758;
wire  _GEN24986 = io_x[38] ? _GEN24985 : _GEN21871;
wire  _GEN24987 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN24988 = io_x[38] ? _GEN24987 : _GEN21833;
wire  _GEN24989 = io_x[34] ? _GEN24988 : _GEN24986;
wire  _GEN24990 = io_x[39] ? _GEN24989 : _GEN24981;
wire  _GEN24991 = io_x[46] ? _GEN24990 : _GEN24957;
wire  _GEN24992 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24993 = io_x[27] ? _GEN24992 : _GEN21739;
wire  _GEN24994 = io_x[29] ? _GEN24993 : _GEN21743;
wire  _GEN24995 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN24996 = io_x[75] ? _GEN24995 : _GEN24994;
wire  _GEN24997 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24998 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN24999 = io_x[27] ? _GEN24998 : _GEN24997;
wire  _GEN25000 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25001 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25002 = io_x[27] ? _GEN25001 : _GEN25000;
wire  _GEN25003 = io_x[29] ? _GEN25002 : _GEN24999;
wire  _GEN25004 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25005 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25006 = io_x[27] ? _GEN25005 : _GEN25004;
wire  _GEN25007 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25008 = io_x[29] ? _GEN25007 : _GEN25006;
wire  _GEN25009 = io_x[75] ? _GEN25008 : _GEN25003;
wire  _GEN25010 = io_x[38] ? _GEN25009 : _GEN24996;
wire  _GEN25011 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25012 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25013 = io_x[27] ? _GEN25012 : _GEN25011;
wire  _GEN25014 = io_x[29] ? _GEN25013 : _GEN21743;
wire  _GEN25015 = io_x[75] ? _GEN21772 : _GEN25014;
wire  _GEN25016 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25017 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25018 = io_x[27] ? _GEN25017 : _GEN25016;
wire  _GEN25019 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25020 = io_x[27] ? _GEN25019 : _GEN21739;
wire  _GEN25021 = io_x[29] ? _GEN25020 : _GEN25018;
wire  _GEN25022 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25023 = io_x[29] ? _GEN21743 : _GEN25022;
wire  _GEN25024 = io_x[75] ? _GEN25023 : _GEN25021;
wire  _GEN25025 = io_x[38] ? _GEN25024 : _GEN25015;
wire  _GEN25026 = io_x[34] ? _GEN25025 : _GEN25010;
wire  _GEN25027 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25028 = io_x[27] ? _GEN21750 : _GEN25027;
wire  _GEN25029 = io_x[29] ? _GEN21744 : _GEN25028;
wire  _GEN25030 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25031 = io_x[27] ? _GEN21750 : _GEN25030;
wire  _GEN25032 = io_x[29] ? _GEN21743 : _GEN25031;
wire  _GEN25033 = io_x[75] ? _GEN25032 : _GEN25029;
wire  _GEN25034 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25035 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25036 = io_x[27] ? _GEN25035 : _GEN25034;
wire  _GEN25037 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25038 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25039 = io_x[27] ? _GEN25038 : _GEN25037;
wire  _GEN25040 = io_x[29] ? _GEN25039 : _GEN25036;
wire  _GEN25041 = io_x[75] ? _GEN21772 : _GEN25040;
wire  _GEN25042 = io_x[38] ? _GEN25041 : _GEN25033;
wire  _GEN25043 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25044 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25045 = io_x[27] ? _GEN25044 : _GEN25043;
wire  _GEN25046 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25047 = io_x[27] ? _GEN21739 : _GEN25046;
wire  _GEN25048 = io_x[29] ? _GEN25047 : _GEN25045;
wire  _GEN25049 = io_x[75] ? _GEN21772 : _GEN25048;
wire  _GEN25050 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25051 = io_x[27] ? _GEN25050 : _GEN21739;
wire  _GEN25052 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25053 = io_x[27] ? _GEN25052 : _GEN21750;
wire  _GEN25054 = io_x[29] ? _GEN25053 : _GEN25051;
wire  _GEN25055 = io_x[75] ? _GEN21758 : _GEN25054;
wire  _GEN25056 = io_x[38] ? _GEN25055 : _GEN25049;
wire  _GEN25057 = io_x[34] ? _GEN25056 : _GEN25042;
wire  _GEN25058 = io_x[39] ? _GEN25057 : _GEN25026;
wire  _GEN25059 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25060 = io_x[27] ? _GEN21739 : _GEN25059;
wire  _GEN25061 = io_x[29] ? _GEN21744 : _GEN25060;
wire  _GEN25062 = io_x[75] ? _GEN25061 : _GEN21758;
wire  _GEN25063 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25064 = io_x[27] ? _GEN25063 : _GEN21739;
wire  _GEN25065 = io_x[29] ? _GEN21744 : _GEN25064;
wire  _GEN25066 = io_x[75] ? _GEN25065 : _GEN21758;
wire  _GEN25067 = io_x[38] ? _GEN25066 : _GEN25062;
wire  _GEN25068 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25069 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25070 = io_x[27] ? _GEN25069 : _GEN25068;
wire  _GEN25071 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25072 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25073 = io_x[27] ? _GEN25072 : _GEN25071;
wire  _GEN25074 = io_x[29] ? _GEN25073 : _GEN25070;
wire  _GEN25075 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25076 = io_x[29] ? _GEN25075 : _GEN21743;
wire  _GEN25077 = io_x[75] ? _GEN25076 : _GEN25074;
wire  _GEN25078 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25079 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25080 = io_x[27] ? _GEN25079 : _GEN25078;
wire  _GEN25081 = io_x[29] ? _GEN21743 : _GEN25080;
wire  _GEN25082 = io_x[75] ? _GEN25081 : _GEN21758;
wire  _GEN25083 = io_x[38] ? _GEN25082 : _GEN25077;
wire  _GEN25084 = io_x[34] ? _GEN25083 : _GEN25067;
wire  _GEN25085 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25086 = io_x[27] ? _GEN21750 : _GEN25085;
wire  _GEN25087 = io_x[29] ? _GEN21743 : _GEN25086;
wire  _GEN25088 = io_x[75] ? _GEN25087 : _GEN21758;
wire  _GEN25089 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25090 = io_x[27] ? _GEN25089 : _GEN21739;
wire  _GEN25091 = io_x[29] ? _GEN21743 : _GEN25090;
wire  _GEN25092 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25093 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25094 = io_x[27] ? _GEN25093 : _GEN21750;
wire  _GEN25095 = io_x[29] ? _GEN25094 : _GEN25092;
wire  _GEN25096 = io_x[75] ? _GEN25095 : _GEN25091;
wire  _GEN25097 = io_x[38] ? _GEN25096 : _GEN25088;
wire  _GEN25098 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25099 = io_x[27] ? _GEN21739 : _GEN25098;
wire  _GEN25100 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25101 = io_x[29] ? _GEN25100 : _GEN25099;
wire  _GEN25102 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25103 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25104 = io_x[27] ? _GEN25103 : _GEN25102;
wire  _GEN25105 = io_x[29] ? _GEN21743 : _GEN25104;
wire  _GEN25106 = io_x[75] ? _GEN25105 : _GEN25101;
wire  _GEN25107 = io_x[38] ? _GEN25106 : _GEN21833;
wire  _GEN25108 = io_x[34] ? _GEN25107 : _GEN25097;
wire  _GEN25109 = io_x[39] ? _GEN25108 : _GEN25084;
wire  _GEN25110 = io_x[46] ? _GEN25109 : _GEN25058;
wire  _GEN25111 = io_x[18] ? _GEN25110 : _GEN24991;
wire  _GEN25112 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25113 = io_x[27] ? _GEN25112 : _GEN21739;
wire  _GEN25114 = io_x[29] ? _GEN25113 : _GEN21743;
wire  _GEN25115 = io_x[75] ? _GEN21758 : _GEN25114;
wire  _GEN25116 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25117 = io_x[27] ? _GEN21750 : _GEN25116;
wire  _GEN25118 = io_x[29] ? _GEN25117 : _GEN21744;
wire  _GEN25119 = io_x[75] ? _GEN21758 : _GEN25118;
wire  _GEN25120 = io_x[38] ? _GEN25119 : _GEN25115;
wire  _GEN25121 = io_x[34] ? _GEN21927 : _GEN25120;
wire  _GEN25122 = io_x[39] ? _GEN21910 : _GEN25121;
wire  _GEN25123 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN25124 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN25125 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN25126 = io_x[38] ? _GEN25125 : _GEN25124;
wire  _GEN25127 = io_x[34] ? _GEN25126 : _GEN25123;
wire  _GEN25128 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN25129 = io_x[38] ? _GEN21833 : _GEN25128;
wire  _GEN25130 = io_x[34] ? _GEN25129 : _GEN21766;
wire  _GEN25131 = io_x[39] ? _GEN25130 : _GEN25127;
wire  _GEN25132 = io_x[46] ? _GEN25131 : _GEN25122;
wire  _GEN25133 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25134 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25135 = io_x[29] ? _GEN25134 : _GEN25133;
wire  _GEN25136 = io_x[75] ? _GEN21758 : _GEN25135;
wire  _GEN25137 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25138 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25139 = io_x[27] ? _GEN25138 : _GEN25137;
wire  _GEN25140 = io_x[29] ? _GEN21744 : _GEN25139;
wire  _GEN25141 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25142 = io_x[27] ? _GEN25141 : _GEN21739;
wire  _GEN25143 = io_x[29] ? _GEN25142 : _GEN21743;
wire  _GEN25144 = io_x[75] ? _GEN25143 : _GEN25140;
wire  _GEN25145 = io_x[38] ? _GEN25144 : _GEN25136;
wire  _GEN25146 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN25147 = io_x[75] ? _GEN25146 : _GEN21758;
wire  _GEN25148 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25149 = io_x[27] ? _GEN21739 : _GEN25148;
wire  _GEN25150 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25151 = io_x[27] ? _GEN25150 : _GEN21739;
wire  _GEN25152 = io_x[29] ? _GEN25151 : _GEN25149;
wire  _GEN25153 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25154 = io_x[27] ? _GEN21739 : _GEN25153;
wire  _GEN25155 = io_x[29] ? _GEN21743 : _GEN25154;
wire  _GEN25156 = io_x[75] ? _GEN25155 : _GEN25152;
wire  _GEN25157 = io_x[38] ? _GEN25156 : _GEN25147;
wire  _GEN25158 = io_x[34] ? _GEN25157 : _GEN25145;
wire  _GEN25159 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN25160 = io_x[38] ? _GEN21833 : _GEN25159;
wire  _GEN25161 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN25162 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25163 = io_x[29] ? _GEN21743 : _GEN25162;
wire  _GEN25164 = io_x[75] ? _GEN25163 : _GEN25161;
wire  _GEN25165 = io_x[38] ? _GEN21833 : _GEN25164;
wire  _GEN25166 = io_x[34] ? _GEN25165 : _GEN25160;
wire  _GEN25167 = io_x[39] ? _GEN25166 : _GEN25158;
wire  _GEN25168 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25169 = io_x[27] ? _GEN21739 : _GEN25168;
wire  _GEN25170 = io_x[29] ? _GEN21743 : _GEN25169;
wire  _GEN25171 = io_x[75] ? _GEN21758 : _GEN25170;
wire  _GEN25172 = io_x[38] ? _GEN21871 : _GEN25171;
wire  _GEN25173 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN25174 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25175 = io_x[29] ? _GEN21743 : _GEN25174;
wire  _GEN25176 = io_x[75] ? _GEN21758 : _GEN25175;
wire  _GEN25177 = io_x[38] ? _GEN25176 : _GEN25173;
wire  _GEN25178 = io_x[34] ? _GEN25177 : _GEN25172;
wire  _GEN25179 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25180 = io_x[27] ? _GEN21739 : _GEN25179;
wire  _GEN25181 = io_x[29] ? _GEN21743 : _GEN25180;
wire  _GEN25182 = io_x[75] ? _GEN21758 : _GEN25181;
wire  _GEN25183 = io_x[38] ? _GEN21871 : _GEN25182;
wire  _GEN25184 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25185 = io_x[27] ? _GEN21739 : _GEN25184;
wire  _GEN25186 = io_x[29] ? _GEN21744 : _GEN25185;
wire  _GEN25187 = io_x[75] ? _GEN25186 : _GEN21758;
wire  _GEN25188 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25189 = io_x[27] ? _GEN21739 : _GEN25188;
wire  _GEN25190 = io_x[29] ? _GEN21743 : _GEN25189;
wire  _GEN25191 = io_x[75] ? _GEN25190 : _GEN21758;
wire  _GEN25192 = io_x[38] ? _GEN25191 : _GEN25187;
wire  _GEN25193 = io_x[34] ? _GEN25192 : _GEN25183;
wire  _GEN25194 = io_x[39] ? _GEN25193 : _GEN25178;
wire  _GEN25195 = io_x[46] ? _GEN25194 : _GEN25167;
wire  _GEN25196 = io_x[18] ? _GEN25195 : _GEN25132;
wire  _GEN25197 = io_x[49] ? _GEN25196 : _GEN25111;
wire  _GEN25198 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25199 = io_x[27] ? _GEN25198 : _GEN21739;
wire  _GEN25200 = io_x[29] ? _GEN25199 : _GEN21743;
wire  _GEN25201 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25202 = io_x[27] ? _GEN25201 : _GEN21739;
wire  _GEN25203 = io_x[29] ? _GEN21743 : _GEN25202;
wire  _GEN25204 = io_x[75] ? _GEN25203 : _GEN25200;
wire  _GEN25205 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25206 = io_x[27] ? _GEN25205 : _GEN21739;
wire  _GEN25207 = io_x[29] ? _GEN25206 : _GEN21743;
wire  _GEN25208 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25209 = io_x[27] ? _GEN25208 : _GEN21739;
wire  _GEN25210 = io_x[29] ? _GEN25209 : _GEN21743;
wire  _GEN25211 = io_x[75] ? _GEN25210 : _GEN25207;
wire  _GEN25212 = io_x[38] ? _GEN25211 : _GEN25204;
wire  _GEN25213 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25214 = io_x[27] ? _GEN25213 : _GEN21739;
wire  _GEN25215 = io_x[29] ? _GEN25214 : _GEN21743;
wire  _GEN25216 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25217 = io_x[27] ? _GEN21739 : _GEN25216;
wire  _GEN25218 = io_x[29] ? _GEN25217 : _GEN21743;
wire  _GEN25219 = io_x[75] ? _GEN25218 : _GEN25215;
wire  _GEN25220 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25221 = io_x[27] ? _GEN25220 : _GEN21739;
wire  _GEN25222 = io_x[29] ? _GEN25221 : _GEN21744;
wire  _GEN25223 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25224 = io_x[27] ? _GEN25223 : _GEN21739;
wire  _GEN25225 = io_x[29] ? _GEN25224 : _GEN21743;
wire  _GEN25226 = io_x[75] ? _GEN25225 : _GEN25222;
wire  _GEN25227 = io_x[38] ? _GEN25226 : _GEN25219;
wire  _GEN25228 = io_x[34] ? _GEN25227 : _GEN25212;
wire  _GEN25229 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25230 = io_x[27] ? _GEN25229 : _GEN21750;
wire  _GEN25231 = io_x[29] ? _GEN25230 : _GEN21744;
wire  _GEN25232 = io_x[75] ? _GEN21758 : _GEN25231;
wire  _GEN25233 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25234 = io_x[27] ? _GEN25233 : _GEN21750;
wire  _GEN25235 = io_x[29] ? _GEN25234 : _GEN21744;
wire  _GEN25236 = io_x[75] ? _GEN21758 : _GEN25235;
wire  _GEN25237 = io_x[38] ? _GEN25236 : _GEN25232;
wire  _GEN25238 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25239 = io_x[27] ? _GEN25238 : _GEN21739;
wire  _GEN25240 = io_x[29] ? _GEN25239 : _GEN21743;
wire  _GEN25241 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25242 = io_x[27] ? _GEN25241 : _GEN21739;
wire  _GEN25243 = io_x[29] ? _GEN25242 : _GEN21743;
wire  _GEN25244 = io_x[75] ? _GEN25243 : _GEN25240;
wire  _GEN25245 = io_x[38] ? _GEN21871 : _GEN25244;
wire  _GEN25246 = io_x[34] ? _GEN25245 : _GEN25237;
wire  _GEN25247 = io_x[39] ? _GEN25246 : _GEN25228;
wire  _GEN25248 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN25249 = io_x[75] ? _GEN25248 : _GEN21758;
wire  _GEN25250 = io_x[38] ? _GEN21833 : _GEN25249;
wire  _GEN25251 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25252 = io_x[27] ? _GEN21739 : _GEN25251;
wire  _GEN25253 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25254 = io_x[27] ? _GEN21739 : _GEN25253;
wire  _GEN25255 = io_x[29] ? _GEN25254 : _GEN25252;
wire  _GEN25256 = io_x[75] ? _GEN21758 : _GEN25255;
wire  _GEN25257 = io_x[38] ? _GEN21833 : _GEN25256;
wire  _GEN25258 = io_x[34] ? _GEN25257 : _GEN25250;
wire  _GEN25259 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN25260 = io_x[34] ? _GEN25259 : _GEN21927;
wire  _GEN25261 = io_x[39] ? _GEN25260 : _GEN25258;
wire  _GEN25262 = io_x[46] ? _GEN25261 : _GEN25247;
wire  _GEN25263 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25264 = io_x[27] ? _GEN25263 : _GEN21750;
wire  _GEN25265 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25266 = io_x[27] ? _GEN25265 : _GEN21739;
wire  _GEN25267 = io_x[29] ? _GEN25266 : _GEN25264;
wire  _GEN25268 = io_x[75] ? _GEN21772 : _GEN25267;
wire  _GEN25269 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25270 = io_x[27] ? _GEN25269 : _GEN21739;
wire  _GEN25271 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25272 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25273 = io_x[27] ? _GEN25272 : _GEN25271;
wire  _GEN25274 = io_x[29] ? _GEN25273 : _GEN25270;
wire  _GEN25275 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25276 = io_x[27] ? _GEN25275 : _GEN21739;
wire  _GEN25277 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25278 = io_x[27] ? _GEN25277 : _GEN21739;
wire  _GEN25279 = io_x[29] ? _GEN25278 : _GEN25276;
wire  _GEN25280 = io_x[75] ? _GEN25279 : _GEN25274;
wire  _GEN25281 = io_x[38] ? _GEN25280 : _GEN25268;
wire  _GEN25282 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25283 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25284 = io_x[27] ? _GEN25283 : _GEN21739;
wire  _GEN25285 = io_x[29] ? _GEN25284 : _GEN25282;
wire  _GEN25286 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25287 = io_x[27] ? _GEN25286 : _GEN21750;
wire  _GEN25288 = io_x[29] ? _GEN25287 : _GEN21743;
wire  _GEN25289 = io_x[75] ? _GEN25288 : _GEN25285;
wire  _GEN25290 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25291 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25292 = io_x[27] ? _GEN25291 : _GEN25290;
wire  _GEN25293 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25294 = io_x[27] ? _GEN25293 : _GEN21739;
wire  _GEN25295 = io_x[29] ? _GEN25294 : _GEN25292;
wire  _GEN25296 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25297 = io_x[27] ? _GEN25296 : _GEN21739;
wire  _GEN25298 = io_x[29] ? _GEN25297 : _GEN21743;
wire  _GEN25299 = io_x[75] ? _GEN25298 : _GEN25295;
wire  _GEN25300 = io_x[38] ? _GEN25299 : _GEN25289;
wire  _GEN25301 = io_x[34] ? _GEN25300 : _GEN25281;
wire  _GEN25302 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25303 = io_x[27] ? _GEN25302 : _GEN21750;
wire  _GEN25304 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25305 = io_x[27] ? _GEN25304 : _GEN21750;
wire  _GEN25306 = io_x[29] ? _GEN25305 : _GEN25303;
wire  _GEN25307 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25308 = io_x[29] ? _GEN25307 : _GEN21743;
wire  _GEN25309 = io_x[75] ? _GEN25308 : _GEN25306;
wire  _GEN25310 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25311 = io_x[27] ? _GEN25310 : _GEN21750;
wire  _GEN25312 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25313 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25314 = io_x[27] ? _GEN25313 : _GEN25312;
wire  _GEN25315 = io_x[29] ? _GEN25314 : _GEN25311;
wire  _GEN25316 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25317 = io_x[27] ? _GEN25316 : _GEN21739;
wire  _GEN25318 = io_x[29] ? _GEN25317 : _GEN21744;
wire  _GEN25319 = io_x[75] ? _GEN25318 : _GEN25315;
wire  _GEN25320 = io_x[38] ? _GEN25319 : _GEN25309;
wire  _GEN25321 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25322 = io_x[27] ? _GEN21739 : _GEN25321;
wire  _GEN25323 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25324 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25325 = io_x[27] ? _GEN25324 : _GEN25323;
wire  _GEN25326 = io_x[29] ? _GEN25325 : _GEN25322;
wire  _GEN25327 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25328 = io_x[27] ? _GEN25327 : _GEN21739;
wire  _GEN25329 = io_x[29] ? _GEN25328 : _GEN21743;
wire  _GEN25330 = io_x[75] ? _GEN25329 : _GEN25326;
wire  _GEN25331 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25332 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25333 = io_x[27] ? _GEN25332 : _GEN21739;
wire  _GEN25334 = io_x[29] ? _GEN25333 : _GEN25331;
wire  _GEN25335 = io_x[75] ? _GEN21758 : _GEN25334;
wire  _GEN25336 = io_x[38] ? _GEN25335 : _GEN25330;
wire  _GEN25337 = io_x[34] ? _GEN25336 : _GEN25320;
wire  _GEN25338 = io_x[39] ? _GEN25337 : _GEN25301;
wire  _GEN25339 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25340 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25341 = io_x[27] ? _GEN25340 : _GEN25339;
wire  _GEN25342 = io_x[29] ? _GEN25341 : _GEN21743;
wire  _GEN25343 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25344 = io_x[27] ? _GEN21750 : _GEN25343;
wire  _GEN25345 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25346 = io_x[27] ? _GEN25345 : _GEN21750;
wire  _GEN25347 = io_x[29] ? _GEN25346 : _GEN25344;
wire  _GEN25348 = io_x[75] ? _GEN25347 : _GEN25342;
wire  _GEN25349 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25350 = io_x[27] ? _GEN21739 : _GEN25349;
wire  _GEN25351 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25352 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25353 = io_x[27] ? _GEN25352 : _GEN25351;
wire  _GEN25354 = io_x[29] ? _GEN25353 : _GEN25350;
wire  _GEN25355 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25356 = io_x[27] ? _GEN21739 : _GEN25355;
wire  _GEN25357 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25358 = io_x[27] ? _GEN25357 : _GEN21750;
wire  _GEN25359 = io_x[29] ? _GEN25358 : _GEN25356;
wire  _GEN25360 = io_x[75] ? _GEN25359 : _GEN25354;
wire  _GEN25361 = io_x[38] ? _GEN25360 : _GEN25348;
wire  _GEN25362 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25363 = io_x[27] ? _GEN21739 : _GEN25362;
wire  _GEN25364 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25365 = io_x[27] ? _GEN25364 : _GEN21750;
wire  _GEN25366 = io_x[29] ? _GEN25365 : _GEN25363;
wire  _GEN25367 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25368 = io_x[27] ? _GEN25367 : _GEN21739;
wire  _GEN25369 = io_x[29] ? _GEN25368 : _GEN21743;
wire  _GEN25370 = io_x[75] ? _GEN25369 : _GEN25366;
wire  _GEN25371 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25372 = io_x[27] ? _GEN25371 : _GEN21739;
wire  _GEN25373 = io_x[29] ? _GEN25372 : _GEN21743;
wire  _GEN25374 = io_x[75] ? _GEN21772 : _GEN25373;
wire  _GEN25375 = io_x[38] ? _GEN25374 : _GEN25370;
wire  _GEN25376 = io_x[34] ? _GEN25375 : _GEN25361;
wire  _GEN25377 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25378 = io_x[27] ? _GEN21739 : _GEN25377;
wire  _GEN25379 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25380 = io_x[27] ? _GEN25379 : _GEN21739;
wire  _GEN25381 = io_x[29] ? _GEN25380 : _GEN25378;
wire  _GEN25382 = io_x[75] ? _GEN25381 : _GEN21758;
wire  _GEN25383 = io_x[38] ? _GEN25382 : _GEN21833;
wire  _GEN25384 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN25385 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25386 = io_x[27] ? _GEN25385 : _GEN21739;
wire  _GEN25387 = io_x[29] ? _GEN25386 : _GEN21744;
wire  _GEN25388 = io_x[75] ? _GEN25387 : _GEN25384;
wire  _GEN25389 = io_x[38] ? _GEN25388 : _GEN21833;
wire  _GEN25390 = io_x[34] ? _GEN25389 : _GEN25383;
wire  _GEN25391 = io_x[39] ? _GEN25390 : _GEN25376;
wire  _GEN25392 = io_x[46] ? _GEN25391 : _GEN25338;
wire  _GEN25393 = io_x[18] ? _GEN25392 : _GEN25262;
wire  _GEN25394 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25395 = io_x[27] ? _GEN21739 : _GEN25394;
wire  _GEN25396 = io_x[29] ? _GEN25395 : _GEN21743;
wire  _GEN25397 = io_x[75] ? _GEN21758 : _GEN25396;
wire  _GEN25398 = io_x[38] ? _GEN25397 : _GEN21871;
wire  _GEN25399 = io_x[34] ? _GEN21766 : _GEN25398;
wire  _GEN25400 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN25401 = io_x[38] ? _GEN21871 : _GEN25400;
wire  _GEN25402 = io_x[34] ? _GEN21927 : _GEN25401;
wire  _GEN25403 = io_x[39] ? _GEN25402 : _GEN25399;
wire  _GEN25404 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN25405 = io_x[75] ? _GEN21772 : _GEN25404;
wire  _GEN25406 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN25407 = io_x[38] ? _GEN25406 : _GEN25405;
wire  _GEN25408 = io_x[34] ? _GEN25407 : _GEN21766;
wire  _GEN25409 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25410 = io_x[27] ? _GEN25409 : _GEN21750;
wire  _GEN25411 = io_x[29] ? _GEN25410 : _GEN21743;
wire  _GEN25412 = io_x[75] ? _GEN25411 : _GEN21758;
wire  _GEN25413 = io_x[38] ? _GEN21833 : _GEN25412;
wire  _GEN25414 = io_x[34] ? _GEN25413 : _GEN21766;
wire  _GEN25415 = io_x[39] ? _GEN25414 : _GEN25408;
wire  _GEN25416 = io_x[46] ? _GEN25415 : _GEN25403;
wire  _GEN25417 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25418 = io_x[27] ? _GEN21750 : _GEN25417;
wire  _GEN25419 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25420 = io_x[27] ? _GEN21750 : _GEN25419;
wire  _GEN25421 = io_x[29] ? _GEN25420 : _GEN25418;
wire  _GEN25422 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25423 = io_x[27] ? _GEN21750 : _GEN25422;
wire  _GEN25424 = io_x[29] ? _GEN25423 : _GEN21743;
wire  _GEN25425 = io_x[75] ? _GEN25424 : _GEN25421;
wire  _GEN25426 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25427 = io_x[27] ? _GEN21750 : _GEN25426;
wire  _GEN25428 = io_x[29] ? _GEN25427 : _GEN21744;
wire  _GEN25429 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25430 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25431 = io_x[27] ? _GEN25430 : _GEN25429;
wire  _GEN25432 = io_x[29] ? _GEN25431 : _GEN21743;
wire  _GEN25433 = io_x[75] ? _GEN25432 : _GEN25428;
wire  _GEN25434 = io_x[38] ? _GEN25433 : _GEN25425;
wire  _GEN25435 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25436 = io_x[27] ? _GEN25435 : _GEN21739;
wire  _GEN25437 = io_x[29] ? _GEN25436 : _GEN21743;
wire  _GEN25438 = io_x[75] ? _GEN25437 : _GEN21772;
wire  _GEN25439 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25440 = io_x[27] ? _GEN21739 : _GEN25439;
wire  _GEN25441 = io_x[29] ? _GEN25440 : _GEN21743;
wire  _GEN25442 = io_x[75] ? _GEN25441 : _GEN21772;
wire  _GEN25443 = io_x[38] ? _GEN25442 : _GEN25438;
wire  _GEN25444 = io_x[34] ? _GEN25443 : _GEN25434;
wire  _GEN25445 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25446 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25447 = io_x[27] ? _GEN25446 : _GEN25445;
wire  _GEN25448 = io_x[29] ? _GEN25447 : _GEN21744;
wire  _GEN25449 = io_x[75] ? _GEN21772 : _GEN25448;
wire  _GEN25450 = io_x[38] ? _GEN21833 : _GEN25449;
wire  _GEN25451 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25452 = io_x[27] ? _GEN21739 : _GEN25451;
wire  _GEN25453 = io_x[29] ? _GEN25452 : _GEN21743;
wire  _GEN25454 = io_x[75] ? _GEN21758 : _GEN25453;
wire  _GEN25455 = io_x[38] ? _GEN21871 : _GEN25454;
wire  _GEN25456 = io_x[34] ? _GEN25455 : _GEN25450;
wire  _GEN25457 = io_x[39] ? _GEN25456 : _GEN25444;
wire  _GEN25458 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN25459 = io_x[75] ? _GEN21758 : _GEN25458;
wire  _GEN25460 = io_x[38] ? _GEN21871 : _GEN25459;
wire  _GEN25461 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25462 = io_x[27] ? _GEN21739 : _GEN25461;
wire  _GEN25463 = io_x[29] ? _GEN21743 : _GEN25462;
wire  _GEN25464 = io_x[75] ? _GEN21758 : _GEN25463;
wire  _GEN25465 = io_x[38] ? _GEN25464 : _GEN21871;
wire  _GEN25466 = io_x[34] ? _GEN25465 : _GEN25460;
wire  _GEN25467 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25468 = io_x[29] ? _GEN25467 : _GEN21743;
wire  _GEN25469 = io_x[75] ? _GEN25468 : _GEN21758;
wire  _GEN25470 = io_x[38] ? _GEN21833 : _GEN25469;
wire  _GEN25471 = io_x[34] ? _GEN25470 : _GEN21927;
wire  _GEN25472 = io_x[39] ? _GEN25471 : _GEN25466;
wire  _GEN25473 = io_x[46] ? _GEN25472 : _GEN25457;
wire  _GEN25474 = io_x[18] ? _GEN25473 : _GEN25416;
wire  _GEN25475 = io_x[49] ? _GEN25474 : _GEN25393;
wire  _GEN25476 = io_x[24] ? _GEN25475 : _GEN25197;
wire  _GEN25477 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25478 = io_x[27] ? _GEN21750 : _GEN25477;
wire  _GEN25479 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25480 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25481 = io_x[27] ? _GEN25480 : _GEN25479;
wire  _GEN25482 = io_x[29] ? _GEN25481 : _GEN25478;
wire  _GEN25483 = io_x[75] ? _GEN25482 : _GEN21758;
wire  _GEN25484 = io_x[38] ? _GEN21871 : _GEN25483;
wire  _GEN25485 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN25486 = io_x[75] ? _GEN25485 : _GEN21758;
wire  _GEN25487 = io_x[38] ? _GEN21833 : _GEN25486;
wire  _GEN25488 = io_x[34] ? _GEN25487 : _GEN25484;
wire  _GEN25489 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25490 = io_x[29] ? _GEN21744 : _GEN25489;
wire  _GEN25491 = io_x[75] ? _GEN21758 : _GEN25490;
wire  _GEN25492 = io_x[38] ? _GEN21833 : _GEN25491;
wire  _GEN25493 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN25494 = io_x[38] ? _GEN21833 : _GEN25493;
wire  _GEN25495 = io_x[34] ? _GEN25494 : _GEN25492;
wire  _GEN25496 = io_x[39] ? _GEN25495 : _GEN25488;
wire  _GEN25497 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN25498 = io_x[34] ? _GEN21766 : _GEN25497;
wire  _GEN25499 = io_x[39] ? _GEN21910 : _GEN25498;
wire  _GEN25500 = io_x[46] ? _GEN25499 : _GEN25496;
wire  _GEN25501 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25502 = io_x[27] ? _GEN21750 : _GEN25501;
wire  _GEN25503 = io_x[29] ? _GEN21743 : _GEN25502;
wire  _GEN25504 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25505 = io_x[27] ? _GEN21739 : _GEN25504;
wire  _GEN25506 = io_x[29] ? _GEN21743 : _GEN25505;
wire  _GEN25507 = io_x[75] ? _GEN25506 : _GEN25503;
wire  _GEN25508 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25509 = io_x[27] ? _GEN21739 : _GEN25508;
wire  _GEN25510 = io_x[29] ? _GEN21744 : _GEN25509;
wire  _GEN25511 = io_x[75] ? _GEN21758 : _GEN25510;
wire  _GEN25512 = io_x[38] ? _GEN25511 : _GEN25507;
wire  _GEN25513 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN25514 = io_x[38] ? _GEN21871 : _GEN25513;
wire  _GEN25515 = io_x[34] ? _GEN25514 : _GEN25512;
wire  _GEN25516 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN25517 = io_x[75] ? _GEN25516 : _GEN21758;
wire  _GEN25518 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25519 = io_x[29] ? _GEN21743 : _GEN25518;
wire  _GEN25520 = io_x[75] ? _GEN21758 : _GEN25519;
wire  _GEN25521 = io_x[38] ? _GEN25520 : _GEN25517;
wire  _GEN25522 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25523 = io_x[27] ? _GEN21739 : _GEN25522;
wire  _GEN25524 = io_x[29] ? _GEN21743 : _GEN25523;
wire  _GEN25525 = io_x[75] ? _GEN21758 : _GEN25524;
wire  _GEN25526 = io_x[38] ? _GEN25525 : _GEN21833;
wire  _GEN25527 = io_x[34] ? _GEN25526 : _GEN25521;
wire  _GEN25528 = io_x[39] ? _GEN25527 : _GEN25515;
wire  _GEN25529 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN25530 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25531 = io_x[27] ? _GEN21750 : _GEN25530;
wire  _GEN25532 = io_x[29] ? _GEN21743 : _GEN25531;
wire  _GEN25533 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN25534 = io_x[75] ? _GEN25533 : _GEN25532;
wire  _GEN25535 = io_x[38] ? _GEN21871 : _GEN25534;
wire  _GEN25536 = io_x[34] ? _GEN25535 : _GEN25529;
wire  _GEN25537 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN25538 = io_x[75] ? _GEN21758 : _GEN25537;
wire  _GEN25539 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25540 = io_x[27] ? _GEN21750 : _GEN25539;
wire  _GEN25541 = io_x[29] ? _GEN21743 : _GEN25540;
wire  _GEN25542 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25543 = io_x[27] ? _GEN21739 : _GEN25542;
wire  _GEN25544 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25545 = io_x[27] ? _GEN25544 : _GEN21739;
wire  _GEN25546 = io_x[29] ? _GEN25545 : _GEN25543;
wire  _GEN25547 = io_x[75] ? _GEN25546 : _GEN25541;
wire  _GEN25548 = io_x[38] ? _GEN25547 : _GEN25538;
wire  _GEN25549 = io_x[34] ? _GEN25548 : _GEN21766;
wire  _GEN25550 = io_x[39] ? _GEN25549 : _GEN25536;
wire  _GEN25551 = io_x[46] ? _GEN25550 : _GEN25528;
wire  _GEN25552 = io_x[18] ? _GEN25551 : _GEN25500;
wire  _GEN25553 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25554 = io_x[29] ? _GEN21743 : _GEN25553;
wire  _GEN25555 = io_x[75] ? _GEN25554 : _GEN21758;
wire  _GEN25556 = io_x[38] ? _GEN25555 : _GEN21833;
wire  _GEN25557 = io_x[34] ? _GEN25556 : _GEN21927;
wire  _GEN25558 = io_x[39] ? _GEN22327 : _GEN25557;
wire  _GEN25559 = io_x[46] ? _GEN22145 : _GEN25558;
wire  _GEN25560 = io_x[18] ? _GEN25559 : _GEN23503;
wire  _GEN25561 = io_x[49] ? _GEN25560 : _GEN25552;
wire  _GEN25562 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25563 = io_x[27] ? _GEN25562 : _GEN21739;
wire  _GEN25564 = io_x[29] ? _GEN25563 : _GEN21743;
wire  _GEN25565 = io_x[75] ? _GEN21758 : _GEN25564;
wire  _GEN25566 = io_x[38] ? _GEN21871 : _GEN25565;
wire  _GEN25567 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25568 = io_x[27] ? _GEN25567 : _GEN21750;
wire  _GEN25569 = io_x[29] ? _GEN21744 : _GEN25568;
wire  _GEN25570 = io_x[75] ? _GEN25569 : _GEN21758;
wire  _GEN25571 = io_x[38] ? _GEN21871 : _GEN25570;
wire  _GEN25572 = io_x[34] ? _GEN25571 : _GEN25566;
wire  _GEN25573 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25574 = io_x[27] ? _GEN25573 : _GEN21739;
wire  _GEN25575 = io_x[29] ? _GEN25574 : _GEN21744;
wire  _GEN25576 = io_x[75] ? _GEN21758 : _GEN25575;
wire  _GEN25577 = io_x[38] ? _GEN21833 : _GEN25576;
wire  _GEN25578 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN25579 = io_x[34] ? _GEN25578 : _GEN25577;
wire  _GEN25580 = io_x[39] ? _GEN25579 : _GEN25572;
wire  _GEN25581 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN25582 = io_x[38] ? _GEN25581 : _GEN21833;
wire  _GEN25583 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25584 = io_x[27] ? _GEN25583 : _GEN21739;
wire  _GEN25585 = io_x[29] ? _GEN25584 : _GEN21743;
wire  _GEN25586 = io_x[75] ? _GEN21758 : _GEN25585;
wire  _GEN25587 = io_x[38] ? _GEN21871 : _GEN25586;
wire  _GEN25588 = io_x[34] ? _GEN25587 : _GEN25582;
wire  _GEN25589 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN25590 = io_x[75] ? _GEN25589 : _GEN21758;
wire  _GEN25591 = io_x[38] ? _GEN25590 : _GEN21833;
wire  _GEN25592 = io_x[34] ? _GEN25591 : _GEN21766;
wire  _GEN25593 = io_x[39] ? _GEN25592 : _GEN25588;
wire  _GEN25594 = io_x[46] ? _GEN25593 : _GEN25580;
wire  _GEN25595 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25596 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25597 = io_x[27] ? _GEN25596 : _GEN25595;
wire  _GEN25598 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25599 = io_x[27] ? _GEN25598 : _GEN21739;
wire  _GEN25600 = io_x[29] ? _GEN25599 : _GEN25597;
wire  _GEN25601 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25602 = io_x[27] ? _GEN21739 : _GEN25601;
wire  _GEN25603 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25604 = io_x[27] ? _GEN25603 : _GEN21739;
wire  _GEN25605 = io_x[29] ? _GEN25604 : _GEN25602;
wire  _GEN25606 = io_x[75] ? _GEN25605 : _GEN25600;
wire  _GEN25607 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25608 = io_x[27] ? _GEN25607 : _GEN21739;
wire  _GEN25609 = io_x[29] ? _GEN25608 : _GEN21743;
wire  _GEN25610 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25611 = io_x[27] ? _GEN21750 : _GEN25610;
wire  _GEN25612 = io_x[29] ? _GEN25611 : _GEN21744;
wire  _GEN25613 = io_x[75] ? _GEN25612 : _GEN25609;
wire  _GEN25614 = io_x[38] ? _GEN25613 : _GEN25606;
wire  _GEN25615 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25616 = io_x[27] ? _GEN21739 : _GEN25615;
wire  _GEN25617 = io_x[29] ? _GEN21744 : _GEN25616;
wire  _GEN25618 = io_x[75] ? _GEN25617 : _GEN21772;
wire  _GEN25619 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25620 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25621 = io_x[27] ? _GEN25620 : _GEN21739;
wire  _GEN25622 = io_x[29] ? _GEN25621 : _GEN25619;
wire  _GEN25623 = io_x[75] ? _GEN21758 : _GEN25622;
wire  _GEN25624 = io_x[38] ? _GEN25623 : _GEN25618;
wire  _GEN25625 = io_x[34] ? _GEN25624 : _GEN25614;
wire  _GEN25626 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25627 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25628 = io_x[27] ? _GEN25627 : _GEN25626;
wire  _GEN25629 = io_x[29] ? _GEN25628 : _GEN21743;
wire  _GEN25630 = io_x[75] ? _GEN25629 : _GEN21758;
wire  _GEN25631 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25632 = io_x[27] ? _GEN25631 : _GEN21739;
wire  _GEN25633 = io_x[29] ? _GEN25632 : _GEN21743;
wire  _GEN25634 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25635 = io_x[27] ? _GEN21739 : _GEN25634;
wire  _GEN25636 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25637 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25638 = io_x[27] ? _GEN25637 : _GEN25636;
wire  _GEN25639 = io_x[29] ? _GEN25638 : _GEN25635;
wire  _GEN25640 = io_x[75] ? _GEN25639 : _GEN25633;
wire  _GEN25641 = io_x[38] ? _GEN25640 : _GEN25630;
wire  _GEN25642 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN25643 = io_x[75] ? _GEN25642 : _GEN21758;
wire  _GEN25644 = io_x[38] ? _GEN21833 : _GEN25643;
wire  _GEN25645 = io_x[34] ? _GEN25644 : _GEN25641;
wire  _GEN25646 = io_x[39] ? _GEN25645 : _GEN25625;
wire  _GEN25647 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN25648 = io_x[38] ? _GEN25647 : _GEN21871;
wire  _GEN25649 = io_x[34] ? _GEN21927 : _GEN25648;
wire  _GEN25650 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25651 = io_x[27] ? _GEN21739 : _GEN25650;
wire  _GEN25652 = io_x[29] ? _GEN25651 : _GEN21743;
wire  _GEN25653 = io_x[75] ? _GEN21758 : _GEN25652;
wire  _GEN25654 = io_x[38] ? _GEN25653 : _GEN21833;
wire  _GEN25655 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25656 = io_x[27] ? _GEN25655 : _GEN21739;
wire  _GEN25657 = io_x[29] ? _GEN25656 : _GEN21743;
wire  _GEN25658 = io_x[75] ? _GEN25657 : _GEN21758;
wire  _GEN25659 = io_x[38] ? _GEN25658 : _GEN21833;
wire  _GEN25660 = io_x[34] ? _GEN25659 : _GEN25654;
wire  _GEN25661 = io_x[39] ? _GEN25660 : _GEN25649;
wire  _GEN25662 = io_x[46] ? _GEN25661 : _GEN25646;
wire  _GEN25663 = io_x[18] ? _GEN25662 : _GEN25594;
wire  _GEN25664 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN25665 = io_x[34] ? _GEN21927 : _GEN25664;
wire  _GEN25666 = io_x[39] ? _GEN21910 : _GEN25665;
wire  _GEN25667 = io_x[46] ? _GEN22145 : _GEN25666;
wire  _GEN25668 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN25669 = io_x[34] ? _GEN25668 : _GEN21927;
wire  _GEN25670 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN25671 = io_x[38] ? _GEN21871 : _GEN25670;
wire  _GEN25672 = io_x[34] ? _GEN21927 : _GEN25671;
wire  _GEN25673 = io_x[39] ? _GEN25672 : _GEN25669;
wire  _GEN25674 = io_x[46] ? _GEN22145 : _GEN25673;
wire  _GEN25675 = io_x[18] ? _GEN25674 : _GEN25667;
wire  _GEN25676 = io_x[49] ? _GEN25675 : _GEN25663;
wire  _GEN25677 = io_x[24] ? _GEN25676 : _GEN25561;
wire  _GEN25678 = io_x[80] ? _GEN25677 : _GEN25476;
wire  _GEN25679 = io_x[16] ? _GEN25678 : _GEN24923;
wire  _GEN25680 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25681 = io_x[27] ? _GEN21739 : _GEN25680;
wire  _GEN25682 = io_x[29] ? _GEN21743 : _GEN25681;
wire  _GEN25683 = io_x[75] ? _GEN21772 : _GEN25682;
wire  _GEN25684 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN25685 = io_x[38] ? _GEN25684 : _GEN25683;
wire  _GEN25686 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25687 = io_x[27] ? _GEN25686 : _GEN21739;
wire  _GEN25688 = io_x[29] ? _GEN25687 : _GEN21743;
wire  _GEN25689 = io_x[75] ? _GEN21758 : _GEN25688;
wire  _GEN25690 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25691 = io_x[27] ? _GEN25690 : _GEN21750;
wire  _GEN25692 = io_x[29] ? _GEN25691 : _GEN21744;
wire  _GEN25693 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN25694 = io_x[75] ? _GEN25693 : _GEN25692;
wire  _GEN25695 = io_x[38] ? _GEN25694 : _GEN25689;
wire  _GEN25696 = io_x[34] ? _GEN25695 : _GEN25685;
wire  _GEN25697 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25698 = io_x[27] ? _GEN25697 : _GEN21750;
wire  _GEN25699 = io_x[29] ? _GEN25698 : _GEN21744;
wire  _GEN25700 = io_x[75] ? _GEN21772 : _GEN25699;
wire  _GEN25701 = io_x[38] ? _GEN21871 : _GEN25700;
wire  _GEN25702 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25703 = io_x[27] ? _GEN21739 : _GEN25702;
wire  _GEN25704 = io_x[29] ? _GEN21743 : _GEN25703;
wire  _GEN25705 = io_x[75] ? _GEN21772 : _GEN25704;
wire  _GEN25706 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25707 = io_x[29] ? _GEN21743 : _GEN25706;
wire  _GEN25708 = io_x[75] ? _GEN21758 : _GEN25707;
wire  _GEN25709 = io_x[38] ? _GEN25708 : _GEN25705;
wire  _GEN25710 = io_x[34] ? _GEN25709 : _GEN25701;
wire  _GEN25711 = io_x[39] ? _GEN25710 : _GEN25696;
wire  _GEN25712 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25713 = io_x[27] ? _GEN21739 : _GEN25712;
wire  _GEN25714 = io_x[29] ? _GEN21743 : _GEN25713;
wire  _GEN25715 = io_x[75] ? _GEN21758 : _GEN25714;
wire  _GEN25716 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25717 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25718 = io_x[27] ? _GEN25717 : _GEN25716;
wire  _GEN25719 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25720 = io_x[27] ? _GEN21750 : _GEN25719;
wire  _GEN25721 = io_x[29] ? _GEN25720 : _GEN25718;
wire  _GEN25722 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25723 = io_x[27] ? _GEN25722 : _GEN21739;
wire  _GEN25724 = io_x[29] ? _GEN25723 : _GEN21743;
wire  _GEN25725 = io_x[75] ? _GEN25724 : _GEN25721;
wire  _GEN25726 = io_x[38] ? _GEN25725 : _GEN25715;
wire  _GEN25727 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25728 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25729 = io_x[27] ? _GEN25728 : _GEN25727;
wire  _GEN25730 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25731 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25732 = io_x[27] ? _GEN25731 : _GEN25730;
wire  _GEN25733 = io_x[29] ? _GEN25732 : _GEN25729;
wire  _GEN25734 = io_x[75] ? _GEN21758 : _GEN25733;
wire  _GEN25735 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25736 = io_x[27] ? _GEN21739 : _GEN25735;
wire  _GEN25737 = io_x[29] ? _GEN21743 : _GEN25736;
wire  _GEN25738 = io_x[75] ? _GEN21758 : _GEN25737;
wire  _GEN25739 = io_x[38] ? _GEN25738 : _GEN25734;
wire  _GEN25740 = io_x[34] ? _GEN25739 : _GEN25726;
wire  _GEN25741 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN25742 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN25743 = io_x[38] ? _GEN25742 : _GEN21833;
wire  _GEN25744 = io_x[34] ? _GEN25743 : _GEN25741;
wire  _GEN25745 = io_x[39] ? _GEN25744 : _GEN25740;
wire  _GEN25746 = io_x[46] ? _GEN25745 : _GEN25711;
wire  _GEN25747 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25748 = io_x[27] ? _GEN21739 : _GEN25747;
wire  _GEN25749 = io_x[29] ? _GEN21743 : _GEN25748;
wire  _GEN25750 = io_x[75] ? _GEN21772 : _GEN25749;
wire  _GEN25751 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25752 = io_x[27] ? _GEN21739 : _GEN25751;
wire  _GEN25753 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25754 = io_x[29] ? _GEN25753 : _GEN25752;
wire  _GEN25755 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25756 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25757 = io_x[27] ? _GEN25756 : _GEN25755;
wire  _GEN25758 = io_x[29] ? _GEN21743 : _GEN25757;
wire  _GEN25759 = io_x[75] ? _GEN25758 : _GEN25754;
wire  _GEN25760 = io_x[38] ? _GEN25759 : _GEN25750;
wire  _GEN25761 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN25762 = io_x[75] ? _GEN21772 : _GEN25761;
wire  _GEN25763 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25764 = io_x[27] ? _GEN25763 : _GEN21750;
wire  _GEN25765 = io_x[29] ? _GEN25764 : _GEN21744;
wire  _GEN25766 = io_x[75] ? _GEN21758 : _GEN25765;
wire  _GEN25767 = io_x[38] ? _GEN25766 : _GEN25762;
wire  _GEN25768 = io_x[34] ? _GEN25767 : _GEN25760;
wire  _GEN25769 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25770 = io_x[27] ? _GEN21750 : _GEN25769;
wire  _GEN25771 = io_x[29] ? _GEN25770 : _GEN21744;
wire  _GEN25772 = io_x[75] ? _GEN21758 : _GEN25771;
wire  _GEN25773 = io_x[38] ? _GEN21871 : _GEN25772;
wire  _GEN25774 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25775 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25776 = io_x[27] ? _GEN25775 : _GEN25774;
wire  _GEN25777 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25778 = io_x[27] ? _GEN25777 : _GEN21739;
wire  _GEN25779 = io_x[29] ? _GEN25778 : _GEN25776;
wire  _GEN25780 = io_x[75] ? _GEN21772 : _GEN25779;
wire  _GEN25781 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25782 = io_x[29] ? _GEN21743 : _GEN25781;
wire  _GEN25783 = io_x[75] ? _GEN21758 : _GEN25782;
wire  _GEN25784 = io_x[38] ? _GEN25783 : _GEN25780;
wire  _GEN25785 = io_x[34] ? _GEN25784 : _GEN25773;
wire  _GEN25786 = io_x[39] ? _GEN25785 : _GEN25768;
wire  _GEN25787 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25788 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25789 = io_x[27] ? _GEN25788 : _GEN25787;
wire  _GEN25790 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25791 = io_x[27] ? _GEN25790 : _GEN21739;
wire  _GEN25792 = io_x[29] ? _GEN25791 : _GEN25789;
wire  _GEN25793 = io_x[75] ? _GEN21758 : _GEN25792;
wire  _GEN25794 = io_x[38] ? _GEN25793 : _GEN21833;
wire  _GEN25795 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25796 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25797 = io_x[27] ? _GEN25796 : _GEN25795;
wire  _GEN25798 = io_x[29] ? _GEN21743 : _GEN25797;
wire  _GEN25799 = io_x[75] ? _GEN21758 : _GEN25798;
wire  _GEN25800 = io_x[38] ? _GEN21833 : _GEN25799;
wire  _GEN25801 = io_x[34] ? _GEN25800 : _GEN25794;
wire  _GEN25802 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25803 = io_x[27] ? _GEN21739 : _GEN25802;
wire  _GEN25804 = io_x[29] ? _GEN21743 : _GEN25803;
wire  _GEN25805 = io_x[75] ? _GEN21758 : _GEN25804;
wire  _GEN25806 = io_x[38] ? _GEN25805 : _GEN21871;
wire  _GEN25807 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25808 = io_x[29] ? _GEN25807 : _GEN21744;
wire  _GEN25809 = io_x[75] ? _GEN25808 : _GEN21758;
wire  _GEN25810 = io_x[38] ? _GEN25809 : _GEN21833;
wire  _GEN25811 = io_x[34] ? _GEN25810 : _GEN25806;
wire  _GEN25812 = io_x[39] ? _GEN25811 : _GEN25801;
wire  _GEN25813 = io_x[46] ? _GEN25812 : _GEN25786;
wire  _GEN25814 = io_x[18] ? _GEN25813 : _GEN25746;
wire  _GEN25815 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25816 = io_x[29] ? _GEN21744 : _GEN25815;
wire  _GEN25817 = io_x[75] ? _GEN21758 : _GEN25816;
wire  _GEN25818 = io_x[38] ? _GEN25817 : _GEN21833;
wire  _GEN25819 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25820 = io_x[29] ? _GEN21743 : _GEN25819;
wire  _GEN25821 = io_x[75] ? _GEN21758 : _GEN25820;
wire  _GEN25822 = io_x[38] ? _GEN25821 : _GEN21833;
wire  _GEN25823 = io_x[34] ? _GEN25822 : _GEN25818;
wire  _GEN25824 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN25825 = io_x[75] ? _GEN25824 : _GEN21772;
wire  _GEN25826 = io_x[38] ? _GEN21871 : _GEN25825;
wire  _GEN25827 = io_x[34] ? _GEN25826 : _GEN21927;
wire  _GEN25828 = io_x[39] ? _GEN25827 : _GEN25823;
wire  _GEN25829 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25830 = io_x[27] ? _GEN25829 : _GEN21739;
wire  _GEN25831 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25832 = io_x[29] ? _GEN25831 : _GEN25830;
wire  _GEN25833 = io_x[75] ? _GEN21758 : _GEN25832;
wire  _GEN25834 = io_x[38] ? _GEN21871 : _GEN25833;
wire  _GEN25835 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN25836 = io_x[38] ? _GEN25835 : _GEN21833;
wire  _GEN25837 = io_x[34] ? _GEN25836 : _GEN25834;
wire  _GEN25838 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25839 = io_x[27] ? _GEN25838 : _GEN21739;
wire  _GEN25840 = io_x[29] ? _GEN25839 : _GEN21743;
wire  _GEN25841 = io_x[75] ? _GEN25840 : _GEN21758;
wire  _GEN25842 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25843 = io_x[29] ? _GEN21743 : _GEN25842;
wire  _GEN25844 = io_x[75] ? _GEN25843 : _GEN21758;
wire  _GEN25845 = io_x[38] ? _GEN25844 : _GEN25841;
wire  _GEN25846 = io_x[34] ? _GEN25845 : _GEN21927;
wire  _GEN25847 = io_x[39] ? _GEN25846 : _GEN25837;
wire  _GEN25848 = io_x[46] ? _GEN25847 : _GEN25828;
wire  _GEN25849 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25850 = io_x[27] ? _GEN21739 : _GEN25849;
wire  _GEN25851 = io_x[29] ? _GEN21743 : _GEN25850;
wire  _GEN25852 = io_x[75] ? _GEN21758 : _GEN25851;
wire  _GEN25853 = io_x[38] ? _GEN25852 : _GEN21833;
wire  _GEN25854 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN25855 = io_x[75] ? _GEN25854 : _GEN21772;
wire  _GEN25856 = io_x[38] ? _GEN21871 : _GEN25855;
wire  _GEN25857 = io_x[34] ? _GEN25856 : _GEN25853;
wire  _GEN25858 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN25859 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25860 = io_x[27] ? _GEN25859 : _GEN21739;
wire  _GEN25861 = io_x[29] ? _GEN21744 : _GEN25860;
wire  _GEN25862 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25863 = io_x[27] ? _GEN25862 : _GEN21739;
wire  _GEN25864 = io_x[29] ? _GEN25863 : _GEN21743;
wire  _GEN25865 = io_x[75] ? _GEN25864 : _GEN25861;
wire  _GEN25866 = io_x[38] ? _GEN25865 : _GEN25858;
wire  _GEN25867 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25868 = io_x[27] ? _GEN25867 : _GEN21750;
wire  _GEN25869 = io_x[29] ? _GEN25868 : _GEN21744;
wire  _GEN25870 = io_x[75] ? _GEN25869 : _GEN21758;
wire  _GEN25871 = io_x[38] ? _GEN21833 : _GEN25870;
wire  _GEN25872 = io_x[34] ? _GEN25871 : _GEN25866;
wire  _GEN25873 = io_x[39] ? _GEN25872 : _GEN25857;
wire  _GEN25874 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25875 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25876 = io_x[27] ? _GEN25875 : _GEN25874;
wire  _GEN25877 = io_x[29] ? _GEN21743 : _GEN25876;
wire  _GEN25878 = io_x[75] ? _GEN21772 : _GEN25877;
wire  _GEN25879 = io_x[38] ? _GEN21871 : _GEN25878;
wire  _GEN25880 = io_x[34] ? _GEN21927 : _GEN25879;
wire  _GEN25881 = io_x[39] ? _GEN21910 : _GEN25880;
wire  _GEN25882 = io_x[46] ? _GEN25881 : _GEN25873;
wire  _GEN25883 = io_x[18] ? _GEN25882 : _GEN25848;
wire  _GEN25884 = io_x[49] ? _GEN25883 : _GEN25814;
wire  _GEN25885 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25886 = io_x[27] ? _GEN25885 : _GEN21739;
wire  _GEN25887 = io_x[29] ? _GEN25886 : _GEN21743;
wire  _GEN25888 = io_x[75] ? _GEN21772 : _GEN25887;
wire  _GEN25889 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25890 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25891 = io_x[27] ? _GEN25890 : _GEN25889;
wire  _GEN25892 = io_x[29] ? _GEN25891 : _GEN21743;
wire  _GEN25893 = io_x[75] ? _GEN21772 : _GEN25892;
wire  _GEN25894 = io_x[38] ? _GEN25893 : _GEN25888;
wire  _GEN25895 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25896 = io_x[27] ? _GEN25895 : _GEN21739;
wire  _GEN25897 = io_x[29] ? _GEN25896 : _GEN21743;
wire  _GEN25898 = io_x[75] ? _GEN21758 : _GEN25897;
wire  _GEN25899 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25900 = io_x[27] ? _GEN25899 : _GEN21750;
wire  _GEN25901 = io_x[29] ? _GEN25900 : _GEN21744;
wire  _GEN25902 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN25903 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25904 = io_x[27] ? _GEN25903 : _GEN21750;
wire  _GEN25905 = io_x[29] ? _GEN25904 : _GEN25902;
wire  _GEN25906 = io_x[75] ? _GEN25905 : _GEN25901;
wire  _GEN25907 = io_x[38] ? _GEN25906 : _GEN25898;
wire  _GEN25908 = io_x[34] ? _GEN25907 : _GEN25894;
wire  _GEN25909 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25910 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25911 = io_x[27] ? _GEN25910 : _GEN25909;
wire  _GEN25912 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25913 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25914 = io_x[27] ? _GEN25913 : _GEN25912;
wire  _GEN25915 = io_x[29] ? _GEN25914 : _GEN25911;
wire  _GEN25916 = io_x[75] ? _GEN21758 : _GEN25915;
wire  _GEN25917 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN25918 = io_x[29] ? _GEN21744 : _GEN25917;
wire  _GEN25919 = io_x[75] ? _GEN21758 : _GEN25918;
wire  _GEN25920 = io_x[38] ? _GEN25919 : _GEN25916;
wire  _GEN25921 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25922 = io_x[27] ? _GEN21750 : _GEN25921;
wire  _GEN25923 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25924 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25925 = io_x[27] ? _GEN25924 : _GEN25923;
wire  _GEN25926 = io_x[29] ? _GEN25925 : _GEN25922;
wire  _GEN25927 = io_x[75] ? _GEN21772 : _GEN25926;
wire  _GEN25928 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25929 = io_x[27] ? _GEN25928 : _GEN21739;
wire  _GEN25930 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25931 = io_x[27] ? _GEN25930 : _GEN21739;
wire  _GEN25932 = io_x[29] ? _GEN25931 : _GEN25929;
wire  _GEN25933 = io_x[75] ? _GEN21758 : _GEN25932;
wire  _GEN25934 = io_x[38] ? _GEN25933 : _GEN25927;
wire  _GEN25935 = io_x[34] ? _GEN25934 : _GEN25920;
wire  _GEN25936 = io_x[39] ? _GEN25935 : _GEN25908;
wire  _GEN25937 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25938 = io_x[27] ? _GEN25937 : _GEN21739;
wire  _GEN25939 = io_x[29] ? _GEN25938 : _GEN21743;
wire  _GEN25940 = io_x[75] ? _GEN25939 : _GEN21758;
wire  _GEN25941 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25942 = io_x[27] ? _GEN21739 : _GEN25941;
wire  _GEN25943 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25944 = io_x[27] ? _GEN21739 : _GEN25943;
wire  _GEN25945 = io_x[29] ? _GEN25944 : _GEN25942;
wire  _GEN25946 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25947 = io_x[27] ? _GEN21739 : _GEN25946;
wire  _GEN25948 = io_x[29] ? _GEN25947 : _GEN21743;
wire  _GEN25949 = io_x[75] ? _GEN25948 : _GEN25945;
wire  _GEN25950 = io_x[38] ? _GEN25949 : _GEN25940;
wire  _GEN25951 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25952 = io_x[27] ? _GEN21750 : _GEN25951;
wire  _GEN25953 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25954 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25955 = io_x[27] ? _GEN25954 : _GEN25953;
wire  _GEN25956 = io_x[29] ? _GEN25955 : _GEN25952;
wire  _GEN25957 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25958 = io_x[27] ? _GEN25957 : _GEN21739;
wire  _GEN25959 = io_x[29] ? _GEN25958 : _GEN21743;
wire  _GEN25960 = io_x[75] ? _GEN25959 : _GEN25956;
wire  _GEN25961 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25962 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25963 = io_x[27] ? _GEN25962 : _GEN25961;
wire  _GEN25964 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25965 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25966 = io_x[27] ? _GEN25965 : _GEN25964;
wire  _GEN25967 = io_x[29] ? _GEN25966 : _GEN25963;
wire  _GEN25968 = io_x[75] ? _GEN21758 : _GEN25967;
wire  _GEN25969 = io_x[38] ? _GEN25968 : _GEN25960;
wire  _GEN25970 = io_x[34] ? _GEN25969 : _GEN25950;
wire  _GEN25971 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25972 = io_x[27] ? _GEN25971 : _GEN21750;
wire  _GEN25973 = io_x[29] ? _GEN25972 : _GEN21743;
wire  _GEN25974 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN25975 = io_x[75] ? _GEN25974 : _GEN25973;
wire  _GEN25976 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25977 = io_x[27] ? _GEN25976 : _GEN21739;
wire  _GEN25978 = io_x[29] ? _GEN25977 : _GEN21743;
wire  _GEN25979 = io_x[75] ? _GEN25978 : _GEN21758;
wire  _GEN25980 = io_x[38] ? _GEN25979 : _GEN25975;
wire  _GEN25981 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN25982 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25983 = io_x[27] ? _GEN25982 : _GEN21739;
wire  _GEN25984 = io_x[29] ? _GEN25983 : _GEN21743;
wire  _GEN25985 = io_x[75] ? _GEN25984 : _GEN25981;
wire  _GEN25986 = io_x[38] ? _GEN25985 : _GEN21833;
wire  _GEN25987 = io_x[34] ? _GEN25986 : _GEN25980;
wire  _GEN25988 = io_x[39] ? _GEN25987 : _GEN25970;
wire  _GEN25989 = io_x[46] ? _GEN25988 : _GEN25936;
wire  _GEN25990 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25991 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25992 = io_x[27] ? _GEN25991 : _GEN25990;
wire  _GEN25993 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25994 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25995 = io_x[27] ? _GEN25994 : _GEN25993;
wire  _GEN25996 = io_x[29] ? _GEN25995 : _GEN25992;
wire  _GEN25997 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN25998 = io_x[27] ? _GEN21739 : _GEN25997;
wire  _GEN25999 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26000 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26001 = io_x[27] ? _GEN26000 : _GEN25999;
wire  _GEN26002 = io_x[29] ? _GEN26001 : _GEN25998;
wire  _GEN26003 = io_x[75] ? _GEN26002 : _GEN25996;
wire  _GEN26004 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26005 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26006 = io_x[27] ? _GEN26005 : _GEN26004;
wire  _GEN26007 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26008 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26009 = io_x[27] ? _GEN26008 : _GEN26007;
wire  _GEN26010 = io_x[29] ? _GEN26009 : _GEN26006;
wire  _GEN26011 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26012 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26013 = io_x[27] ? _GEN26012 : _GEN26011;
wire  _GEN26014 = io_x[29] ? _GEN26013 : _GEN21744;
wire  _GEN26015 = io_x[75] ? _GEN26014 : _GEN26010;
wire  _GEN26016 = io_x[38] ? _GEN26015 : _GEN26003;
wire  _GEN26017 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26018 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26019 = io_x[27] ? _GEN26018 : _GEN26017;
wire  _GEN26020 = io_x[29] ? _GEN26019 : _GEN21743;
wire  _GEN26021 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26022 = io_x[27] ? _GEN26021 : _GEN21739;
wire  _GEN26023 = io_x[29] ? _GEN26022 : _GEN21743;
wire  _GEN26024 = io_x[75] ? _GEN26023 : _GEN26020;
wire  _GEN26025 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26026 = io_x[27] ? _GEN26025 : _GEN21750;
wire  _GEN26027 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26028 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26029 = io_x[27] ? _GEN26028 : _GEN26027;
wire  _GEN26030 = io_x[29] ? _GEN26029 : _GEN26026;
wire  _GEN26031 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26032 = io_x[27] ? _GEN26031 : _GEN21739;
wire  _GEN26033 = io_x[29] ? _GEN26032 : _GEN21743;
wire  _GEN26034 = io_x[75] ? _GEN26033 : _GEN26030;
wire  _GEN26035 = io_x[38] ? _GEN26034 : _GEN26024;
wire  _GEN26036 = io_x[34] ? _GEN26035 : _GEN26016;
wire  _GEN26037 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26038 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26039 = io_x[27] ? _GEN26038 : _GEN26037;
wire  _GEN26040 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26041 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26042 = io_x[27] ? _GEN26041 : _GEN26040;
wire  _GEN26043 = io_x[29] ? _GEN26042 : _GEN26039;
wire  _GEN26044 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26045 = io_x[27] ? _GEN26044 : _GEN21750;
wire  _GEN26046 = io_x[29] ? _GEN26045 : _GEN21744;
wire  _GEN26047 = io_x[75] ? _GEN26046 : _GEN26043;
wire  _GEN26048 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26049 = io_x[27] ? _GEN21750 : _GEN26048;
wire  _GEN26050 = io_x[29] ? _GEN26049 : _GEN21744;
wire  _GEN26051 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26052 = io_x[27] ? _GEN26051 : _GEN21739;
wire  _GEN26053 = io_x[29] ? _GEN26052 : _GEN21743;
wire  _GEN26054 = io_x[75] ? _GEN26053 : _GEN26050;
wire  _GEN26055 = io_x[38] ? _GEN26054 : _GEN26047;
wire  _GEN26056 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26057 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26058 = io_x[27] ? _GEN26057 : _GEN26056;
wire  _GEN26059 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26060 = io_x[27] ? _GEN26059 : _GEN21739;
wire  _GEN26061 = io_x[29] ? _GEN26060 : _GEN26058;
wire  _GEN26062 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26063 = io_x[27] ? _GEN26062 : _GEN21750;
wire  _GEN26064 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26065 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26066 = io_x[27] ? _GEN26065 : _GEN26064;
wire  _GEN26067 = io_x[29] ? _GEN26066 : _GEN26063;
wire  _GEN26068 = io_x[75] ? _GEN26067 : _GEN26061;
wire  _GEN26069 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26070 = io_x[27] ? _GEN26069 : _GEN21739;
wire  _GEN26071 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26072 = io_x[27] ? _GEN26071 : _GEN21739;
wire  _GEN26073 = io_x[29] ? _GEN26072 : _GEN26070;
wire  _GEN26074 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26075 = io_x[27] ? _GEN26074 : _GEN21739;
wire  _GEN26076 = io_x[29] ? _GEN26075 : _GEN21743;
wire  _GEN26077 = io_x[75] ? _GEN26076 : _GEN26073;
wire  _GEN26078 = io_x[38] ? _GEN26077 : _GEN26068;
wire  _GEN26079 = io_x[34] ? _GEN26078 : _GEN26055;
wire  _GEN26080 = io_x[39] ? _GEN26079 : _GEN26036;
wire  _GEN26081 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26082 = io_x[27] ? _GEN26081 : _GEN21739;
wire  _GEN26083 = io_x[29] ? _GEN26082 : _GEN21743;
wire  _GEN26084 = io_x[75] ? _GEN26083 : _GEN21758;
wire  _GEN26085 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26086 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26087 = io_x[27] ? _GEN26086 : _GEN26085;
wire  _GEN26088 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26089 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26090 = io_x[27] ? _GEN26089 : _GEN26088;
wire  _GEN26091 = io_x[29] ? _GEN26090 : _GEN26087;
wire  _GEN26092 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26093 = io_x[27] ? _GEN26092 : _GEN21739;
wire  _GEN26094 = io_x[29] ? _GEN26093 : _GEN21743;
wire  _GEN26095 = io_x[75] ? _GEN26094 : _GEN26091;
wire  _GEN26096 = io_x[38] ? _GEN26095 : _GEN26084;
wire  _GEN26097 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26098 = io_x[27] ? _GEN21739 : _GEN26097;
wire  _GEN26099 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26100 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26101 = io_x[27] ? _GEN26100 : _GEN26099;
wire  _GEN26102 = io_x[29] ? _GEN26101 : _GEN26098;
wire  _GEN26103 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26104 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26105 = io_x[27] ? _GEN26104 : _GEN26103;
wire  _GEN26106 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26107 = io_x[27] ? _GEN26106 : _GEN21739;
wire  _GEN26108 = io_x[29] ? _GEN26107 : _GEN26105;
wire  _GEN26109 = io_x[75] ? _GEN26108 : _GEN26102;
wire  _GEN26110 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26111 = io_x[27] ? _GEN26110 : _GEN21739;
wire  _GEN26112 = io_x[29] ? _GEN26111 : _GEN21743;
wire  _GEN26113 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26114 = io_x[27] ? _GEN26113 : _GEN21739;
wire  _GEN26115 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26116 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26117 = io_x[27] ? _GEN26116 : _GEN26115;
wire  _GEN26118 = io_x[29] ? _GEN26117 : _GEN26114;
wire  _GEN26119 = io_x[75] ? _GEN26118 : _GEN26112;
wire  _GEN26120 = io_x[38] ? _GEN26119 : _GEN26109;
wire  _GEN26121 = io_x[34] ? _GEN26120 : _GEN26096;
wire  _GEN26122 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26123 = io_x[27] ? _GEN26122 : _GEN21739;
wire  _GEN26124 = io_x[29] ? _GEN26123 : _GEN21743;
wire  _GEN26125 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26126 = io_x[27] ? _GEN26125 : _GEN21750;
wire  _GEN26127 = io_x[29] ? _GEN26126 : _GEN21744;
wire  _GEN26128 = io_x[75] ? _GEN26127 : _GEN26124;
wire  _GEN26129 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26130 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26131 = io_x[27] ? _GEN26130 : _GEN26129;
wire  _GEN26132 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26133 = io_x[27] ? _GEN26132 : _GEN21739;
wire  _GEN26134 = io_x[29] ? _GEN26133 : _GEN26131;
wire  _GEN26135 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26136 = io_x[27] ? _GEN26135 : _GEN21739;
wire  _GEN26137 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26138 = io_x[27] ? _GEN26137 : _GEN21739;
wire  _GEN26139 = io_x[29] ? _GEN26138 : _GEN26136;
wire  _GEN26140 = io_x[75] ? _GEN26139 : _GEN26134;
wire  _GEN26141 = io_x[38] ? _GEN26140 : _GEN26128;
wire  _GEN26142 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26143 = io_x[27] ? _GEN26142 : _GEN21739;
wire  _GEN26144 = io_x[29] ? _GEN26143 : _GEN21743;
wire  _GEN26145 = io_x[75] ? _GEN21758 : _GEN26144;
wire  _GEN26146 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26147 = io_x[27] ? _GEN26146 : _GEN21739;
wire  _GEN26148 = io_x[29] ? _GEN26147 : _GEN21743;
wire  _GEN26149 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN26150 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26151 = io_x[27] ? _GEN26150 : _GEN21739;
wire  _GEN26152 = io_x[29] ? _GEN26151 : _GEN26149;
wire  _GEN26153 = io_x[75] ? _GEN26152 : _GEN26148;
wire  _GEN26154 = io_x[38] ? _GEN26153 : _GEN26145;
wire  _GEN26155 = io_x[34] ? _GEN26154 : _GEN26141;
wire  _GEN26156 = io_x[39] ? _GEN26155 : _GEN26121;
wire  _GEN26157 = io_x[46] ? _GEN26156 : _GEN26080;
wire  _GEN26158 = io_x[18] ? _GEN26157 : _GEN25989;
wire  _GEN26159 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26160 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26161 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26162 = io_x[27] ? _GEN26161 : _GEN26160;
wire  _GEN26163 = io_x[29] ? _GEN26162 : _GEN26159;
wire  _GEN26164 = io_x[75] ? _GEN21758 : _GEN26163;
wire  _GEN26165 = io_x[38] ? _GEN26164 : _GEN21833;
wire  _GEN26166 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN26167 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN26168 = io_x[38] ? _GEN26167 : _GEN26166;
wire  _GEN26169 = io_x[34] ? _GEN26168 : _GEN26165;
wire  _GEN26170 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26171 = io_x[27] ? _GEN26170 : _GEN21739;
wire  _GEN26172 = io_x[29] ? _GEN26171 : _GEN21743;
wire  _GEN26173 = io_x[75] ? _GEN26172 : _GEN21758;
wire  _GEN26174 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26175 = io_x[27] ? _GEN21750 : _GEN26174;
wire  _GEN26176 = io_x[29] ? _GEN21744 : _GEN26175;
wire  _GEN26177 = io_x[75] ? _GEN21758 : _GEN26176;
wire  _GEN26178 = io_x[38] ? _GEN26177 : _GEN26173;
wire  _GEN26179 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN26180 = io_x[75] ? _GEN26179 : _GEN21772;
wire  _GEN26181 = io_x[38] ? _GEN21871 : _GEN26180;
wire  _GEN26182 = io_x[34] ? _GEN26181 : _GEN26178;
wire  _GEN26183 = io_x[39] ? _GEN26182 : _GEN26169;
wire  _GEN26184 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26185 = io_x[27] ? _GEN21739 : _GEN26184;
wire  _GEN26186 = io_x[29] ? _GEN21743 : _GEN26185;
wire  _GEN26187 = io_x[75] ? _GEN21772 : _GEN26186;
wire  _GEN26188 = io_x[38] ? _GEN21871 : _GEN26187;
wire  _GEN26189 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN26190 = io_x[38] ? _GEN26189 : _GEN21833;
wire  _GEN26191 = io_x[34] ? _GEN26190 : _GEN26188;
wire  _GEN26192 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26193 = io_x[27] ? _GEN26192 : _GEN21739;
wire  _GEN26194 = io_x[29] ? _GEN26193 : _GEN21743;
wire  _GEN26195 = io_x[75] ? _GEN26194 : _GEN21758;
wire  _GEN26196 = io_x[38] ? _GEN26195 : _GEN21833;
wire  _GEN26197 = io_x[34] ? _GEN26196 : _GEN21927;
wire  _GEN26198 = io_x[39] ? _GEN26197 : _GEN26191;
wire  _GEN26199 = io_x[46] ? _GEN26198 : _GEN26183;
wire  _GEN26200 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26201 = io_x[27] ? _GEN26200 : _GEN21739;
wire  _GEN26202 = io_x[29] ? _GEN26201 : _GEN21743;
wire  _GEN26203 = io_x[75] ? _GEN21758 : _GEN26202;
wire  _GEN26204 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26205 = io_x[27] ? _GEN26204 : _GEN21750;
wire  _GEN26206 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26207 = io_x[27] ? _GEN26206 : _GEN21739;
wire  _GEN26208 = io_x[29] ? _GEN26207 : _GEN26205;
wire  _GEN26209 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26210 = io_x[27] ? _GEN26209 : _GEN21739;
wire  _GEN26211 = io_x[29] ? _GEN26210 : _GEN21743;
wire  _GEN26212 = io_x[75] ? _GEN26211 : _GEN26208;
wire  _GEN26213 = io_x[38] ? _GEN26212 : _GEN26203;
wire  _GEN26214 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26215 = io_x[27] ? _GEN21750 : _GEN26214;
wire  _GEN26216 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26217 = io_x[27] ? _GEN26216 : _GEN21750;
wire  _GEN26218 = io_x[29] ? _GEN26217 : _GEN26215;
wire  _GEN26219 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26220 = io_x[27] ? _GEN26219 : _GEN21739;
wire  _GEN26221 = io_x[29] ? _GEN26220 : _GEN21744;
wire  _GEN26222 = io_x[75] ? _GEN26221 : _GEN26218;
wire  _GEN26223 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26224 = io_x[27] ? _GEN21750 : _GEN26223;
wire  _GEN26225 = io_x[29] ? _GEN21744 : _GEN26224;
wire  _GEN26226 = io_x[75] ? _GEN26225 : _GEN21772;
wire  _GEN26227 = io_x[38] ? _GEN26226 : _GEN26222;
wire  _GEN26228 = io_x[34] ? _GEN26227 : _GEN26213;
wire  _GEN26229 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26230 = io_x[27] ? _GEN21750 : _GEN26229;
wire  _GEN26231 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26232 = io_x[27] ? _GEN26231 : _GEN21739;
wire  _GEN26233 = io_x[29] ? _GEN26232 : _GEN26230;
wire  _GEN26234 = io_x[75] ? _GEN26233 : _GEN21772;
wire  _GEN26235 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26236 = io_x[27] ? _GEN26235 : _GEN21750;
wire  _GEN26237 = io_x[29] ? _GEN26236 : _GEN21744;
wire  _GEN26238 = io_x[75] ? _GEN21758 : _GEN26237;
wire  _GEN26239 = io_x[38] ? _GEN26238 : _GEN26234;
wire  _GEN26240 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26241 = io_x[27] ? _GEN26240 : _GEN21739;
wire  _GEN26242 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN26243 = io_x[29] ? _GEN26242 : _GEN26241;
wire  _GEN26244 = io_x[75] ? _GEN26243 : _GEN21772;
wire  _GEN26245 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26246 = io_x[27] ? _GEN26245 : _GEN21739;
wire  _GEN26247 = io_x[29] ? _GEN26246 : _GEN21743;
wire  _GEN26248 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26249 = io_x[27] ? _GEN26248 : _GEN21739;
wire  _GEN26250 = io_x[29] ? _GEN26249 : _GEN21743;
wire  _GEN26251 = io_x[75] ? _GEN26250 : _GEN26247;
wire  _GEN26252 = io_x[38] ? _GEN26251 : _GEN26244;
wire  _GEN26253 = io_x[34] ? _GEN26252 : _GEN26239;
wire  _GEN26254 = io_x[39] ? _GEN26253 : _GEN26228;
wire  _GEN26255 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26256 = io_x[27] ? _GEN26255 : _GEN21739;
wire  _GEN26257 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26258 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26259 = io_x[27] ? _GEN26258 : _GEN26257;
wire  _GEN26260 = io_x[29] ? _GEN26259 : _GEN26256;
wire  _GEN26261 = io_x[75] ? _GEN21758 : _GEN26260;
wire  _GEN26262 = io_x[38] ? _GEN21871 : _GEN26261;
wire  _GEN26263 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN26264 = io_x[38] ? _GEN26263 : _GEN21833;
wire  _GEN26265 = io_x[34] ? _GEN26264 : _GEN26262;
wire  _GEN26266 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26267 = io_x[27] ? _GEN21750 : _GEN26266;
wire  _GEN26268 = io_x[29] ? _GEN21744 : _GEN26267;
wire  _GEN26269 = io_x[75] ? _GEN26268 : _GEN21758;
wire  _GEN26270 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26271 = io_x[27] ? _GEN26270 : _GEN21739;
wire  _GEN26272 = io_x[29] ? _GEN26271 : _GEN21743;
wire  _GEN26273 = io_x[75] ? _GEN26272 : _GEN21758;
wire  _GEN26274 = io_x[38] ? _GEN26273 : _GEN26269;
wire  _GEN26275 = io_x[34] ? _GEN26274 : _GEN21927;
wire  _GEN26276 = io_x[39] ? _GEN26275 : _GEN26265;
wire  _GEN26277 = io_x[46] ? _GEN26276 : _GEN26254;
wire  _GEN26278 = io_x[18] ? _GEN26277 : _GEN26199;
wire  _GEN26279 = io_x[49] ? _GEN26278 : _GEN26158;
wire  _GEN26280 = io_x[24] ? _GEN26279 : _GEN25884;
wire  _GEN26281 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26282 = io_x[27] ? _GEN26281 : _GEN21739;
wire  _GEN26283 = io_x[29] ? _GEN21743 : _GEN26282;
wire  _GEN26284 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26285 = io_x[27] ? _GEN21739 : _GEN26284;
wire  _GEN26286 = io_x[29] ? _GEN26285 : _GEN21743;
wire  _GEN26287 = io_x[75] ? _GEN26286 : _GEN26283;
wire  _GEN26288 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26289 = io_x[27] ? _GEN26288 : _GEN21739;
wire  _GEN26290 = io_x[29] ? _GEN21743 : _GEN26289;
wire  _GEN26291 = io_x[75] ? _GEN21758 : _GEN26290;
wire  _GEN26292 = io_x[38] ? _GEN26291 : _GEN26287;
wire  _GEN26293 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26294 = io_x[27] ? _GEN21750 : _GEN26293;
wire  _GEN26295 = io_x[29] ? _GEN21744 : _GEN26294;
wire  _GEN26296 = io_x[75] ? _GEN26295 : _GEN21758;
wire  _GEN26297 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26298 = io_x[27] ? _GEN26297 : _GEN21739;
wire  _GEN26299 = io_x[29] ? _GEN26298 : _GEN21743;
wire  _GEN26300 = io_x[75] ? _GEN21758 : _GEN26299;
wire  _GEN26301 = io_x[38] ? _GEN26300 : _GEN26296;
wire  _GEN26302 = io_x[34] ? _GEN26301 : _GEN26292;
wire  _GEN26303 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN26304 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26305 = io_x[29] ? _GEN26304 : _GEN26303;
wire  _GEN26306 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN26307 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26308 = io_x[27] ? _GEN21750 : _GEN26307;
wire  _GEN26309 = io_x[29] ? _GEN26308 : _GEN26306;
wire  _GEN26310 = io_x[75] ? _GEN26309 : _GEN26305;
wire  _GEN26311 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26312 = io_x[27] ? _GEN26311 : _GEN21739;
wire  _GEN26313 = io_x[29] ? _GEN21743 : _GEN26312;
wire  _GEN26314 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN26315 = io_x[29] ? _GEN26314 : _GEN21743;
wire  _GEN26316 = io_x[75] ? _GEN26315 : _GEN26313;
wire  _GEN26317 = io_x[38] ? _GEN26316 : _GEN26310;
wire  _GEN26318 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26319 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26320 = io_x[27] ? _GEN26319 : _GEN21739;
wire  _GEN26321 = io_x[29] ? _GEN26320 : _GEN26318;
wire  _GEN26322 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26323 = io_x[27] ? _GEN21739 : _GEN26322;
wire  _GEN26324 = io_x[29] ? _GEN26323 : _GEN21743;
wire  _GEN26325 = io_x[75] ? _GEN26324 : _GEN26321;
wire  _GEN26326 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN26327 = io_x[75] ? _GEN21758 : _GEN26326;
wire  _GEN26328 = io_x[38] ? _GEN26327 : _GEN26325;
wire  _GEN26329 = io_x[34] ? _GEN26328 : _GEN26317;
wire  _GEN26330 = io_x[39] ? _GEN26329 : _GEN26302;
wire  _GEN26331 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26332 = io_x[27] ? _GEN21739 : _GEN26331;
wire  _GEN26333 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26334 = io_x[27] ? _GEN26333 : _GEN21739;
wire  _GEN26335 = io_x[29] ? _GEN26334 : _GEN26332;
wire  _GEN26336 = io_x[75] ? _GEN21772 : _GEN26335;
wire  _GEN26337 = io_x[38] ? _GEN26336 : _GEN21833;
wire  _GEN26338 = io_x[34] ? _GEN21927 : _GEN26337;
wire  _GEN26339 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26340 = io_x[27] ? _GEN21739 : _GEN26339;
wire  _GEN26341 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26342 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26343 = io_x[27] ? _GEN26342 : _GEN26341;
wire  _GEN26344 = io_x[29] ? _GEN26343 : _GEN26340;
wire  _GEN26345 = io_x[75] ? _GEN21772 : _GEN26344;
wire  _GEN26346 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN26347 = io_x[29] ? _GEN26346 : _GEN21744;
wire  _GEN26348 = io_x[75] ? _GEN26347 : _GEN21772;
wire  _GEN26349 = io_x[38] ? _GEN26348 : _GEN26345;
wire  _GEN26350 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26351 = io_x[29] ? _GEN21743 : _GEN26350;
wire  _GEN26352 = io_x[75] ? _GEN21758 : _GEN26351;
wire  _GEN26353 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26354 = io_x[27] ? _GEN21739 : _GEN26353;
wire  _GEN26355 = io_x[29] ? _GEN26354 : _GEN21743;
wire  _GEN26356 = io_x[75] ? _GEN26355 : _GEN21758;
wire  _GEN26357 = io_x[38] ? _GEN26356 : _GEN26352;
wire  _GEN26358 = io_x[34] ? _GEN26357 : _GEN26349;
wire  _GEN26359 = io_x[39] ? _GEN26358 : _GEN26338;
wire  _GEN26360 = io_x[46] ? _GEN26359 : _GEN26330;
wire  _GEN26361 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26362 = io_x[27] ? _GEN21739 : _GEN26361;
wire  _GEN26363 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26364 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26365 = io_x[27] ? _GEN26364 : _GEN26363;
wire  _GEN26366 = io_x[29] ? _GEN26365 : _GEN26362;
wire  _GEN26367 = io_x[75] ? _GEN21772 : _GEN26366;
wire  _GEN26368 = io_x[38] ? _GEN21833 : _GEN26367;
wire  _GEN26369 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26370 = io_x[27] ? _GEN21739 : _GEN26369;
wire  _GEN26371 = io_x[29] ? _GEN21744 : _GEN26370;
wire  _GEN26372 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN26373 = io_x[75] ? _GEN26372 : _GEN26371;
wire  _GEN26374 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN26375 = io_x[29] ? _GEN26374 : _GEN21743;
wire  _GEN26376 = io_x[75] ? _GEN21758 : _GEN26375;
wire  _GEN26377 = io_x[38] ? _GEN26376 : _GEN26373;
wire  _GEN26378 = io_x[34] ? _GEN26377 : _GEN26368;
wire  _GEN26379 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN26380 = io_x[39] ? _GEN26379 : _GEN26378;
wire  _GEN26381 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26382 = io_x[27] ? _GEN21739 : _GEN26381;
wire  _GEN26383 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26384 = io_x[27] ? _GEN21739 : _GEN26383;
wire  _GEN26385 = io_x[29] ? _GEN26384 : _GEN26382;
wire  _GEN26386 = io_x[75] ? _GEN21758 : _GEN26385;
wire  _GEN26387 = io_x[38] ? _GEN26386 : _GEN21833;
wire  _GEN26388 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN26389 = io_x[34] ? _GEN26388 : _GEN26387;
wire  _GEN26390 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26391 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26392 = io_x[27] ? _GEN26391 : _GEN26390;
wire  _GEN26393 = io_x[29] ? _GEN26392 : _GEN21744;
wire  _GEN26394 = io_x[75] ? _GEN21758 : _GEN26393;
wire  _GEN26395 = io_x[38] ? _GEN21871 : _GEN26394;
wire  _GEN26396 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26397 = io_x[27] ? _GEN21739 : _GEN26396;
wire  _GEN26398 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26399 = io_x[27] ? _GEN21739 : _GEN26398;
wire  _GEN26400 = io_x[29] ? _GEN26399 : _GEN26397;
wire  _GEN26401 = io_x[75] ? _GEN21758 : _GEN26400;
wire  _GEN26402 = io_x[38] ? _GEN21833 : _GEN26401;
wire  _GEN26403 = io_x[34] ? _GEN26402 : _GEN26395;
wire  _GEN26404 = io_x[39] ? _GEN26403 : _GEN26389;
wire  _GEN26405 = io_x[46] ? _GEN26404 : _GEN26380;
wire  _GEN26406 = io_x[18] ? _GEN26405 : _GEN26360;
wire  _GEN26407 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN26408 = io_x[29] ? _GEN21744 : _GEN26407;
wire  _GEN26409 = io_x[75] ? _GEN26408 : _GEN21758;
wire  _GEN26410 = io_x[38] ? _GEN26409 : _GEN21833;
wire  _GEN26411 = io_x[34] ? _GEN26410 : _GEN21766;
wire  _GEN26412 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN26413 = io_x[34] ? _GEN26412 : _GEN21766;
wire  _GEN26414 = io_x[39] ? _GEN26413 : _GEN26411;
wire  _GEN26415 = io_x[46] ? _GEN22145 : _GEN26414;
wire  _GEN26416 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN26417 = io_x[39] ? _GEN22327 : _GEN26416;
wire  _GEN26418 = io_x[46] ? _GEN22145 : _GEN26417;
wire  _GEN26419 = io_x[18] ? _GEN26418 : _GEN26415;
wire  _GEN26420 = io_x[49] ? _GEN26419 : _GEN26406;
wire  _GEN26421 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN26422 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN26423 = io_x[29] ? _GEN26422 : _GEN21743;
wire  _GEN26424 = io_x[75] ? _GEN26423 : _GEN26421;
wire  _GEN26425 = io_x[38] ? _GEN21871 : _GEN26424;
wire  _GEN26426 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26427 = io_x[29] ? _GEN26426 : _GEN21743;
wire  _GEN26428 = io_x[75] ? _GEN21758 : _GEN26427;
wire  _GEN26429 = io_x[38] ? _GEN21833 : _GEN26428;
wire  _GEN26430 = io_x[34] ? _GEN26429 : _GEN26425;
wire  _GEN26431 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN26432 = io_x[75] ? _GEN26431 : _GEN21758;
wire  _GEN26433 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26434 = io_x[27] ? _GEN21739 : _GEN26433;
wire  _GEN26435 = io_x[29] ? _GEN26434 : _GEN21743;
wire  _GEN26436 = io_x[75] ? _GEN21758 : _GEN26435;
wire  _GEN26437 = io_x[38] ? _GEN26436 : _GEN26432;
wire  _GEN26438 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN26439 = io_x[34] ? _GEN26438 : _GEN26437;
wire  _GEN26440 = io_x[39] ? _GEN26439 : _GEN26430;
wire  _GEN26441 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26442 = io_x[27] ? _GEN21750 : _GEN26441;
wire  _GEN26443 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26444 = io_x[27] ? _GEN26443 : _GEN21750;
wire  _GEN26445 = io_x[29] ? _GEN26444 : _GEN26442;
wire  _GEN26446 = io_x[75] ? _GEN21758 : _GEN26445;
wire  _GEN26447 = io_x[38] ? _GEN26446 : _GEN21833;
wire  _GEN26448 = io_x[34] ? _GEN21927 : _GEN26447;
wire  _GEN26449 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26450 = io_x[27] ? _GEN21739 : _GEN26449;
wire  _GEN26451 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26452 = io_x[27] ? _GEN26451 : _GEN21750;
wire  _GEN26453 = io_x[29] ? _GEN26452 : _GEN26450;
wire  _GEN26454 = io_x[75] ? _GEN21758 : _GEN26453;
wire  _GEN26455 = io_x[38] ? _GEN21871 : _GEN26454;
wire  _GEN26456 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26457 = io_x[27] ? _GEN21739 : _GEN26456;
wire  _GEN26458 = io_x[29] ? _GEN21743 : _GEN26457;
wire  _GEN26459 = io_x[75] ? _GEN21758 : _GEN26458;
wire  _GEN26460 = io_x[38] ? _GEN21871 : _GEN26459;
wire  _GEN26461 = io_x[34] ? _GEN26460 : _GEN26455;
wire  _GEN26462 = io_x[39] ? _GEN26461 : _GEN26448;
wire  _GEN26463 = io_x[46] ? _GEN26462 : _GEN26440;
wire  _GEN26464 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26465 = io_x[27] ? _GEN26464 : _GEN21739;
wire  _GEN26466 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26467 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26468 = io_x[27] ? _GEN26467 : _GEN26466;
wire  _GEN26469 = io_x[29] ? _GEN26468 : _GEN26465;
wire  _GEN26470 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN26471 = io_x[29] ? _GEN26470 : _GEN21743;
wire  _GEN26472 = io_x[75] ? _GEN26471 : _GEN26469;
wire  _GEN26473 = io_x[38] ? _GEN21871 : _GEN26472;
wire  _GEN26474 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26475 = io_x[27] ? _GEN26474 : _GEN21739;
wire  _GEN26476 = io_x[29] ? _GEN26475 : _GEN21743;
wire  _GEN26477 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN26478 = io_x[75] ? _GEN26477 : _GEN26476;
wire  _GEN26479 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26480 = io_x[27] ? _GEN26479 : _GEN21739;
wire  _GEN26481 = io_x[29] ? _GEN26480 : _GEN21743;
wire  _GEN26482 = io_x[75] ? _GEN26481 : _GEN21758;
wire  _GEN26483 = io_x[38] ? _GEN26482 : _GEN26478;
wire  _GEN26484 = io_x[34] ? _GEN26483 : _GEN26473;
wire  _GEN26485 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26486 = io_x[27] ? _GEN26485 : _GEN21739;
wire  _GEN26487 = io_x[29] ? _GEN26486 : _GEN21743;
wire  _GEN26488 = io_x[75] ? _GEN21772 : _GEN26487;
wire  _GEN26489 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26490 = io_x[27] ? _GEN26489 : _GEN21739;
wire  _GEN26491 = io_x[29] ? _GEN26490 : _GEN21743;
wire  _GEN26492 = io_x[75] ? _GEN26491 : _GEN21758;
wire  _GEN26493 = io_x[38] ? _GEN26492 : _GEN26488;
wire  _GEN26494 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN26495 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26496 = io_x[27] ? _GEN26495 : _GEN21739;
wire  _GEN26497 = io_x[29] ? _GEN26496 : _GEN21743;
wire  _GEN26498 = io_x[75] ? _GEN21758 : _GEN26497;
wire  _GEN26499 = io_x[38] ? _GEN26498 : _GEN26494;
wire  _GEN26500 = io_x[34] ? _GEN26499 : _GEN26493;
wire  _GEN26501 = io_x[39] ? _GEN26500 : _GEN26484;
wire  _GEN26502 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26503 = io_x[27] ? _GEN21739 : _GEN26502;
wire  _GEN26504 = io_x[29] ? _GEN21743 : _GEN26503;
wire  _GEN26505 = io_x[75] ? _GEN26504 : _GEN21758;
wire  _GEN26506 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26507 = io_x[27] ? _GEN21739 : _GEN26506;
wire  _GEN26508 = io_x[29] ? _GEN21743 : _GEN26507;
wire  _GEN26509 = io_x[75] ? _GEN21758 : _GEN26508;
wire  _GEN26510 = io_x[38] ? _GEN26509 : _GEN26505;
wire  _GEN26511 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN26512 = io_x[34] ? _GEN26511 : _GEN26510;
wire  _GEN26513 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26514 = io_x[27] ? _GEN21750 : _GEN26513;
wire  _GEN26515 = io_x[29] ? _GEN21744 : _GEN26514;
wire  _GEN26516 = io_x[75] ? _GEN21758 : _GEN26515;
wire  _GEN26517 = io_x[38] ? _GEN21833 : _GEN26516;
wire  _GEN26518 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26519 = io_x[27] ? _GEN21739 : _GEN26518;
wire  _GEN26520 = io_x[29] ? _GEN21743 : _GEN26519;
wire  _GEN26521 = io_x[75] ? _GEN21758 : _GEN26520;
wire  _GEN26522 = io_x[38] ? _GEN21833 : _GEN26521;
wire  _GEN26523 = io_x[34] ? _GEN26522 : _GEN26517;
wire  _GEN26524 = io_x[39] ? _GEN26523 : _GEN26512;
wire  _GEN26525 = io_x[46] ? _GEN26524 : _GEN26501;
wire  _GEN26526 = io_x[18] ? _GEN26525 : _GEN26463;
wire  _GEN26527 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26528 = io_x[29] ? _GEN26527 : _GEN21743;
wire  _GEN26529 = io_x[75] ? _GEN26528 : _GEN21758;
wire  _GEN26530 = io_x[38] ? _GEN26529 : _GEN21833;
wire  _GEN26531 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26532 = io_x[29] ? _GEN26531 : _GEN21743;
wire  _GEN26533 = io_x[75] ? _GEN26532 : _GEN21758;
wire  _GEN26534 = io_x[38] ? _GEN21833 : _GEN26533;
wire  _GEN26535 = io_x[34] ? _GEN26534 : _GEN26530;
wire  _GEN26536 = io_x[39] ? _GEN26535 : _GEN21910;
wire  _GEN26537 = io_x[46] ? _GEN22145 : _GEN26536;
wire  _GEN26538 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN26539 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26540 = io_x[29] ? _GEN26539 : _GEN21743;
wire  _GEN26541 = io_x[75] ? _GEN26540 : _GEN21758;
wire  _GEN26542 = io_x[38] ? _GEN26541 : _GEN21833;
wire  _GEN26543 = io_x[34] ? _GEN26542 : _GEN26538;
wire  _GEN26544 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26545 = io_x[27] ? _GEN26544 : _GEN21750;
wire  _GEN26546 = io_x[29] ? _GEN26545 : _GEN21744;
wire  _GEN26547 = io_x[75] ? _GEN26546 : _GEN21758;
wire  _GEN26548 = io_x[38] ? _GEN26547 : _GEN21833;
wire  _GEN26549 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN26550 = io_x[75] ? _GEN21758 : _GEN26549;
wire  _GEN26551 = io_x[38] ? _GEN21833 : _GEN26550;
wire  _GEN26552 = io_x[34] ? _GEN26551 : _GEN26548;
wire  _GEN26553 = io_x[39] ? _GEN26552 : _GEN26543;
wire  _GEN26554 = io_x[46] ? _GEN22145 : _GEN26553;
wire  _GEN26555 = io_x[18] ? _GEN26554 : _GEN26537;
wire  _GEN26556 = io_x[49] ? _GEN26555 : _GEN26526;
wire  _GEN26557 = io_x[24] ? _GEN26556 : _GEN26420;
wire  _GEN26558 = io_x[80] ? _GEN26557 : _GEN26280;
wire  _GEN26559 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26560 = io_x[27] ? _GEN26559 : _GEN21739;
wire  _GEN26561 = io_x[29] ? _GEN26560 : _GEN21743;
wire  _GEN26562 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN26563 = io_x[75] ? _GEN26562 : _GEN26561;
wire  _GEN26564 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26565 = io_x[27] ? _GEN26564 : _GEN21739;
wire  _GEN26566 = io_x[29] ? _GEN26565 : _GEN21744;
wire  _GEN26567 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26568 = io_x[27] ? _GEN26567 : _GEN21739;
wire  _GEN26569 = io_x[29] ? _GEN26568 : _GEN21743;
wire  _GEN26570 = io_x[75] ? _GEN26569 : _GEN26566;
wire  _GEN26571 = io_x[38] ? _GEN26570 : _GEN26563;
wire  _GEN26572 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26573 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26574 = io_x[27] ? _GEN26573 : _GEN21739;
wire  _GEN26575 = io_x[29] ? _GEN26574 : _GEN26572;
wire  _GEN26576 = io_x[75] ? _GEN21772 : _GEN26575;
wire  _GEN26577 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26578 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26579 = io_x[27] ? _GEN26578 : _GEN26577;
wire  _GEN26580 = io_x[29] ? _GEN26579 : _GEN21744;
wire  _GEN26581 = io_x[75] ? _GEN21772 : _GEN26580;
wire  _GEN26582 = io_x[38] ? _GEN26581 : _GEN26576;
wire  _GEN26583 = io_x[34] ? _GEN26582 : _GEN26571;
wire  _GEN26584 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26585 = io_x[27] ? _GEN21750 : _GEN26584;
wire  _GEN26586 = io_x[29] ? _GEN21744 : _GEN26585;
wire  _GEN26587 = io_x[75] ? _GEN21772 : _GEN26586;
wire  _GEN26588 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26589 = io_x[27] ? _GEN21739 : _GEN26588;
wire  _GEN26590 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26591 = io_x[27] ? _GEN26590 : _GEN21739;
wire  _GEN26592 = io_x[29] ? _GEN26591 : _GEN26589;
wire  _GEN26593 = io_x[75] ? _GEN21758 : _GEN26592;
wire  _GEN26594 = io_x[38] ? _GEN26593 : _GEN26587;
wire  _GEN26595 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26596 = io_x[27] ? _GEN26595 : _GEN21739;
wire  _GEN26597 = io_x[29] ? _GEN26596 : _GEN21744;
wire  _GEN26598 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26599 = io_x[27] ? _GEN26598 : _GEN21739;
wire  _GEN26600 = io_x[29] ? _GEN26599 : _GEN21743;
wire  _GEN26601 = io_x[75] ? _GEN26600 : _GEN26597;
wire  _GEN26602 = io_x[38] ? _GEN21833 : _GEN26601;
wire  _GEN26603 = io_x[34] ? _GEN26602 : _GEN26594;
wire  _GEN26604 = io_x[39] ? _GEN26603 : _GEN26583;
wire  _GEN26605 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN26606 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26607 = io_x[27] ? _GEN21739 : _GEN26606;
wire  _GEN26608 = io_x[29] ? _GEN21743 : _GEN26607;
wire  _GEN26609 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26610 = io_x[27] ? _GEN21739 : _GEN26609;
wire  _GEN26611 = io_x[29] ? _GEN21743 : _GEN26610;
wire  _GEN26612 = io_x[75] ? _GEN26611 : _GEN26608;
wire  _GEN26613 = io_x[38] ? _GEN26612 : _GEN26605;
wire  _GEN26614 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26615 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26616 = io_x[27] ? _GEN26615 : _GEN26614;
wire  _GEN26617 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26618 = io_x[27] ? _GEN21739 : _GEN26617;
wire  _GEN26619 = io_x[29] ? _GEN26618 : _GEN26616;
wire  _GEN26620 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26621 = io_x[27] ? _GEN21739 : _GEN26620;
wire  _GEN26622 = io_x[29] ? _GEN21743 : _GEN26621;
wire  _GEN26623 = io_x[75] ? _GEN26622 : _GEN26619;
wire  _GEN26624 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26625 = io_x[27] ? _GEN21739 : _GEN26624;
wire  _GEN26626 = io_x[29] ? _GEN21744 : _GEN26625;
wire  _GEN26627 = io_x[75] ? _GEN26626 : _GEN21758;
wire  _GEN26628 = io_x[38] ? _GEN26627 : _GEN26623;
wire  _GEN26629 = io_x[34] ? _GEN26628 : _GEN26613;
wire  _GEN26630 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN26631 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26632 = io_x[27] ? _GEN21739 : _GEN26631;
wire  _GEN26633 = io_x[29] ? _GEN21743 : _GEN26632;
wire  _GEN26634 = io_x[75] ? _GEN26633 : _GEN21758;
wire  _GEN26635 = io_x[38] ? _GEN26634 : _GEN26630;
wire  _GEN26636 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26637 = io_x[27] ? _GEN21739 : _GEN26636;
wire  _GEN26638 = io_x[29] ? _GEN21743 : _GEN26637;
wire  _GEN26639 = io_x[75] ? _GEN26638 : _GEN21758;
wire  _GEN26640 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26641 = io_x[27] ? _GEN21750 : _GEN26640;
wire  _GEN26642 = io_x[29] ? _GEN21743 : _GEN26641;
wire  _GEN26643 = io_x[75] ? _GEN26642 : _GEN21758;
wire  _GEN26644 = io_x[38] ? _GEN26643 : _GEN26639;
wire  _GEN26645 = io_x[34] ? _GEN26644 : _GEN26635;
wire  _GEN26646 = io_x[39] ? _GEN26645 : _GEN26629;
wire  _GEN26647 = io_x[46] ? _GEN26646 : _GEN26604;
wire  _GEN26648 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26649 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26650 = io_x[27] ? _GEN26649 : _GEN26648;
wire  _GEN26651 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26652 = io_x[27] ? _GEN26651 : _GEN21739;
wire  _GEN26653 = io_x[29] ? _GEN26652 : _GEN26650;
wire  _GEN26654 = io_x[75] ? _GEN21772 : _GEN26653;
wire  _GEN26655 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26656 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26657 = io_x[27] ? _GEN26656 : _GEN26655;
wire  _GEN26658 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26659 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26660 = io_x[27] ? _GEN26659 : _GEN26658;
wire  _GEN26661 = io_x[29] ? _GEN26660 : _GEN26657;
wire  _GEN26662 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26663 = io_x[27] ? _GEN21739 : _GEN26662;
wire  _GEN26664 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26665 = io_x[27] ? _GEN26664 : _GEN21739;
wire  _GEN26666 = io_x[29] ? _GEN26665 : _GEN26663;
wire  _GEN26667 = io_x[75] ? _GEN26666 : _GEN26661;
wire  _GEN26668 = io_x[38] ? _GEN26667 : _GEN26654;
wire  _GEN26669 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26670 = io_x[27] ? _GEN26669 : _GEN21739;
wire  _GEN26671 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26672 = io_x[27] ? _GEN26671 : _GEN21739;
wire  _GEN26673 = io_x[29] ? _GEN26672 : _GEN26670;
wire  _GEN26674 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN26675 = io_x[75] ? _GEN26674 : _GEN26673;
wire  _GEN26676 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26677 = io_x[27] ? _GEN21739 : _GEN26676;
wire  _GEN26678 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26679 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26680 = io_x[27] ? _GEN26679 : _GEN26678;
wire  _GEN26681 = io_x[29] ? _GEN26680 : _GEN26677;
wire  _GEN26682 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26683 = io_x[27] ? _GEN26682 : _GEN21739;
wire  _GEN26684 = io_x[29] ? _GEN26683 : _GEN21743;
wire  _GEN26685 = io_x[75] ? _GEN26684 : _GEN26681;
wire  _GEN26686 = io_x[38] ? _GEN26685 : _GEN26675;
wire  _GEN26687 = io_x[34] ? _GEN26686 : _GEN26668;
wire  _GEN26688 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26689 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26690 = io_x[27] ? _GEN26689 : _GEN26688;
wire  _GEN26691 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26692 = io_x[27] ? _GEN26691 : _GEN21750;
wire  _GEN26693 = io_x[29] ? _GEN26692 : _GEN26690;
wire  _GEN26694 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26695 = io_x[27] ? _GEN21739 : _GEN26694;
wire  _GEN26696 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26697 = io_x[27] ? _GEN26696 : _GEN21739;
wire  _GEN26698 = io_x[29] ? _GEN26697 : _GEN26695;
wire  _GEN26699 = io_x[75] ? _GEN26698 : _GEN26693;
wire  _GEN26700 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26701 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26702 = io_x[27] ? _GEN26701 : _GEN26700;
wire  _GEN26703 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26704 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26705 = io_x[27] ? _GEN26704 : _GEN26703;
wire  _GEN26706 = io_x[29] ? _GEN26705 : _GEN26702;
wire  _GEN26707 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26708 = io_x[27] ? _GEN26707 : _GEN21739;
wire  _GEN26709 = io_x[29] ? _GEN26708 : _GEN21743;
wire  _GEN26710 = io_x[75] ? _GEN26709 : _GEN26706;
wire  _GEN26711 = io_x[38] ? _GEN26710 : _GEN26699;
wire  _GEN26712 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26713 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26714 = io_x[27] ? _GEN26713 : _GEN26712;
wire  _GEN26715 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26716 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26717 = io_x[27] ? _GEN26716 : _GEN26715;
wire  _GEN26718 = io_x[29] ? _GEN26717 : _GEN26714;
wire  _GEN26719 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26720 = io_x[27] ? _GEN26719 : _GEN21739;
wire  _GEN26721 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26722 = io_x[27] ? _GEN26721 : _GEN21739;
wire  _GEN26723 = io_x[29] ? _GEN26722 : _GEN26720;
wire  _GEN26724 = io_x[75] ? _GEN26723 : _GEN26718;
wire  _GEN26725 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN26726 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26727 = io_x[27] ? _GEN26726 : _GEN21739;
wire  _GEN26728 = io_x[29] ? _GEN26727 : _GEN21744;
wire  _GEN26729 = io_x[75] ? _GEN26728 : _GEN26725;
wire  _GEN26730 = io_x[38] ? _GEN26729 : _GEN26724;
wire  _GEN26731 = io_x[34] ? _GEN26730 : _GEN26711;
wire  _GEN26732 = io_x[39] ? _GEN26731 : _GEN26687;
wire  _GEN26733 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26734 = io_x[27] ? _GEN26733 : _GEN21739;
wire  _GEN26735 = io_x[29] ? _GEN26734 : _GEN21743;
wire  _GEN26736 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26737 = io_x[27] ? _GEN21750 : _GEN26736;
wire  _GEN26738 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26739 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26740 = io_x[27] ? _GEN26739 : _GEN26738;
wire  _GEN26741 = io_x[29] ? _GEN26740 : _GEN26737;
wire  _GEN26742 = io_x[75] ? _GEN26741 : _GEN26735;
wire  _GEN26743 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26744 = io_x[27] ? _GEN21739 : _GEN26743;
wire  _GEN26745 = io_x[29] ? _GEN21743 : _GEN26744;
wire  _GEN26746 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26747 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26748 = io_x[27] ? _GEN26747 : _GEN21750;
wire  _GEN26749 = io_x[29] ? _GEN26748 : _GEN26746;
wire  _GEN26750 = io_x[75] ? _GEN26749 : _GEN26745;
wire  _GEN26751 = io_x[38] ? _GEN26750 : _GEN26742;
wire  _GEN26752 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26753 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26754 = io_x[27] ? _GEN26753 : _GEN26752;
wire  _GEN26755 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26756 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26757 = io_x[27] ? _GEN26756 : _GEN26755;
wire  _GEN26758 = io_x[29] ? _GEN26757 : _GEN26754;
wire  _GEN26759 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26760 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26761 = io_x[27] ? _GEN26760 : _GEN26759;
wire  _GEN26762 = io_x[29] ? _GEN26761 : _GEN21743;
wire  _GEN26763 = io_x[75] ? _GEN26762 : _GEN26758;
wire  _GEN26764 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26765 = io_x[27] ? _GEN26764 : _GEN21739;
wire  _GEN26766 = io_x[29] ? _GEN26765 : _GEN21743;
wire  _GEN26767 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26768 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26769 = io_x[27] ? _GEN26768 : _GEN26767;
wire  _GEN26770 = io_x[29] ? _GEN26769 : _GEN21744;
wire  _GEN26771 = io_x[75] ? _GEN26770 : _GEN26766;
wire  _GEN26772 = io_x[38] ? _GEN26771 : _GEN26763;
wire  _GEN26773 = io_x[34] ? _GEN26772 : _GEN26751;
wire  _GEN26774 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN26775 = io_x[29] ? _GEN21744 : _GEN26774;
wire  _GEN26776 = io_x[75] ? _GEN26775 : _GEN21758;
wire  _GEN26777 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN26778 = io_x[29] ? _GEN26777 : _GEN21743;
wire  _GEN26779 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26780 = io_x[27] ? _GEN21739 : _GEN26779;
wire  _GEN26781 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26782 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26783 = io_x[27] ? _GEN26782 : _GEN26781;
wire  _GEN26784 = io_x[29] ? _GEN26783 : _GEN26780;
wire  _GEN26785 = io_x[75] ? _GEN26784 : _GEN26778;
wire  _GEN26786 = io_x[38] ? _GEN26785 : _GEN26776;
wire  _GEN26787 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26788 = io_x[27] ? _GEN26787 : _GEN21739;
wire  _GEN26789 = io_x[29] ? _GEN26788 : _GEN21743;
wire  _GEN26790 = io_x[75] ? _GEN21758 : _GEN26789;
wire  _GEN26791 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26792 = io_x[27] ? _GEN21739 : _GEN26791;
wire  _GEN26793 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26794 = io_x[27] ? _GEN26793 : _GEN21739;
wire  _GEN26795 = io_x[29] ? _GEN26794 : _GEN26792;
wire  _GEN26796 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26797 = io_x[27] ? _GEN21739 : _GEN26796;
wire  _GEN26798 = io_x[29] ? _GEN26797 : _GEN21744;
wire  _GEN26799 = io_x[75] ? _GEN26798 : _GEN26795;
wire  _GEN26800 = io_x[38] ? _GEN26799 : _GEN26790;
wire  _GEN26801 = io_x[34] ? _GEN26800 : _GEN26786;
wire  _GEN26802 = io_x[39] ? _GEN26801 : _GEN26773;
wire  _GEN26803 = io_x[46] ? _GEN26802 : _GEN26732;
wire  _GEN26804 = io_x[18] ? _GEN26803 : _GEN26647;
wire  _GEN26805 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN26806 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN26807 = io_x[38] ? _GEN26806 : _GEN26805;
wire  _GEN26808 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN26809 = io_x[38] ? _GEN21871 : _GEN26808;
wire  _GEN26810 = io_x[34] ? _GEN26809 : _GEN26807;
wire  _GEN26811 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN26812 = io_x[75] ? _GEN21758 : _GEN26811;
wire  _GEN26813 = io_x[38] ? _GEN21833 : _GEN26812;
wire  _GEN26814 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN26815 = io_x[38] ? _GEN21871 : _GEN26814;
wire  _GEN26816 = io_x[34] ? _GEN26815 : _GEN26813;
wire  _GEN26817 = io_x[39] ? _GEN26816 : _GEN26810;
wire  _GEN26818 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26819 = io_x[29] ? _GEN21743 : _GEN26818;
wire  _GEN26820 = io_x[75] ? _GEN26819 : _GEN21758;
wire  _GEN26821 = io_x[38] ? _GEN26820 : _GEN21871;
wire  _GEN26822 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN26823 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN26824 = io_x[38] ? _GEN26823 : _GEN26822;
wire  _GEN26825 = io_x[34] ? _GEN26824 : _GEN26821;
wire  _GEN26826 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN26827 = io_x[75] ? _GEN26826 : _GEN21758;
wire  _GEN26828 = io_x[38] ? _GEN21833 : _GEN26827;
wire  _GEN26829 = io_x[34] ? _GEN26828 : _GEN21927;
wire  _GEN26830 = io_x[39] ? _GEN26829 : _GEN26825;
wire  _GEN26831 = io_x[46] ? _GEN26830 : _GEN26817;
wire  _GEN26832 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26833 = io_x[29] ? _GEN21744 : _GEN26832;
wire  _GEN26834 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26835 = io_x[29] ? _GEN26834 : _GEN21744;
wire  _GEN26836 = io_x[75] ? _GEN26835 : _GEN26833;
wire  _GEN26837 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26838 = io_x[27] ? _GEN21750 : _GEN26837;
wire  _GEN26839 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26840 = io_x[27] ? _GEN26839 : _GEN21739;
wire  _GEN26841 = io_x[29] ? _GEN26840 : _GEN26838;
wire  _GEN26842 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26843 = io_x[27] ? _GEN21750 : _GEN26842;
wire  _GEN26844 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26845 = io_x[27] ? _GEN26844 : _GEN21750;
wire  _GEN26846 = io_x[29] ? _GEN26845 : _GEN26843;
wire  _GEN26847 = io_x[75] ? _GEN26846 : _GEN26841;
wire  _GEN26848 = io_x[38] ? _GEN26847 : _GEN26836;
wire  _GEN26849 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN26850 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26851 = io_x[27] ? _GEN21750 : _GEN26850;
wire  _GEN26852 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26853 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26854 = io_x[27] ? _GEN26853 : _GEN26852;
wire  _GEN26855 = io_x[29] ? _GEN26854 : _GEN26851;
wire  _GEN26856 = io_x[75] ? _GEN26855 : _GEN26849;
wire  _GEN26857 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26858 = io_x[27] ? _GEN26857 : _GEN21750;
wire  _GEN26859 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26860 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26861 = io_x[27] ? _GEN26860 : _GEN26859;
wire  _GEN26862 = io_x[29] ? _GEN26861 : _GEN26858;
wire  _GEN26863 = io_x[75] ? _GEN21772 : _GEN26862;
wire  _GEN26864 = io_x[38] ? _GEN26863 : _GEN26856;
wire  _GEN26865 = io_x[34] ? _GEN26864 : _GEN26848;
wire  _GEN26866 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26867 = io_x[27] ? _GEN26866 : _GEN21739;
wire  _GEN26868 = io_x[29] ? _GEN26867 : _GEN21743;
wire  _GEN26869 = io_x[75] ? _GEN21772 : _GEN26868;
wire  _GEN26870 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26871 = io_x[29] ? _GEN21743 : _GEN26870;
wire  _GEN26872 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26873 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26874 = io_x[27] ? _GEN26873 : _GEN21750;
wire  _GEN26875 = io_x[29] ? _GEN26874 : _GEN26872;
wire  _GEN26876 = io_x[75] ? _GEN26875 : _GEN26871;
wire  _GEN26877 = io_x[38] ? _GEN26876 : _GEN26869;
wire  _GEN26878 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26879 = io_x[27] ? _GEN26878 : _GEN21739;
wire  _GEN26880 = io_x[29] ? _GEN21743 : _GEN26879;
wire  _GEN26881 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26882 = io_x[27] ? _GEN26881 : _GEN21739;
wire  _GEN26883 = io_x[29] ? _GEN26882 : _GEN21744;
wire  _GEN26884 = io_x[75] ? _GEN26883 : _GEN26880;
wire  _GEN26885 = io_x[38] ? _GEN21833 : _GEN26884;
wire  _GEN26886 = io_x[34] ? _GEN26885 : _GEN26877;
wire  _GEN26887 = io_x[39] ? _GEN26886 : _GEN26865;
wire  _GEN26888 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26889 = io_x[27] ? _GEN21750 : _GEN26888;
wire  _GEN26890 = io_x[29] ? _GEN21744 : _GEN26889;
wire  _GEN26891 = io_x[75] ? _GEN21772 : _GEN26890;
wire  _GEN26892 = io_x[38] ? _GEN21871 : _GEN26891;
wire  _GEN26893 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN26894 = io_x[34] ? _GEN26893 : _GEN26892;
wire  _GEN26895 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26896 = io_x[27] ? _GEN21739 : _GEN26895;
wire  _GEN26897 = io_x[29] ? _GEN21743 : _GEN26896;
wire  _GEN26898 = io_x[75] ? _GEN26897 : _GEN21758;
wire  _GEN26899 = io_x[38] ? _GEN26898 : _GEN21833;
wire  _GEN26900 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26901 = io_x[29] ? _GEN26900 : _GEN21743;
wire  _GEN26902 = io_x[75] ? _GEN26901 : _GEN21758;
wire  _GEN26903 = io_x[38] ? _GEN21833 : _GEN26902;
wire  _GEN26904 = io_x[34] ? _GEN26903 : _GEN26899;
wire  _GEN26905 = io_x[39] ? _GEN26904 : _GEN26894;
wire  _GEN26906 = io_x[46] ? _GEN26905 : _GEN26887;
wire  _GEN26907 = io_x[18] ? _GEN26906 : _GEN26831;
wire  _GEN26908 = io_x[49] ? _GEN26907 : _GEN26804;
wire  _GEN26909 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26910 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26911 = io_x[27] ? _GEN26910 : _GEN26909;
wire  _GEN26912 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26913 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26914 = io_x[27] ? _GEN26913 : _GEN26912;
wire  _GEN26915 = io_x[29] ? _GEN26914 : _GEN26911;
wire  _GEN26916 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26917 = io_x[27] ? _GEN26916 : _GEN21739;
wire  _GEN26918 = io_x[29] ? _GEN26917 : _GEN21743;
wire  _GEN26919 = io_x[75] ? _GEN26918 : _GEN26915;
wire  _GEN26920 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26921 = io_x[27] ? _GEN26920 : _GEN21739;
wire  _GEN26922 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26923 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26924 = io_x[27] ? _GEN26923 : _GEN26922;
wire  _GEN26925 = io_x[29] ? _GEN26924 : _GEN26921;
wire  _GEN26926 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26927 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26928 = io_x[27] ? _GEN26927 : _GEN26926;
wire  _GEN26929 = io_x[29] ? _GEN26928 : _GEN21743;
wire  _GEN26930 = io_x[75] ? _GEN26929 : _GEN26925;
wire  _GEN26931 = io_x[38] ? _GEN26930 : _GEN26919;
wire  _GEN26932 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN26933 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26934 = io_x[27] ? _GEN26933 : _GEN21750;
wire  _GEN26935 = io_x[29] ? _GEN26934 : _GEN26932;
wire  _GEN26936 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26937 = io_x[27] ? _GEN26936 : _GEN21750;
wire  _GEN26938 = io_x[29] ? _GEN26937 : _GEN21743;
wire  _GEN26939 = io_x[75] ? _GEN26938 : _GEN26935;
wire  _GEN26940 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26941 = io_x[27] ? _GEN21739 : _GEN26940;
wire  _GEN26942 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26943 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26944 = io_x[27] ? _GEN26943 : _GEN26942;
wire  _GEN26945 = io_x[29] ? _GEN26944 : _GEN26941;
wire  _GEN26946 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26947 = io_x[27] ? _GEN26946 : _GEN21739;
wire  _GEN26948 = io_x[29] ? _GEN26947 : _GEN21743;
wire  _GEN26949 = io_x[75] ? _GEN26948 : _GEN26945;
wire  _GEN26950 = io_x[38] ? _GEN26949 : _GEN26939;
wire  _GEN26951 = io_x[34] ? _GEN26950 : _GEN26931;
wire  _GEN26952 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26953 = io_x[27] ? _GEN26952 : _GEN21739;
wire  _GEN26954 = io_x[29] ? _GEN26953 : _GEN21743;
wire  _GEN26955 = io_x[75] ? _GEN26954 : _GEN21772;
wire  _GEN26956 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26957 = io_x[27] ? _GEN26956 : _GEN21750;
wire  _GEN26958 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26959 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26960 = io_x[27] ? _GEN26959 : _GEN26958;
wire  _GEN26961 = io_x[29] ? _GEN26960 : _GEN26957;
wire  _GEN26962 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26963 = io_x[27] ? _GEN26962 : _GEN21739;
wire  _GEN26964 = io_x[29] ? _GEN26963 : _GEN21744;
wire  _GEN26965 = io_x[75] ? _GEN26964 : _GEN26961;
wire  _GEN26966 = io_x[38] ? _GEN26965 : _GEN26955;
wire  _GEN26967 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26968 = io_x[27] ? _GEN26967 : _GEN21739;
wire  _GEN26969 = io_x[29] ? _GEN26968 : _GEN21743;
wire  _GEN26970 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26971 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26972 = io_x[27] ? _GEN26971 : _GEN26970;
wire  _GEN26973 = io_x[29] ? _GEN26972 : _GEN21743;
wire  _GEN26974 = io_x[75] ? _GEN26973 : _GEN26969;
wire  _GEN26975 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26976 = io_x[27] ? _GEN26975 : _GEN21739;
wire  _GEN26977 = io_x[29] ? _GEN26976 : _GEN21744;
wire  _GEN26978 = io_x[75] ? _GEN21758 : _GEN26977;
wire  _GEN26979 = io_x[38] ? _GEN26978 : _GEN26974;
wire  _GEN26980 = io_x[34] ? _GEN26979 : _GEN26966;
wire  _GEN26981 = io_x[39] ? _GEN26980 : _GEN26951;
wire  _GEN26982 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26983 = io_x[27] ? _GEN26982 : _GEN21739;
wire  _GEN26984 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26985 = io_x[27] ? _GEN26984 : _GEN21750;
wire  _GEN26986 = io_x[29] ? _GEN26985 : _GEN26983;
wire  _GEN26987 = io_x[75] ? _GEN26986 : _GEN21758;
wire  _GEN26988 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26989 = io_x[27] ? _GEN21739 : _GEN26988;
wire  _GEN26990 = io_x[29] ? _GEN21743 : _GEN26989;
wire  _GEN26991 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26992 = io_x[27] ? _GEN26991 : _GEN21739;
wire  _GEN26993 = io_x[29] ? _GEN26992 : _GEN21743;
wire  _GEN26994 = io_x[75] ? _GEN26993 : _GEN26990;
wire  _GEN26995 = io_x[38] ? _GEN26994 : _GEN26987;
wire  _GEN26996 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26997 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN26998 = io_x[27] ? _GEN26997 : _GEN26996;
wire  _GEN26999 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27000 = io_x[27] ? _GEN26999 : _GEN21739;
wire  _GEN27001 = io_x[29] ? _GEN27000 : _GEN26998;
wire  _GEN27002 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN27003 = io_x[75] ? _GEN27002 : _GEN27001;
wire  _GEN27004 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27005 = io_x[27] ? _GEN27004 : _GEN21739;
wire  _GEN27006 = io_x[29] ? _GEN27005 : _GEN21743;
wire  _GEN27007 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN27008 = io_x[29] ? _GEN27007 : _GEN21743;
wire  _GEN27009 = io_x[75] ? _GEN27008 : _GEN27006;
wire  _GEN27010 = io_x[38] ? _GEN27009 : _GEN27003;
wire  _GEN27011 = io_x[34] ? _GEN27010 : _GEN26995;
wire  _GEN27012 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27013 = io_x[27] ? _GEN27012 : _GEN21750;
wire  _GEN27014 = io_x[29] ? _GEN27013 : _GEN21744;
wire  _GEN27015 = io_x[75] ? _GEN27014 : _GEN21758;
wire  _GEN27016 = io_x[38] ? _GEN27015 : _GEN21833;
wire  _GEN27017 = io_x[34] ? _GEN27016 : _GEN21927;
wire  _GEN27018 = io_x[39] ? _GEN27017 : _GEN27011;
wire  _GEN27019 = io_x[46] ? _GEN27018 : _GEN26981;
wire  _GEN27020 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27021 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27022 = io_x[27] ? _GEN27021 : _GEN27020;
wire  _GEN27023 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27024 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27025 = io_x[27] ? _GEN27024 : _GEN27023;
wire  _GEN27026 = io_x[29] ? _GEN27025 : _GEN27022;
wire  _GEN27027 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27028 = io_x[27] ? _GEN27027 : _GEN21750;
wire  _GEN27029 = io_x[29] ? _GEN27028 : _GEN21744;
wire  _GEN27030 = io_x[75] ? _GEN27029 : _GEN27026;
wire  _GEN27031 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27032 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27033 = io_x[27] ? _GEN27032 : _GEN27031;
wire  _GEN27034 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27035 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27036 = io_x[27] ? _GEN27035 : _GEN27034;
wire  _GEN27037 = io_x[29] ? _GEN27036 : _GEN27033;
wire  _GEN27038 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27039 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27040 = io_x[27] ? _GEN27039 : _GEN27038;
wire  _GEN27041 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27042 = io_x[27] ? _GEN27041 : _GEN21739;
wire  _GEN27043 = io_x[29] ? _GEN27042 : _GEN27040;
wire  _GEN27044 = io_x[75] ? _GEN27043 : _GEN27037;
wire  _GEN27045 = io_x[38] ? _GEN27044 : _GEN27030;
wire  _GEN27046 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27047 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27048 = io_x[27] ? _GEN27047 : _GEN27046;
wire  _GEN27049 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27050 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27051 = io_x[27] ? _GEN27050 : _GEN27049;
wire  _GEN27052 = io_x[29] ? _GEN27051 : _GEN27048;
wire  _GEN27053 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27054 = io_x[27] ? _GEN27053 : _GEN21750;
wire  _GEN27055 = io_x[29] ? _GEN27054 : _GEN21744;
wire  _GEN27056 = io_x[75] ? _GEN27055 : _GEN27052;
wire  _GEN27057 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27058 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27059 = io_x[27] ? _GEN27058 : _GEN27057;
wire  _GEN27060 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27061 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27062 = io_x[27] ? _GEN27061 : _GEN27060;
wire  _GEN27063 = io_x[29] ? _GEN27062 : _GEN27059;
wire  _GEN27064 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27065 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27066 = io_x[27] ? _GEN27065 : _GEN27064;
wire  _GEN27067 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27068 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27069 = io_x[27] ? _GEN27068 : _GEN27067;
wire  _GEN27070 = io_x[29] ? _GEN27069 : _GEN27066;
wire  _GEN27071 = io_x[75] ? _GEN27070 : _GEN27063;
wire  _GEN27072 = io_x[38] ? _GEN27071 : _GEN27056;
wire  _GEN27073 = io_x[34] ? _GEN27072 : _GEN27045;
wire  _GEN27074 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27075 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27076 = io_x[27] ? _GEN27075 : _GEN27074;
wire  _GEN27077 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27078 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27079 = io_x[27] ? _GEN27078 : _GEN27077;
wire  _GEN27080 = io_x[29] ? _GEN27079 : _GEN27076;
wire  _GEN27081 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27082 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27083 = io_x[27] ? _GEN27082 : _GEN27081;
wire  _GEN27084 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27085 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27086 = io_x[27] ? _GEN27085 : _GEN27084;
wire  _GEN27087 = io_x[29] ? _GEN27086 : _GEN27083;
wire  _GEN27088 = io_x[75] ? _GEN27087 : _GEN27080;
wire  _GEN27089 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27090 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27091 = io_x[27] ? _GEN27090 : _GEN27089;
wire  _GEN27092 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27093 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27094 = io_x[27] ? _GEN27093 : _GEN27092;
wire  _GEN27095 = io_x[29] ? _GEN27094 : _GEN27091;
wire  _GEN27096 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27097 = io_x[27] ? _GEN27096 : _GEN21750;
wire  _GEN27098 = io_x[29] ? _GEN27097 : _GEN21744;
wire  _GEN27099 = io_x[75] ? _GEN27098 : _GEN27095;
wire  _GEN27100 = io_x[38] ? _GEN27099 : _GEN27088;
wire  _GEN27101 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27102 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27103 = io_x[27] ? _GEN27102 : _GEN27101;
wire  _GEN27104 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27105 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27106 = io_x[27] ? _GEN27105 : _GEN27104;
wire  _GEN27107 = io_x[29] ? _GEN27106 : _GEN27103;
wire  _GEN27108 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27109 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27110 = io_x[27] ? _GEN27109 : _GEN27108;
wire  _GEN27111 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27112 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27113 = io_x[27] ? _GEN27112 : _GEN27111;
wire  _GEN27114 = io_x[29] ? _GEN27113 : _GEN27110;
wire  _GEN27115 = io_x[75] ? _GEN27114 : _GEN27107;
wire  _GEN27116 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27117 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27118 = io_x[27] ? _GEN27117 : _GEN27116;
wire  _GEN27119 = io_x[29] ? _GEN27118 : _GEN21743;
wire  _GEN27120 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27121 = io_x[27] ? _GEN27120 : _GEN21739;
wire  _GEN27122 = io_x[29] ? _GEN27121 : _GEN21743;
wire  _GEN27123 = io_x[75] ? _GEN27122 : _GEN27119;
wire  _GEN27124 = io_x[38] ? _GEN27123 : _GEN27115;
wire  _GEN27125 = io_x[34] ? _GEN27124 : _GEN27100;
wire  _GEN27126 = io_x[39] ? _GEN27125 : _GEN27073;
wire  _GEN27127 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27128 = io_x[27] ? _GEN27127 : _GEN21739;
wire  _GEN27129 = io_x[29] ? _GEN27128 : _GEN21743;
wire  _GEN27130 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27131 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27132 = io_x[27] ? _GEN27131 : _GEN27130;
wire  _GEN27133 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27134 = io_x[27] ? _GEN27133 : _GEN21750;
wire  _GEN27135 = io_x[29] ? _GEN27134 : _GEN27132;
wire  _GEN27136 = io_x[75] ? _GEN27135 : _GEN27129;
wire  _GEN27137 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27138 = io_x[27] ? _GEN27137 : _GEN21739;
wire  _GEN27139 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27140 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27141 = io_x[27] ? _GEN27140 : _GEN27139;
wire  _GEN27142 = io_x[29] ? _GEN27141 : _GEN27138;
wire  _GEN27143 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27144 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27145 = io_x[27] ? _GEN27144 : _GEN27143;
wire  _GEN27146 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27147 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27148 = io_x[27] ? _GEN27147 : _GEN27146;
wire  _GEN27149 = io_x[29] ? _GEN27148 : _GEN27145;
wire  _GEN27150 = io_x[75] ? _GEN27149 : _GEN27142;
wire  _GEN27151 = io_x[38] ? _GEN27150 : _GEN27136;
wire  _GEN27152 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN27153 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27154 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27155 = io_x[27] ? _GEN27154 : _GEN27153;
wire  _GEN27156 = io_x[29] ? _GEN27155 : _GEN27152;
wire  _GEN27157 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27158 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27159 = io_x[27] ? _GEN27158 : _GEN27157;
wire  _GEN27160 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27161 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27162 = io_x[27] ? _GEN27161 : _GEN27160;
wire  _GEN27163 = io_x[29] ? _GEN27162 : _GEN27159;
wire  _GEN27164 = io_x[75] ? _GEN27163 : _GEN27156;
wire  _GEN27165 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27166 = io_x[27] ? _GEN27165 : _GEN21739;
wire  _GEN27167 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27168 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27169 = io_x[27] ? _GEN27168 : _GEN27167;
wire  _GEN27170 = io_x[29] ? _GEN27169 : _GEN27166;
wire  _GEN27171 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27172 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27173 = io_x[27] ? _GEN27172 : _GEN27171;
wire  _GEN27174 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27175 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27176 = io_x[27] ? _GEN27175 : _GEN27174;
wire  _GEN27177 = io_x[29] ? _GEN27176 : _GEN27173;
wire  _GEN27178 = io_x[75] ? _GEN27177 : _GEN27170;
wire  _GEN27179 = io_x[38] ? _GEN27178 : _GEN27164;
wire  _GEN27180 = io_x[34] ? _GEN27179 : _GEN27151;
wire  _GEN27181 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27182 = io_x[27] ? _GEN21739 : _GEN27181;
wire  _GEN27183 = io_x[29] ? _GEN27182 : _GEN21743;
wire  _GEN27184 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27185 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27186 = io_x[27] ? _GEN27185 : _GEN27184;
wire  _GEN27187 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27188 = io_x[27] ? _GEN27187 : _GEN21739;
wire  _GEN27189 = io_x[29] ? _GEN27188 : _GEN27186;
wire  _GEN27190 = io_x[75] ? _GEN27189 : _GEN27183;
wire  _GEN27191 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27192 = io_x[27] ? _GEN21750 : _GEN27191;
wire  _GEN27193 = io_x[29] ? _GEN21744 : _GEN27192;
wire  _GEN27194 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27195 = io_x[27] ? _GEN27194 : _GEN21739;
wire  _GEN27196 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27197 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27198 = io_x[27] ? _GEN27197 : _GEN27196;
wire  _GEN27199 = io_x[29] ? _GEN27198 : _GEN27195;
wire  _GEN27200 = io_x[75] ? _GEN27199 : _GEN27193;
wire  _GEN27201 = io_x[38] ? _GEN27200 : _GEN27190;
wire  _GEN27202 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27203 = io_x[27] ? _GEN21739 : _GEN27202;
wire  _GEN27204 = io_x[29] ? _GEN27203 : _GEN21743;
wire  _GEN27205 = io_x[75] ? _GEN21758 : _GEN27204;
wire  _GEN27206 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27207 = io_x[27] ? _GEN21739 : _GEN27206;
wire  _GEN27208 = io_x[29] ? _GEN21743 : _GEN27207;
wire  _GEN27209 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27210 = io_x[27] ? _GEN21739 : _GEN27209;
wire  _GEN27211 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27212 = io_x[27] ? _GEN27211 : _GEN21739;
wire  _GEN27213 = io_x[29] ? _GEN27212 : _GEN27210;
wire  _GEN27214 = io_x[75] ? _GEN27213 : _GEN27208;
wire  _GEN27215 = io_x[38] ? _GEN27214 : _GEN27205;
wire  _GEN27216 = io_x[34] ? _GEN27215 : _GEN27201;
wire  _GEN27217 = io_x[39] ? _GEN27216 : _GEN27180;
wire  _GEN27218 = io_x[46] ? _GEN27217 : _GEN27126;
wire  _GEN27219 = io_x[18] ? _GEN27218 : _GEN27019;
wire  _GEN27220 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN27221 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27222 = io_x[27] ? _GEN21739 : _GEN27221;
wire  _GEN27223 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27224 = io_x[27] ? _GEN27223 : _GEN21739;
wire  _GEN27225 = io_x[29] ? _GEN27224 : _GEN27222;
wire  _GEN27226 = io_x[75] ? _GEN21772 : _GEN27225;
wire  _GEN27227 = io_x[38] ? _GEN27226 : _GEN27220;
wire  _GEN27228 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27229 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27230 = io_x[27] ? _GEN27229 : _GEN27228;
wire  _GEN27231 = io_x[29] ? _GEN27230 : _GEN21743;
wire  _GEN27232 = io_x[75] ? _GEN27231 : _GEN21772;
wire  _GEN27233 = io_x[38] ? _GEN21871 : _GEN27232;
wire  _GEN27234 = io_x[34] ? _GEN27233 : _GEN27227;
wire  _GEN27235 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27236 = io_x[27] ? _GEN27235 : _GEN21750;
wire  _GEN27237 = io_x[29] ? _GEN27236 : _GEN21744;
wire  _GEN27238 = io_x[75] ? _GEN27237 : _GEN21758;
wire  _GEN27239 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN27240 = io_x[29] ? _GEN27239 : _GEN21744;
wire  _GEN27241 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27242 = io_x[27] ? _GEN27241 : _GEN21750;
wire  _GEN27243 = io_x[29] ? _GEN27242 : _GEN21743;
wire  _GEN27244 = io_x[75] ? _GEN27243 : _GEN27240;
wire  _GEN27245 = io_x[38] ? _GEN27244 : _GEN27238;
wire  _GEN27246 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27247 = io_x[27] ? _GEN21739 : _GEN27246;
wire  _GEN27248 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27249 = io_x[27] ? _GEN27248 : _GEN21739;
wire  _GEN27250 = io_x[29] ? _GEN27249 : _GEN27247;
wire  _GEN27251 = io_x[75] ? _GEN21758 : _GEN27250;
wire  _GEN27252 = io_x[38] ? _GEN21833 : _GEN27251;
wire  _GEN27253 = io_x[34] ? _GEN27252 : _GEN27245;
wire  _GEN27254 = io_x[39] ? _GEN27253 : _GEN27234;
wire  _GEN27255 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN27256 = io_x[29] ? _GEN27255 : _GEN21744;
wire  _GEN27257 = io_x[75] ? _GEN27256 : _GEN21758;
wire  _GEN27258 = io_x[38] ? _GEN27257 : _GEN21871;
wire  _GEN27259 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN27260 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN27261 = io_x[38] ? _GEN27260 : _GEN27259;
wire  _GEN27262 = io_x[34] ? _GEN27261 : _GEN27258;
wire  _GEN27263 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN27264 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27265 = io_x[27] ? _GEN21750 : _GEN27264;
wire  _GEN27266 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27267 = io_x[29] ? _GEN27266 : _GEN27265;
wire  _GEN27268 = io_x[75] ? _GEN27267 : _GEN21758;
wire  _GEN27269 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN27270 = io_x[38] ? _GEN27269 : _GEN27268;
wire  _GEN27271 = io_x[34] ? _GEN27270 : _GEN27263;
wire  _GEN27272 = io_x[39] ? _GEN27271 : _GEN27262;
wire  _GEN27273 = io_x[46] ? _GEN27272 : _GEN27254;
wire  _GEN27274 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27275 = io_x[27] ? _GEN27274 : _GEN21750;
wire  _GEN27276 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27277 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27278 = io_x[27] ? _GEN27277 : _GEN27276;
wire  _GEN27279 = io_x[29] ? _GEN27278 : _GEN27275;
wire  _GEN27280 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27281 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27282 = io_x[27] ? _GEN27281 : _GEN27280;
wire  _GEN27283 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27284 = io_x[27] ? _GEN27283 : _GEN21739;
wire  _GEN27285 = io_x[29] ? _GEN27284 : _GEN27282;
wire  _GEN27286 = io_x[75] ? _GEN27285 : _GEN27279;
wire  _GEN27287 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27288 = io_x[27] ? _GEN27287 : _GEN21739;
wire  _GEN27289 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27290 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27291 = io_x[27] ? _GEN27290 : _GEN27289;
wire  _GEN27292 = io_x[29] ? _GEN27291 : _GEN27288;
wire  _GEN27293 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27294 = io_x[27] ? _GEN21750 : _GEN27293;
wire  _GEN27295 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27296 = io_x[27] ? _GEN27295 : _GEN21750;
wire  _GEN27297 = io_x[29] ? _GEN27296 : _GEN27294;
wire  _GEN27298 = io_x[75] ? _GEN27297 : _GEN27292;
wire  _GEN27299 = io_x[38] ? _GEN27298 : _GEN27286;
wire  _GEN27300 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27301 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27302 = io_x[27] ? _GEN27301 : _GEN21750;
wire  _GEN27303 = io_x[29] ? _GEN27302 : _GEN27300;
wire  _GEN27304 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27305 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27306 = io_x[27] ? _GEN27305 : _GEN27304;
wire  _GEN27307 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27308 = io_x[27] ? _GEN27307 : _GEN21739;
wire  _GEN27309 = io_x[29] ? _GEN27308 : _GEN27306;
wire  _GEN27310 = io_x[75] ? _GEN27309 : _GEN27303;
wire  _GEN27311 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27312 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27313 = io_x[27] ? _GEN27312 : _GEN27311;
wire  _GEN27314 = io_x[29] ? _GEN27313 : _GEN21744;
wire  _GEN27315 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27316 = io_x[27] ? _GEN27315 : _GEN21739;
wire  _GEN27317 = io_x[29] ? _GEN27316 : _GEN21743;
wire  _GEN27318 = io_x[75] ? _GEN27317 : _GEN27314;
wire  _GEN27319 = io_x[38] ? _GEN27318 : _GEN27310;
wire  _GEN27320 = io_x[34] ? _GEN27319 : _GEN27299;
wire  _GEN27321 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27322 = io_x[27] ? _GEN21750 : _GEN27321;
wire  _GEN27323 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27324 = io_x[27] ? _GEN27323 : _GEN21739;
wire  _GEN27325 = io_x[29] ? _GEN27324 : _GEN27322;
wire  _GEN27326 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27327 = io_x[27] ? _GEN21750 : _GEN27326;
wire  _GEN27328 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27329 = io_x[27] ? _GEN27328 : _GEN21750;
wire  _GEN27330 = io_x[29] ? _GEN27329 : _GEN27327;
wire  _GEN27331 = io_x[75] ? _GEN27330 : _GEN27325;
wire  _GEN27332 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27333 = io_x[27] ? _GEN27332 : _GEN21739;
wire  _GEN27334 = io_x[29] ? _GEN27333 : _GEN21743;
wire  _GEN27335 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN27336 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27337 = io_x[27] ? _GEN27336 : _GEN21739;
wire  _GEN27338 = io_x[29] ? _GEN27337 : _GEN27335;
wire  _GEN27339 = io_x[75] ? _GEN27338 : _GEN27334;
wire  _GEN27340 = io_x[38] ? _GEN27339 : _GEN27331;
wire  _GEN27341 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27342 = io_x[27] ? _GEN27341 : _GEN21739;
wire  _GEN27343 = io_x[29] ? _GEN27342 : _GEN21743;
wire  _GEN27344 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27345 = io_x[27] ? _GEN27344 : _GEN21739;
wire  _GEN27346 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27347 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27348 = io_x[27] ? _GEN27347 : _GEN27346;
wire  _GEN27349 = io_x[29] ? _GEN27348 : _GEN27345;
wire  _GEN27350 = io_x[75] ? _GEN27349 : _GEN27343;
wire  _GEN27351 = io_x[38] ? _GEN21871 : _GEN27350;
wire  _GEN27352 = io_x[34] ? _GEN27351 : _GEN27340;
wire  _GEN27353 = io_x[39] ? _GEN27352 : _GEN27320;
wire  _GEN27354 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27355 = io_x[27] ? _GEN27354 : _GEN21750;
wire  _GEN27356 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27357 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27358 = io_x[27] ? _GEN27357 : _GEN27356;
wire  _GEN27359 = io_x[29] ? _GEN27358 : _GEN27355;
wire  _GEN27360 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27361 = io_x[27] ? _GEN27360 : _GEN21739;
wire  _GEN27362 = io_x[29] ? _GEN27361 : _GEN21744;
wire  _GEN27363 = io_x[75] ? _GEN27362 : _GEN27359;
wire  _GEN27364 = io_x[38] ? _GEN21871 : _GEN27363;
wire  _GEN27365 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27366 = io_x[27] ? _GEN27365 : _GEN21750;
wire  _GEN27367 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27368 = io_x[27] ? _GEN27367 : _GEN21750;
wire  _GEN27369 = io_x[29] ? _GEN27368 : _GEN27366;
wire  _GEN27370 = io_x[75] ? _GEN27369 : _GEN21758;
wire  _GEN27371 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN27372 = io_x[38] ? _GEN27371 : _GEN27370;
wire  _GEN27373 = io_x[34] ? _GEN27372 : _GEN27364;
wire  _GEN27374 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27375 = io_x[29] ? _GEN27374 : _GEN21743;
wire  _GEN27376 = io_x[75] ? _GEN27375 : _GEN21758;
wire  _GEN27377 = io_x[38] ? _GEN27376 : _GEN21833;
wire  _GEN27378 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN27379 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27380 = io_x[27] ? _GEN27379 : _GEN21739;
wire  _GEN27381 = io_x[29] ? _GEN27380 : _GEN27378;
wire  _GEN27382 = io_x[75] ? _GEN27381 : _GEN21758;
wire  _GEN27383 = io_x[38] ? _GEN21833 : _GEN27382;
wire  _GEN27384 = io_x[34] ? _GEN27383 : _GEN27377;
wire  _GEN27385 = io_x[39] ? _GEN27384 : _GEN27373;
wire  _GEN27386 = io_x[46] ? _GEN27385 : _GEN27353;
wire  _GEN27387 = io_x[18] ? _GEN27386 : _GEN27273;
wire  _GEN27388 = io_x[49] ? _GEN27387 : _GEN27219;
wire  _GEN27389 = io_x[24] ? _GEN27388 : _GEN26908;
wire  _GEN27390 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN27391 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27392 = io_x[27] ? _GEN21739 : _GEN27391;
wire  _GEN27393 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27394 = io_x[27] ? _GEN27393 : _GEN21739;
wire  _GEN27395 = io_x[29] ? _GEN27394 : _GEN27392;
wire  _GEN27396 = io_x[75] ? _GEN27395 : _GEN27390;
wire  _GEN27397 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27398 = io_x[27] ? _GEN27397 : _GEN21739;
wire  _GEN27399 = io_x[29] ? _GEN27398 : _GEN21743;
wire  _GEN27400 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27401 = io_x[29] ? _GEN21743 : _GEN27400;
wire  _GEN27402 = io_x[75] ? _GEN27401 : _GEN27399;
wire  _GEN27403 = io_x[38] ? _GEN27402 : _GEN27396;
wire  _GEN27404 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27405 = io_x[27] ? _GEN21750 : _GEN27404;
wire  _GEN27406 = io_x[29] ? _GEN21744 : _GEN27405;
wire  _GEN27407 = io_x[75] ? _GEN27406 : _GEN21772;
wire  _GEN27408 = io_x[38] ? _GEN21871 : _GEN27407;
wire  _GEN27409 = io_x[34] ? _GEN27408 : _GEN27403;
wire  _GEN27410 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27411 = io_x[27] ? _GEN27410 : _GEN21750;
wire  _GEN27412 = io_x[29] ? _GEN27411 : _GEN21744;
wire  _GEN27413 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27414 = io_x[27] ? _GEN21739 : _GEN27413;
wire  _GEN27415 = io_x[29] ? _GEN27414 : _GEN21743;
wire  _GEN27416 = io_x[75] ? _GEN27415 : _GEN27412;
wire  _GEN27417 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27418 = io_x[27] ? _GEN27417 : _GEN21739;
wire  _GEN27419 = io_x[29] ? _GEN27418 : _GEN21743;
wire  _GEN27420 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27421 = io_x[27] ? _GEN27420 : _GEN21750;
wire  _GEN27422 = io_x[29] ? _GEN27421 : _GEN21743;
wire  _GEN27423 = io_x[75] ? _GEN27422 : _GEN27419;
wire  _GEN27424 = io_x[38] ? _GEN27423 : _GEN27416;
wire  _GEN27425 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27426 = io_x[27] ? _GEN21739 : _GEN27425;
wire  _GEN27427 = io_x[29] ? _GEN21743 : _GEN27426;
wire  _GEN27428 = io_x[75] ? _GEN27427 : _GEN21772;
wire  _GEN27429 = io_x[38] ? _GEN21833 : _GEN27428;
wire  _GEN27430 = io_x[34] ? _GEN27429 : _GEN27424;
wire  _GEN27431 = io_x[39] ? _GEN27430 : _GEN27409;
wire  _GEN27432 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN27433 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN27434 = io_x[75] ? _GEN21758 : _GEN27433;
wire  _GEN27435 = io_x[38] ? _GEN27434 : _GEN27432;
wire  _GEN27436 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27437 = io_x[27] ? _GEN21739 : _GEN27436;
wire  _GEN27438 = io_x[29] ? _GEN21743 : _GEN27437;
wire  _GEN27439 = io_x[75] ? _GEN27438 : _GEN21772;
wire  _GEN27440 = io_x[38] ? _GEN21871 : _GEN27439;
wire  _GEN27441 = io_x[34] ? _GEN27440 : _GEN27435;
wire  _GEN27442 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27443 = io_x[27] ? _GEN27442 : _GEN21739;
wire  _GEN27444 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27445 = io_x[29] ? _GEN27444 : _GEN27443;
wire  _GEN27446 = io_x[75] ? _GEN21758 : _GEN27445;
wire  _GEN27447 = io_x[38] ? _GEN27446 : _GEN21871;
wire  _GEN27448 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27449 = io_x[29] ? _GEN21744 : _GEN27448;
wire  _GEN27450 = io_x[75] ? _GEN21758 : _GEN27449;
wire  _GEN27451 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27452 = io_x[27] ? _GEN21750 : _GEN27451;
wire  _GEN27453 = io_x[29] ? _GEN21744 : _GEN27452;
wire  _GEN27454 = io_x[75] ? _GEN21772 : _GEN27453;
wire  _GEN27455 = io_x[38] ? _GEN27454 : _GEN27450;
wire  _GEN27456 = io_x[34] ? _GEN27455 : _GEN27447;
wire  _GEN27457 = io_x[39] ? _GEN27456 : _GEN27441;
wire  _GEN27458 = io_x[46] ? _GEN27457 : _GEN27431;
wire  _GEN27459 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27460 = io_x[27] ? _GEN21739 : _GEN27459;
wire  _GEN27461 = io_x[29] ? _GEN21743 : _GEN27460;
wire  _GEN27462 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27463 = io_x[27] ? _GEN27462 : _GEN21739;
wire  _GEN27464 = io_x[29] ? _GEN27463 : _GEN21744;
wire  _GEN27465 = io_x[75] ? _GEN27464 : _GEN27461;
wire  _GEN27466 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27467 = io_x[27] ? _GEN21739 : _GEN27466;
wire  _GEN27468 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27469 = io_x[27] ? _GEN27468 : _GEN21739;
wire  _GEN27470 = io_x[29] ? _GEN27469 : _GEN27467;
wire  _GEN27471 = io_x[75] ? _GEN21758 : _GEN27470;
wire  _GEN27472 = io_x[38] ? _GEN27471 : _GEN27465;
wire  _GEN27473 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN27474 = io_x[34] ? _GEN27473 : _GEN27472;
wire  _GEN27475 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN27476 = io_x[29] ? _GEN27475 : _GEN21743;
wire  _GEN27477 = io_x[75] ? _GEN21772 : _GEN27476;
wire  _GEN27478 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27479 = io_x[27] ? _GEN21750 : _GEN27478;
wire  _GEN27480 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27481 = io_x[29] ? _GEN27480 : _GEN27479;
wire  _GEN27482 = io_x[75] ? _GEN21758 : _GEN27481;
wire  _GEN27483 = io_x[38] ? _GEN27482 : _GEN27477;
wire  _GEN27484 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27485 = io_x[27] ? _GEN27484 : _GEN21739;
wire  _GEN27486 = io_x[29] ? _GEN27485 : _GEN21743;
wire  _GEN27487 = io_x[75] ? _GEN21758 : _GEN27486;
wire  _GEN27488 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27489 = io_x[27] ? _GEN27488 : _GEN21739;
wire  _GEN27490 = io_x[29] ? _GEN27489 : _GEN21743;
wire  _GEN27491 = io_x[75] ? _GEN21758 : _GEN27490;
wire  _GEN27492 = io_x[38] ? _GEN27491 : _GEN27487;
wire  _GEN27493 = io_x[34] ? _GEN27492 : _GEN27483;
wire  _GEN27494 = io_x[39] ? _GEN27493 : _GEN27474;
wire  _GEN27495 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN27496 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN27497 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27498 = io_x[27] ? _GEN27497 : _GEN21739;
wire  _GEN27499 = io_x[29] ? _GEN21743 : _GEN27498;
wire  _GEN27500 = io_x[75] ? _GEN27499 : _GEN27496;
wire  _GEN27501 = io_x[38] ? _GEN21871 : _GEN27500;
wire  _GEN27502 = io_x[34] ? _GEN27501 : _GEN27495;
wire  _GEN27503 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27504 = io_x[29] ? _GEN27503 : _GEN21744;
wire  _GEN27505 = io_x[75] ? _GEN21772 : _GEN27504;
wire  _GEN27506 = io_x[38] ? _GEN27505 : _GEN21871;
wire  _GEN27507 = io_x[34] ? _GEN21927 : _GEN27506;
wire  _GEN27508 = io_x[39] ? _GEN27507 : _GEN27502;
wire  _GEN27509 = io_x[46] ? _GEN27508 : _GEN27494;
wire  _GEN27510 = io_x[18] ? _GEN27509 : _GEN27458;
wire  _GEN27511 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN27512 = io_x[38] ? _GEN27511 : _GEN21871;
wire  _GEN27513 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN27514 = io_x[34] ? _GEN27513 : _GEN27512;
wire  _GEN27515 = io_x[39] ? _GEN27514 : _GEN21910;
wire  _GEN27516 = io_x[46] ? _GEN22145 : _GEN27515;
wire  _GEN27517 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN27518 = io_x[34] ? _GEN27517 : _GEN21927;
wire  _GEN27519 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27520 = io_x[27] ? _GEN21739 : _GEN27519;
wire  _GEN27521 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27522 = io_x[27] ? _GEN27521 : _GEN21739;
wire  _GEN27523 = io_x[29] ? _GEN27522 : _GEN27520;
wire  _GEN27524 = io_x[75] ? _GEN27523 : _GEN21758;
wire  _GEN27525 = io_x[38] ? _GEN21871 : _GEN27524;
wire  _GEN27526 = io_x[34] ? _GEN21927 : _GEN27525;
wire  _GEN27527 = io_x[39] ? _GEN27526 : _GEN27518;
wire  _GEN27528 = io_x[46] ? _GEN22145 : _GEN27527;
wire  _GEN27529 = io_x[18] ? _GEN27528 : _GEN27516;
wire  _GEN27530 = io_x[49] ? _GEN27529 : _GEN27510;
wire  _GEN27531 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27532 = io_x[27] ? _GEN21739 : _GEN27531;
wire  _GEN27533 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27534 = io_x[27] ? _GEN27533 : _GEN21739;
wire  _GEN27535 = io_x[29] ? _GEN27534 : _GEN27532;
wire  _GEN27536 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27537 = io_x[27] ? _GEN27536 : _GEN21739;
wire  _GEN27538 = io_x[29] ? _GEN27537 : _GEN21743;
wire  _GEN27539 = io_x[75] ? _GEN27538 : _GEN27535;
wire  _GEN27540 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27541 = io_x[29] ? _GEN27540 : _GEN21743;
wire  _GEN27542 = io_x[75] ? _GEN21758 : _GEN27541;
wire  _GEN27543 = io_x[38] ? _GEN27542 : _GEN27539;
wire  _GEN27544 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27545 = io_x[27] ? _GEN27544 : _GEN21750;
wire  _GEN27546 = io_x[29] ? _GEN27545 : _GEN21744;
wire  _GEN27547 = io_x[75] ? _GEN27546 : _GEN21772;
wire  _GEN27548 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27549 = io_x[27] ? _GEN27548 : _GEN21739;
wire  _GEN27550 = io_x[29] ? _GEN27549 : _GEN21743;
wire  _GEN27551 = io_x[75] ? _GEN21758 : _GEN27550;
wire  _GEN27552 = io_x[38] ? _GEN27551 : _GEN27547;
wire  _GEN27553 = io_x[34] ? _GEN27552 : _GEN27543;
wire  _GEN27554 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27555 = io_x[27] ? _GEN27554 : _GEN21750;
wire  _GEN27556 = io_x[29] ? _GEN27555 : _GEN21744;
wire  _GEN27557 = io_x[75] ? _GEN21772 : _GEN27556;
wire  _GEN27558 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27559 = io_x[27] ? _GEN27558 : _GEN21739;
wire  _GEN27560 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27561 = io_x[27] ? _GEN27560 : _GEN21750;
wire  _GEN27562 = io_x[29] ? _GEN27561 : _GEN27559;
wire  _GEN27563 = io_x[75] ? _GEN21758 : _GEN27562;
wire  _GEN27564 = io_x[38] ? _GEN27563 : _GEN27557;
wire  _GEN27565 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN27566 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27567 = io_x[29] ? _GEN27566 : _GEN21743;
wire  _GEN27568 = io_x[75] ? _GEN21758 : _GEN27567;
wire  _GEN27569 = io_x[38] ? _GEN27568 : _GEN27565;
wire  _GEN27570 = io_x[34] ? _GEN27569 : _GEN27564;
wire  _GEN27571 = io_x[39] ? _GEN27570 : _GEN27553;
wire  _GEN27572 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN27573 = io_x[75] ? _GEN27572 : _GEN21758;
wire  _GEN27574 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN27575 = io_x[38] ? _GEN27574 : _GEN27573;
wire  _GEN27576 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN27577 = io_x[75] ? _GEN21758 : _GEN27576;
wire  _GEN27578 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27579 = io_x[27] ? _GEN27578 : _GEN21739;
wire  _GEN27580 = io_x[29] ? _GEN27579 : _GEN21743;
wire  _GEN27581 = io_x[75] ? _GEN27580 : _GEN21758;
wire  _GEN27582 = io_x[38] ? _GEN27581 : _GEN27577;
wire  _GEN27583 = io_x[34] ? _GEN27582 : _GEN27575;
wire  _GEN27584 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN27585 = io_x[75] ? _GEN21758 : _GEN27584;
wire  _GEN27586 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27587 = io_x[27] ? _GEN21750 : _GEN27586;
wire  _GEN27588 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27589 = io_x[27] ? _GEN27588 : _GEN21739;
wire  _GEN27590 = io_x[29] ? _GEN27589 : _GEN27587;
wire  _GEN27591 = io_x[75] ? _GEN27590 : _GEN21772;
wire  _GEN27592 = io_x[38] ? _GEN27591 : _GEN27585;
wire  _GEN27593 = io_x[34] ? _GEN27592 : _GEN21766;
wire  _GEN27594 = io_x[39] ? _GEN27593 : _GEN27583;
wire  _GEN27595 = io_x[46] ? _GEN27594 : _GEN27571;
wire  _GEN27596 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27597 = io_x[27] ? _GEN21739 : _GEN27596;
wire  _GEN27598 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27599 = io_x[27] ? _GEN27598 : _GEN21739;
wire  _GEN27600 = io_x[29] ? _GEN27599 : _GEN27597;
wire  _GEN27601 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27602 = io_x[27] ? _GEN27601 : _GEN21739;
wire  _GEN27603 = io_x[29] ? _GEN27602 : _GEN21744;
wire  _GEN27604 = io_x[75] ? _GEN27603 : _GEN27600;
wire  _GEN27605 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27606 = io_x[27] ? _GEN27605 : _GEN21750;
wire  _GEN27607 = io_x[29] ? _GEN27606 : _GEN21744;
wire  _GEN27608 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27609 = io_x[29] ? _GEN21744 : _GEN27608;
wire  _GEN27610 = io_x[75] ? _GEN27609 : _GEN27607;
wire  _GEN27611 = io_x[38] ? _GEN27610 : _GEN27604;
wire  _GEN27612 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27613 = io_x[27] ? _GEN21750 : _GEN27612;
wire  _GEN27614 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27615 = io_x[27] ? _GEN27614 : _GEN21750;
wire  _GEN27616 = io_x[29] ? _GEN27615 : _GEN27613;
wire  _GEN27617 = io_x[75] ? _GEN27616 : _GEN21772;
wire  _GEN27618 = io_x[38] ? _GEN21833 : _GEN27617;
wire  _GEN27619 = io_x[34] ? _GEN27618 : _GEN27611;
wire  _GEN27620 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27621 = io_x[27] ? _GEN27620 : _GEN21739;
wire  _GEN27622 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27623 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27624 = io_x[27] ? _GEN27623 : _GEN27622;
wire  _GEN27625 = io_x[29] ? _GEN27624 : _GEN27621;
wire  _GEN27626 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27627 = io_x[27] ? _GEN27626 : _GEN21750;
wire  _GEN27628 = io_x[29] ? _GEN27627 : _GEN21743;
wire  _GEN27629 = io_x[75] ? _GEN27628 : _GEN27625;
wire  _GEN27630 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27631 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27632 = io_x[27] ? _GEN27631 : _GEN27630;
wire  _GEN27633 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27634 = io_x[27] ? _GEN27633 : _GEN21750;
wire  _GEN27635 = io_x[29] ? _GEN27634 : _GEN27632;
wire  _GEN27636 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27637 = io_x[27] ? _GEN27636 : _GEN21739;
wire  _GEN27638 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27639 = io_x[27] ? _GEN27638 : _GEN21739;
wire  _GEN27640 = io_x[29] ? _GEN27639 : _GEN27637;
wire  _GEN27641 = io_x[75] ? _GEN27640 : _GEN27635;
wire  _GEN27642 = io_x[38] ? _GEN27641 : _GEN27629;
wire  _GEN27643 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27644 = io_x[27] ? _GEN27643 : _GEN21739;
wire  _GEN27645 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27646 = io_x[27] ? _GEN27645 : _GEN21739;
wire  _GEN27647 = io_x[29] ? _GEN27646 : _GEN27644;
wire  _GEN27648 = io_x[75] ? _GEN27647 : _GEN21758;
wire  _GEN27649 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27650 = io_x[27] ? _GEN27649 : _GEN21739;
wire  _GEN27651 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27652 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27653 = io_x[27] ? _GEN27652 : _GEN27651;
wire  _GEN27654 = io_x[29] ? _GEN27653 : _GEN27650;
wire  _GEN27655 = io_x[75] ? _GEN21758 : _GEN27654;
wire  _GEN27656 = io_x[38] ? _GEN27655 : _GEN27648;
wire  _GEN27657 = io_x[34] ? _GEN27656 : _GEN27642;
wire  _GEN27658 = io_x[39] ? _GEN27657 : _GEN27619;
wire  _GEN27659 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27660 = io_x[27] ? _GEN27659 : _GEN21739;
wire  _GEN27661 = io_x[29] ? _GEN27660 : _GEN21743;
wire  _GEN27662 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27663 = io_x[27] ? _GEN21750 : _GEN27662;
wire  _GEN27664 = io_x[29] ? _GEN21744 : _GEN27663;
wire  _GEN27665 = io_x[75] ? _GEN27664 : _GEN27661;
wire  _GEN27666 = io_x[38] ? _GEN27665 : _GEN21871;
wire  _GEN27667 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27668 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27669 = io_x[27] ? _GEN27668 : _GEN27667;
wire  _GEN27670 = io_x[29] ? _GEN27669 : _GEN21743;
wire  _GEN27671 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27672 = io_x[27] ? _GEN27671 : _GEN21739;
wire  _GEN27673 = io_x[29] ? _GEN27672 : _GEN21743;
wire  _GEN27674 = io_x[75] ? _GEN27673 : _GEN27670;
wire  _GEN27675 = io_x[38] ? _GEN21871 : _GEN27674;
wire  _GEN27676 = io_x[34] ? _GEN27675 : _GEN27666;
wire  _GEN27677 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27678 = io_x[27] ? _GEN27677 : _GEN21750;
wire  _GEN27679 = io_x[29] ? _GEN27678 : _GEN21744;
wire  _GEN27680 = io_x[75] ? _GEN27679 : _GEN21758;
wire  _GEN27681 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27682 = io_x[27] ? _GEN21739 : _GEN27681;
wire  _GEN27683 = io_x[29] ? _GEN27682 : _GEN21743;
wire  _GEN27684 = io_x[75] ? _GEN21758 : _GEN27683;
wire  _GEN27685 = io_x[38] ? _GEN27684 : _GEN27680;
wire  _GEN27686 = io_x[34] ? _GEN21927 : _GEN27685;
wire  _GEN27687 = io_x[39] ? _GEN27686 : _GEN27676;
wire  _GEN27688 = io_x[46] ? _GEN27687 : _GEN27658;
wire  _GEN27689 = io_x[18] ? _GEN27688 : _GEN27595;
wire  _GEN27690 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN27691 = io_x[34] ? _GEN21927 : _GEN27690;
wire  _GEN27692 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27693 = io_x[27] ? _GEN27692 : _GEN21739;
wire  _GEN27694 = io_x[29] ? _GEN27693 : _GEN21744;
wire  _GEN27695 = io_x[75] ? _GEN27694 : _GEN21758;
wire  _GEN27696 = io_x[38] ? _GEN27695 : _GEN21833;
wire  _GEN27697 = io_x[34] ? _GEN21766 : _GEN27696;
wire  _GEN27698 = io_x[39] ? _GEN27697 : _GEN27691;
wire  _GEN27699 = io_x[46] ? _GEN22145 : _GEN27698;
wire  _GEN27700 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN27701 = io_x[34] ? _GEN27700 : _GEN21927;
wire  _GEN27702 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN27703 = io_x[38] ? _GEN21871 : _GEN27702;
wire  _GEN27704 = io_x[34] ? _GEN21927 : _GEN27703;
wire  _GEN27705 = io_x[39] ? _GEN27704 : _GEN27701;
wire  _GEN27706 = io_x[46] ? _GEN22145 : _GEN27705;
wire  _GEN27707 = io_x[18] ? _GEN27706 : _GEN27699;
wire  _GEN27708 = io_x[49] ? _GEN27707 : _GEN27689;
wire  _GEN27709 = io_x[24] ? _GEN27708 : _GEN27530;
wire  _GEN27710 = io_x[80] ? _GEN27709 : _GEN27389;
wire  _GEN27711 = io_x[16] ? _GEN27710 : _GEN26558;
wire  _GEN27712 = io_x[22] ? _GEN27711 : _GEN25679;
wire  _GEN27713 = io_x[20] ? _GEN27712 : _GEN24312;
wire  _GEN27714 = io_x[34] ? _GEN21766 : _GEN21927;
wire  _GEN27715 = io_x[39] ? _GEN21910 : _GEN27714;
wire  _GEN27716 = io_x[46] ? _GEN22145 : _GEN27715;
wire  _GEN27717 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN27718 = io_x[39] ? _GEN27717 : _GEN22327;
wire  _GEN27719 = io_x[46] ? _GEN22145 : _GEN27718;
wire  _GEN27720 = io_x[18] ? _GEN27719 : _GEN27716;
wire  _GEN27721 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN27722 = io_x[34] ? _GEN27721 : _GEN21766;
wire  _GEN27723 = io_x[39] ? _GEN21910 : _GEN27722;
wire  _GEN27724 = io_x[46] ? _GEN27723 : _GEN22145;
wire  _GEN27725 = io_x[39] ? _GEN22327 : _GEN21910;
wire  _GEN27726 = 1'b0;
wire  _GEN27727 = io_x[46] ? _GEN27726 : _GEN27725;
wire  _GEN27728 = io_x[18] ? _GEN27727 : _GEN27724;
wire  _GEN27729 = io_x[49] ? _GEN27728 : _GEN27720;
wire  _GEN27730 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN27731 = io_x[39] ? _GEN21910 : _GEN27730;
wire  _GEN27732 = io_x[46] ? _GEN27731 : _GEN22145;
wire  _GEN27733 = io_x[46] ? _GEN27726 : _GEN22145;
wire  _GEN27734 = io_x[18] ? _GEN27733 : _GEN27732;
wire  _GEN27735 = io_x[49] ? _GEN27734 : _GEN22268;
wire  _GEN27736 = io_x[24] ? _GEN27735 : _GEN27729;
wire  _GEN27737 = 1'b0;
wire  _GEN27738 = io_x[80] ? _GEN27737 : _GEN27736;
wire  _GEN27739 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN27740 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27741 = io_x[27] ? _GEN21739 : _GEN27740;
wire  _GEN27742 = io_x[29] ? _GEN21744 : _GEN27741;
wire  _GEN27743 = io_x[75] ? _GEN21758 : _GEN27742;
wire  _GEN27744 = io_x[38] ? _GEN27743 : _GEN21833;
wire  _GEN27745 = io_x[34] ? _GEN27744 : _GEN27739;
wire  _GEN27746 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN27747 = io_x[75] ? _GEN21758 : _GEN27746;
wire  _GEN27748 = io_x[38] ? _GEN27747 : _GEN21833;
wire  _GEN27749 = io_x[34] ? _GEN27748 : _GEN21766;
wire  _GEN27750 = io_x[39] ? _GEN27749 : _GEN27745;
wire  _GEN27751 = io_x[46] ? _GEN27726 : _GEN27750;
wire  _GEN27752 = io_x[18] ? _GEN27751 : _GEN23503;
wire  _GEN27753 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN27754 = io_x[34] ? _GEN21927 : _GEN27753;
wire  _GEN27755 = io_x[39] ? _GEN21910 : _GEN27754;
wire  _GEN27756 = io_x[46] ? _GEN27755 : _GEN22145;
wire  _GEN27757 = io_x[39] ? _GEN22327 : _GEN21910;
wire  _GEN27758 = io_x[46] ? _GEN27726 : _GEN27757;
wire  _GEN27759 = io_x[18] ? _GEN27758 : _GEN27756;
wire  _GEN27760 = io_x[49] ? _GEN27759 : _GEN27752;
wire  _GEN27761 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN27762 = io_x[75] ? _GEN21772 : _GEN27761;
wire  _GEN27763 = io_x[38] ? _GEN27762 : _GEN21833;
wire  _GEN27764 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27765 = io_x[27] ? _GEN27764 : _GEN21739;
wire  _GEN27766 = io_x[29] ? _GEN21744 : _GEN27765;
wire  _GEN27767 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN27768 = io_x[75] ? _GEN27767 : _GEN27766;
wire  _GEN27769 = io_x[38] ? _GEN27768 : _GEN21833;
wire  _GEN27770 = io_x[34] ? _GEN27769 : _GEN27763;
wire  _GEN27771 = io_x[39] ? _GEN22327 : _GEN27770;
wire  _GEN27772 = io_x[46] ? _GEN22145 : _GEN27771;
wire  _GEN27773 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27774 = io_x[27] ? _GEN21739 : _GEN27773;
wire  _GEN27775 = io_x[29] ? _GEN21743 : _GEN27774;
wire  _GEN27776 = io_x[75] ? _GEN21758 : _GEN27775;
wire  _GEN27777 = io_x[38] ? _GEN27776 : _GEN21833;
wire  _GEN27778 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27779 = io_x[27] ? _GEN21750 : _GEN27778;
wire  _GEN27780 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27781 = io_x[27] ? _GEN27780 : _GEN21739;
wire  _GEN27782 = io_x[29] ? _GEN27781 : _GEN27779;
wire  _GEN27783 = io_x[75] ? _GEN21758 : _GEN27782;
wire  _GEN27784 = io_x[38] ? _GEN27783 : _GEN21871;
wire  _GEN27785 = io_x[34] ? _GEN27784 : _GEN27777;
wire  _GEN27786 = io_x[39] ? _GEN22327 : _GEN27785;
wire  _GEN27787 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN27788 = io_x[39] ? _GEN27787 : _GEN22327;
wire  _GEN27789 = io_x[46] ? _GEN27788 : _GEN27786;
wire  _GEN27790 = io_x[18] ? _GEN27789 : _GEN27772;
wire  _GEN27791 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN27792 = io_x[46] ? _GEN27791 : _GEN22145;
wire  _GEN27793 = io_x[18] ? _GEN27792 : _GEN23503;
wire  _GEN27794 = io_x[49] ? _GEN27793 : _GEN27790;
wire  _GEN27795 = io_x[24] ? _GEN27794 : _GEN27760;
wire  _GEN27796 = io_x[34] ? _GEN21766 : _GEN21927;
wire  _GEN27797 = io_x[39] ? _GEN21910 : _GEN27796;
wire  _GEN27798 = io_x[46] ? _GEN22145 : _GEN27797;
wire  _GEN27799 = io_x[18] ? _GEN27798 : _GEN23503;
wire  _GEN27800 = io_x[49] ? _GEN22268 : _GEN27799;
wire  _GEN27801 = 1'b1;
wire  _GEN27802 = io_x[24] ? _GEN27801 : _GEN27800;
wire  _GEN27803 = io_x[80] ? _GEN27802 : _GEN27795;
wire  _GEN27804 = io_x[16] ? _GEN27803 : _GEN27738;
wire  _GEN27805 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN27806 = io_x[39] ? _GEN21910 : _GEN27805;
wire  _GEN27807 = io_x[46] ? _GEN27806 : _GEN22145;
wire  _GEN27808 = io_x[46] ? _GEN27726 : _GEN22145;
wire  _GEN27809 = io_x[18] ? _GEN27808 : _GEN27807;
wire  _GEN27810 = io_x[49] ? _GEN27809 : _GEN22268;
wire  _GEN27811 = io_x[39] ? _GEN22327 : _GEN21910;
wire  _GEN27812 = io_x[46] ? _GEN22145 : _GEN27811;
wire  _GEN27813 = io_x[39] ? _GEN22327 : _GEN21910;
wire  _GEN27814 = io_x[46] ? _GEN22145 : _GEN27813;
wire  _GEN27815 = io_x[18] ? _GEN27814 : _GEN27812;
wire  _GEN27816 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN27817 = io_x[46] ? _GEN27816 : _GEN22145;
wire  _GEN27818 = io_x[46] ? _GEN27726 : _GEN22145;
wire  _GEN27819 = io_x[18] ? _GEN27818 : _GEN27817;
wire  _GEN27820 = io_x[49] ? _GEN27819 : _GEN27815;
wire  _GEN27821 = io_x[24] ? _GEN27820 : _GEN27810;
wire  _GEN27822 = 1'b0;
wire  _GEN27823 = 1'b1;
wire  _GEN27824 = io_x[49] ? _GEN27823 : _GEN22268;
wire  _GEN27825 = io_x[24] ? _GEN27824 : _GEN27822;
wire  _GEN27826 = io_x[80] ? _GEN27825 : _GEN27821;
wire  _GEN27827 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27828 = io_x[27] ? _GEN27827 : _GEN21739;
wire  _GEN27829 = io_x[29] ? _GEN27828 : _GEN21744;
wire  _GEN27830 = io_x[75] ? _GEN21758 : _GEN27829;
wire  _GEN27831 = io_x[38] ? _GEN27830 : _GEN21833;
wire  _GEN27832 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27833 = io_x[27] ? _GEN27832 : _GEN21739;
wire  _GEN27834 = io_x[29] ? _GEN27833 : _GEN21743;
wire  _GEN27835 = io_x[75] ? _GEN21758 : _GEN27834;
wire  _GEN27836 = io_x[38] ? _GEN27835 : _GEN21833;
wire  _GEN27837 = io_x[34] ? _GEN27836 : _GEN27831;
wire  _GEN27838 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27839 = io_x[29] ? _GEN27838 : _GEN21743;
wire  _GEN27840 = io_x[75] ? _GEN21758 : _GEN27839;
wire  _GEN27841 = io_x[38] ? _GEN27840 : _GEN21833;
wire  _GEN27842 = io_x[34] ? _GEN27841 : _GEN21927;
wire  _GEN27843 = io_x[39] ? _GEN27842 : _GEN27837;
wire  _GEN27844 = io_x[46] ? _GEN22145 : _GEN27843;
wire  _GEN27845 = io_x[34] ? _GEN21766 : _GEN21927;
wire  _GEN27846 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27847 = io_x[27] ? _GEN27846 : _GEN21739;
wire  _GEN27848 = io_x[29] ? _GEN27847 : _GEN21744;
wire  _GEN27849 = io_x[75] ? _GEN21758 : _GEN27848;
wire  _GEN27850 = io_x[38] ? _GEN27849 : _GEN21871;
wire  _GEN27851 = io_x[34] ? _GEN21766 : _GEN27850;
wire  _GEN27852 = io_x[39] ? _GEN27851 : _GEN27845;
wire  _GEN27853 = io_x[46] ? _GEN22145 : _GEN27852;
wire  _GEN27854 = io_x[18] ? _GEN27853 : _GEN27844;
wire  _GEN27855 = io_x[39] ? _GEN22327 : _GEN21910;
wire  _GEN27856 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN27857 = io_x[46] ? _GEN27856 : _GEN27855;
wire  _GEN27858 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN27859 = io_x[46] ? _GEN27858 : _GEN27726;
wire  _GEN27860 = io_x[18] ? _GEN27859 : _GEN27857;
wire  _GEN27861 = io_x[49] ? _GEN27860 : _GEN27854;
wire  _GEN27862 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27863 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27864 = io_x[27] ? _GEN27863 : _GEN21739;
wire  _GEN27865 = io_x[29] ? _GEN27864 : _GEN27862;
wire  _GEN27866 = io_x[75] ? _GEN21758 : _GEN27865;
wire  _GEN27867 = io_x[38] ? _GEN27866 : _GEN21833;
wire  _GEN27868 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27869 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27870 = io_x[27] ? _GEN27869 : _GEN27868;
wire  _GEN27871 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27872 = io_x[27] ? _GEN27871 : _GEN21739;
wire  _GEN27873 = io_x[29] ? _GEN27872 : _GEN27870;
wire  _GEN27874 = io_x[75] ? _GEN21772 : _GEN27873;
wire  _GEN27875 = io_x[38] ? _GEN27874 : _GEN21833;
wire  _GEN27876 = io_x[34] ? _GEN27875 : _GEN27867;
wire  _GEN27877 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN27878 = io_x[29] ? _GEN21743 : _GEN27877;
wire  _GEN27879 = io_x[75] ? _GEN21758 : _GEN27878;
wire  _GEN27880 = io_x[38] ? _GEN27879 : _GEN21833;
wire  _GEN27881 = io_x[34] ? _GEN27880 : _GEN21927;
wire  _GEN27882 = io_x[39] ? _GEN27881 : _GEN27876;
wire  _GEN27883 = io_x[46] ? _GEN22145 : _GEN27882;
wire  _GEN27884 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27885 = io_x[27] ? _GEN21739 : _GEN27884;
wire  _GEN27886 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27887 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27888 = io_x[27] ? _GEN27887 : _GEN27886;
wire  _GEN27889 = io_x[29] ? _GEN27888 : _GEN27885;
wire  _GEN27890 = io_x[75] ? _GEN21758 : _GEN27889;
wire  _GEN27891 = io_x[38] ? _GEN27890 : _GEN21833;
wire  _GEN27892 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27893 = io_x[27] ? _GEN27892 : _GEN21739;
wire  _GEN27894 = io_x[29] ? _GEN27893 : _GEN21743;
wire  _GEN27895 = io_x[75] ? _GEN27894 : _GEN21772;
wire  _GEN27896 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27897 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27898 = io_x[27] ? _GEN27897 : _GEN27896;
wire  _GEN27899 = io_x[29] ? _GEN27898 : _GEN21744;
wire  _GEN27900 = io_x[75] ? _GEN21758 : _GEN27899;
wire  _GEN27901 = io_x[38] ? _GEN27900 : _GEN27895;
wire  _GEN27902 = io_x[34] ? _GEN27901 : _GEN27891;
wire  _GEN27903 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27904 = io_x[27] ? _GEN27903 : _GEN21750;
wire  _GEN27905 = io_x[29] ? _GEN27904 : _GEN21744;
wire  _GEN27906 = io_x[75] ? _GEN21758 : _GEN27905;
wire  _GEN27907 = io_x[38] ? _GEN27906 : _GEN21833;
wire  _GEN27908 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN27909 = io_x[29] ? _GEN27908 : _GEN21743;
wire  _GEN27910 = io_x[75] ? _GEN21758 : _GEN27909;
wire  _GEN27911 = io_x[38] ? _GEN27910 : _GEN21871;
wire  _GEN27912 = io_x[34] ? _GEN27911 : _GEN27907;
wire  _GEN27913 = io_x[39] ? _GEN27912 : _GEN27902;
wire  _GEN27914 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN27915 = io_x[38] ? _GEN21833 : _GEN27914;
wire  _GEN27916 = io_x[34] ? _GEN21927 : _GEN27915;
wire  _GEN27917 = io_x[39] ? _GEN27916 : _GEN22327;
wire  _GEN27918 = io_x[46] ? _GEN27917 : _GEN27913;
wire  _GEN27919 = io_x[18] ? _GEN27918 : _GEN27883;
wire  _GEN27920 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27921 = io_x[27] ? _GEN27920 : _GEN21739;
wire  _GEN27922 = io_x[29] ? _GEN27921 : _GEN21743;
wire  _GEN27923 = io_x[75] ? _GEN21758 : _GEN27922;
wire  _GEN27924 = io_x[38] ? _GEN21833 : _GEN27923;
wire  _GEN27925 = io_x[34] ? _GEN21927 : _GEN27924;
wire  _GEN27926 = io_x[39] ? _GEN27925 : _GEN21910;
wire  _GEN27927 = io_x[46] ? _GEN22145 : _GEN27926;
wire  _GEN27928 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN27929 = io_x[38] ? _GEN21833 : _GEN27928;
wire  _GEN27930 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27931 = io_x[27] ? _GEN27930 : _GEN21739;
wire  _GEN27932 = io_x[29] ? _GEN27931 : _GEN21743;
wire  _GEN27933 = io_x[75] ? _GEN21758 : _GEN27932;
wire  _GEN27934 = io_x[38] ? _GEN27933 : _GEN21833;
wire  _GEN27935 = io_x[34] ? _GEN27934 : _GEN27929;
wire  _GEN27936 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN27937 = io_x[39] ? _GEN27936 : _GEN27935;
wire  _GEN27938 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN27939 = io_x[46] ? _GEN27938 : _GEN27937;
wire  _GEN27940 = io_x[18] ? _GEN27939 : _GEN27927;
wire  _GEN27941 = io_x[49] ? _GEN27940 : _GEN27919;
wire  _GEN27942 = io_x[24] ? _GEN27941 : _GEN27861;
wire  _GEN27943 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN27944 = io_x[38] ? _GEN27943 : _GEN21833;
wire  _GEN27945 = io_x[34] ? _GEN21927 : _GEN27944;
wire  _GEN27946 = io_x[39] ? _GEN27945 : _GEN21910;
wire  _GEN27947 = io_x[46] ? _GEN22145 : _GEN27946;
wire  _GEN27948 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN27949 = io_x[34] ? _GEN21927 : _GEN27948;
wire  _GEN27950 = io_x[39] ? _GEN27949 : _GEN21910;
wire  _GEN27951 = io_x[46] ? _GEN22145 : _GEN27950;
wire  _GEN27952 = io_x[18] ? _GEN27951 : _GEN27947;
wire  _GEN27953 = io_x[49] ? _GEN22268 : _GEN27952;
wire  _GEN27954 = io_x[24] ? _GEN27953 : _GEN27801;
wire  _GEN27955 = io_x[80] ? _GEN27954 : _GEN27942;
wire  _GEN27956 = io_x[16] ? _GEN27955 : _GEN27826;
wire  _GEN27957 = io_x[22] ? _GEN27956 : _GEN27804;
wire  _GEN27958 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN27959 = io_x[34] ? _GEN21927 : _GEN27958;
wire  _GEN27960 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN27961 = io_x[34] ? _GEN27960 : _GEN21927;
wire  _GEN27962 = io_x[39] ? _GEN27961 : _GEN27959;
wire  _GEN27963 = io_x[46] ? _GEN22145 : _GEN27962;
wire  _GEN27964 = io_x[18] ? _GEN27963 : _GEN23503;
wire  _GEN27965 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN27966 = io_x[46] ? _GEN27965 : _GEN22145;
wire  _GEN27967 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN27968 = io_x[46] ? _GEN27967 : _GEN22145;
wire  _GEN27969 = io_x[18] ? _GEN27968 : _GEN27966;
wire  _GEN27970 = io_x[49] ? _GEN27969 : _GEN27964;
wire  _GEN27971 = io_x[46] ? _GEN27726 : _GEN22145;
wire  _GEN27972 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN27973 = io_x[38] ? _GEN27972 : _GEN21833;
wire  _GEN27974 = io_x[34] ? _GEN21927 : _GEN27973;
wire  _GEN27975 = io_x[39] ? _GEN21910 : _GEN27974;
wire  _GEN27976 = io_x[46] ? _GEN27975 : _GEN22145;
wire  _GEN27977 = io_x[18] ? _GEN27976 : _GEN27971;
wire  _GEN27978 = io_x[49] ? _GEN27977 : _GEN22268;
wire  _GEN27979 = io_x[24] ? _GEN27978 : _GEN27970;
wire  _GEN27980 = io_x[18] ? _GEN23503 : _GEN24190;
wire  _GEN27981 = io_x[49] ? _GEN27823 : _GEN27980;
wire  _GEN27982 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN27983 = io_x[39] ? _GEN27982 : _GEN21910;
wire  _GEN27984 = io_x[46] ? _GEN22145 : _GEN27983;
wire  _GEN27985 = io_x[18] ? _GEN27984 : _GEN24190;
wire  _GEN27986 = io_x[49] ? _GEN27823 : _GEN27985;
wire  _GEN27987 = io_x[24] ? _GEN27986 : _GEN27981;
wire  _GEN27988 = io_x[80] ? _GEN27987 : _GEN27979;
wire  _GEN27989 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27990 = io_x[27] ? _GEN27989 : _GEN21739;
wire  _GEN27991 = io_x[29] ? _GEN21743 : _GEN27990;
wire  _GEN27992 = io_x[75] ? _GEN21758 : _GEN27991;
wire  _GEN27993 = io_x[38] ? _GEN27992 : _GEN21833;
wire  _GEN27994 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN27995 = io_x[27] ? _GEN27994 : _GEN21739;
wire  _GEN27996 = io_x[29] ? _GEN27995 : _GEN21744;
wire  _GEN27997 = io_x[75] ? _GEN21758 : _GEN27996;
wire  _GEN27998 = io_x[38] ? _GEN27997 : _GEN21871;
wire  _GEN27999 = io_x[34] ? _GEN27998 : _GEN27993;
wire  _GEN28000 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28001 = io_x[27] ? _GEN21739 : _GEN28000;
wire  _GEN28002 = io_x[29] ? _GEN21744 : _GEN28001;
wire  _GEN28003 = io_x[75] ? _GEN21758 : _GEN28002;
wire  _GEN28004 = io_x[38] ? _GEN28003 : _GEN21871;
wire  _GEN28005 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN28006 = io_x[75] ? _GEN21772 : _GEN28005;
wire  _GEN28007 = io_x[38] ? _GEN21833 : _GEN28006;
wire  _GEN28008 = io_x[34] ? _GEN28007 : _GEN28004;
wire  _GEN28009 = io_x[39] ? _GEN28008 : _GEN27999;
wire  _GEN28010 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN28011 = io_x[38] ? _GEN21833 : _GEN28010;
wire  _GEN28012 = io_x[34] ? _GEN21927 : _GEN28011;
wire  _GEN28013 = io_x[39] ? _GEN28012 : _GEN22327;
wire  _GEN28014 = io_x[46] ? _GEN28013 : _GEN28009;
wire  _GEN28015 = io_x[18] ? _GEN28014 : _GEN23503;
wire  _GEN28016 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN28017 = io_x[46] ? _GEN28016 : _GEN22145;
wire  _GEN28018 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN28019 = io_x[34] ? _GEN28018 : _GEN21766;
wire  _GEN28020 = io_x[39] ? _GEN28019 : _GEN21910;
wire  _GEN28021 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN28022 = io_x[46] ? _GEN28021 : _GEN28020;
wire  _GEN28023 = io_x[18] ? _GEN28022 : _GEN28017;
wire  _GEN28024 = io_x[49] ? _GEN28023 : _GEN28015;
wire  _GEN28025 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN28026 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28027 = io_x[27] ? _GEN28026 : _GEN21739;
wire  _GEN28028 = io_x[29] ? _GEN28027 : _GEN21743;
wire  _GEN28029 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28030 = io_x[27] ? _GEN28029 : _GEN21750;
wire  _GEN28031 = io_x[29] ? _GEN28030 : _GEN21743;
wire  _GEN28032 = io_x[75] ? _GEN28031 : _GEN28028;
wire  _GEN28033 = io_x[38] ? _GEN28032 : _GEN21833;
wire  _GEN28034 = io_x[34] ? _GEN28033 : _GEN28025;
wire  _GEN28035 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28036 = io_x[27] ? _GEN28035 : _GEN21739;
wire  _GEN28037 = io_x[29] ? _GEN28036 : _GEN21743;
wire  _GEN28038 = io_x[75] ? _GEN21758 : _GEN28037;
wire  _GEN28039 = io_x[38] ? _GEN28038 : _GEN21871;
wire  _GEN28040 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28041 = io_x[27] ? _GEN28040 : _GEN21739;
wire  _GEN28042 = io_x[29] ? _GEN28041 : _GEN21743;
wire  _GEN28043 = io_x[75] ? _GEN21758 : _GEN28042;
wire  _GEN28044 = io_x[38] ? _GEN28043 : _GEN21833;
wire  _GEN28045 = io_x[34] ? _GEN28044 : _GEN28039;
wire  _GEN28046 = io_x[39] ? _GEN28045 : _GEN28034;
wire  _GEN28047 = io_x[46] ? _GEN22145 : _GEN28046;
wire  _GEN28048 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28049 = io_x[27] ? _GEN28048 : _GEN21739;
wire  _GEN28050 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28051 = io_x[27] ? _GEN28050 : _GEN21739;
wire  _GEN28052 = io_x[29] ? _GEN28051 : _GEN28049;
wire  _GEN28053 = io_x[75] ? _GEN21758 : _GEN28052;
wire  _GEN28054 = io_x[38] ? _GEN28053 : _GEN21833;
wire  _GEN28055 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28056 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28057 = io_x[27] ? _GEN28056 : _GEN28055;
wire  _GEN28058 = io_x[29] ? _GEN28057 : _GEN21744;
wire  _GEN28059 = io_x[75] ? _GEN21758 : _GEN28058;
wire  _GEN28060 = io_x[38] ? _GEN28059 : _GEN21871;
wire  _GEN28061 = io_x[34] ? _GEN28060 : _GEN28054;
wire  _GEN28062 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28063 = io_x[27] ? _GEN28062 : _GEN21739;
wire  _GEN28064 = io_x[29] ? _GEN28063 : _GEN21743;
wire  _GEN28065 = io_x[75] ? _GEN21758 : _GEN28064;
wire  _GEN28066 = io_x[38] ? _GEN28065 : _GEN21833;
wire  _GEN28067 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28068 = io_x[27] ? _GEN28067 : _GEN21739;
wire  _GEN28069 = io_x[29] ? _GEN28068 : _GEN21743;
wire  _GEN28070 = io_x[75] ? _GEN21758 : _GEN28069;
wire  _GEN28071 = io_x[38] ? _GEN21871 : _GEN28070;
wire  _GEN28072 = io_x[34] ? _GEN28071 : _GEN28066;
wire  _GEN28073 = io_x[39] ? _GEN28072 : _GEN28061;
wire  _GEN28074 = io_x[27] ? _GEN21750 : _GEN21739;
wire  _GEN28075 = io_x[29] ? _GEN28074 : _GEN21743;
wire  _GEN28076 = io_x[75] ? _GEN28075 : _GEN21758;
wire  _GEN28077 = io_x[38] ? _GEN28076 : _GEN21833;
wire  _GEN28078 = io_x[34] ? _GEN28077 : _GEN21927;
wire  _GEN28079 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN28080 = io_x[38] ? _GEN21833 : _GEN28079;
wire  _GEN28081 = io_x[34] ? _GEN21927 : _GEN28080;
wire  _GEN28082 = io_x[39] ? _GEN28081 : _GEN28078;
wire  _GEN28083 = io_x[46] ? _GEN28082 : _GEN28073;
wire  _GEN28084 = io_x[18] ? _GEN28083 : _GEN28047;
wire  _GEN28085 = io_x[46] ? _GEN27726 : _GEN22145;
wire  _GEN28086 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28087 = io_x[27] ? _GEN21739 : _GEN28086;
wire  _GEN28088 = io_x[29] ? _GEN28087 : _GEN21743;
wire  _GEN28089 = io_x[75] ? _GEN28088 : _GEN21758;
wire  _GEN28090 = io_x[38] ? _GEN28089 : _GEN21833;
wire  _GEN28091 = io_x[34] ? _GEN28090 : _GEN21927;
wire  _GEN28092 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN28093 = io_x[39] ? _GEN28092 : _GEN28091;
wire  _GEN28094 = io_x[46] ? _GEN27726 : _GEN28093;
wire  _GEN28095 = io_x[18] ? _GEN28094 : _GEN28085;
wire  _GEN28096 = io_x[49] ? _GEN28095 : _GEN28084;
wire  _GEN28097 = io_x[24] ? _GEN28096 : _GEN28024;
wire  _GEN28098 = io_x[39] ? _GEN22327 : _GEN21910;
wire  _GEN28099 = io_x[46] ? _GEN22145 : _GEN28098;
wire  _GEN28100 = io_x[18] ? _GEN28099 : _GEN24190;
wire  _GEN28101 = io_x[49] ? _GEN28100 : _GEN27823;
wire  _GEN28102 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN28103 = io_x[38] ? _GEN21833 : _GEN28102;
wire  _GEN28104 = io_x[34] ? _GEN21927 : _GEN28103;
wire  _GEN28105 = io_x[39] ? _GEN28104 : _GEN21910;
wire  _GEN28106 = io_x[46] ? _GEN22145 : _GEN28105;
wire  _GEN28107 = io_x[18] ? _GEN28106 : _GEN24190;
wire  _GEN28108 = io_x[49] ? _GEN22268 : _GEN28107;
wire  _GEN28109 = io_x[24] ? _GEN28108 : _GEN28101;
wire  _GEN28110 = io_x[80] ? _GEN28109 : _GEN28097;
wire  _GEN28111 = io_x[16] ? _GEN28110 : _GEN27988;
wire  _GEN28112 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN28113 = io_x[38] ? _GEN28112 : _GEN21833;
wire  _GEN28114 = io_x[34] ? _GEN21927 : _GEN28113;
wire  _GEN28115 = io_x[38] ? _GEN21871 : _GEN21833;
wire  _GEN28116 = io_x[34] ? _GEN21927 : _GEN28115;
wire  _GEN28117 = io_x[39] ? _GEN28116 : _GEN28114;
wire  _GEN28118 = io_x[46] ? _GEN27726 : _GEN28117;
wire  _GEN28119 = io_x[18] ? _GEN28118 : _GEN23503;
wire  _GEN28120 = io_x[46] ? _GEN27726 : _GEN22145;
wire  _GEN28121 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN28122 = io_x[46] ? _GEN28121 : _GEN22145;
wire  _GEN28123 = io_x[18] ? _GEN28122 : _GEN28120;
wire  _GEN28124 = io_x[49] ? _GEN28123 : _GEN28119;
wire  _GEN28125 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN28126 = io_x[38] ? _GEN28125 : _GEN21833;
wire  _GEN28127 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN28128 = io_x[38] ? _GEN28127 : _GEN21833;
wire  _GEN28129 = io_x[34] ? _GEN28128 : _GEN28126;
wire  _GEN28130 = io_x[39] ? _GEN22327 : _GEN28129;
wire  _GEN28131 = io_x[46] ? _GEN27726 : _GEN28130;
wire  _GEN28132 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28133 = io_x[27] ? _GEN28132 : _GEN21739;
wire  _GEN28134 = io_x[29] ? _GEN28133 : _GEN21743;
wire  _GEN28135 = io_x[75] ? _GEN28134 : _GEN21772;
wire  _GEN28136 = io_x[38] ? _GEN28135 : _GEN21871;
wire  _GEN28137 = io_x[34] ? _GEN21927 : _GEN28136;
wire  _GEN28138 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN28139 = io_x[39] ? _GEN28138 : _GEN28137;
wire  _GEN28140 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN28141 = io_x[39] ? _GEN28140 : _GEN21910;
wire  _GEN28142 = io_x[46] ? _GEN28141 : _GEN28139;
wire  _GEN28143 = io_x[18] ? _GEN28142 : _GEN28131;
wire  _GEN28144 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN28145 = io_x[34] ? _GEN21927 : _GEN28144;
wire  _GEN28146 = io_x[39] ? _GEN28145 : _GEN21910;
wire  _GEN28147 = io_x[46] ? _GEN27726 : _GEN28146;
wire  _GEN28148 = io_x[34] ? _GEN21766 : _GEN21927;
wire  _GEN28149 = io_x[39] ? _GEN28148 : _GEN21910;
wire  _GEN28150 = io_x[46] ? _GEN27726 : _GEN28149;
wire  _GEN28151 = io_x[18] ? _GEN28150 : _GEN28147;
wire  _GEN28152 = io_x[49] ? _GEN28151 : _GEN28143;
wire  _GEN28153 = io_x[24] ? _GEN28152 : _GEN28124;
wire  _GEN28154 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN28155 = io_x[46] ? _GEN28154 : _GEN27726;
wire  _GEN28156 = io_x[18] ? _GEN24190 : _GEN28155;
wire  _GEN28157 = io_x[49] ? _GEN22268 : _GEN28156;
wire  _GEN28158 = io_x[24] ? _GEN28157 : _GEN27801;
wire  _GEN28159 = io_x[80] ? _GEN28158 : _GEN28153;
wire  _GEN28160 = io_x[34] ? _GEN21766 : _GEN21927;
wire  _GEN28161 = io_x[29] ? _GEN21744 : _GEN21743;
wire  _GEN28162 = io_x[75] ? _GEN21758 : _GEN28161;
wire  _GEN28163 = io_x[38] ? _GEN28162 : _GEN21833;
wire  _GEN28164 = io_x[34] ? _GEN28163 : _GEN21927;
wire  _GEN28165 = io_x[39] ? _GEN28164 : _GEN28160;
wire  _GEN28166 = io_x[46] ? _GEN22145 : _GEN28165;
wire  _GEN28167 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28168 = io_x[27] ? _GEN28167 : _GEN21739;
wire  _GEN28169 = io_x[29] ? _GEN28168 : _GEN21744;
wire  _GEN28170 = io_x[75] ? _GEN21758 : _GEN28169;
wire  _GEN28171 = io_x[38] ? _GEN28170 : _GEN21833;
wire  _GEN28172 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28173 = io_x[27] ? _GEN28172 : _GEN21750;
wire  _GEN28174 = io_x[29] ? _GEN28173 : _GEN21744;
wire  _GEN28175 = io_x[75] ? _GEN21758 : _GEN28174;
wire  _GEN28176 = io_x[38] ? _GEN28175 : _GEN21871;
wire  _GEN28177 = io_x[34] ? _GEN28176 : _GEN28171;
wire  _GEN28178 = io_x[39] ? _GEN22327 : _GEN28177;
wire  _GEN28179 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN28180 = io_x[38] ? _GEN28179 : _GEN21871;
wire  _GEN28181 = io_x[34] ? _GEN28180 : _GEN21927;
wire  _GEN28182 = io_x[39] ? _GEN21910 : _GEN28181;
wire  _GEN28183 = io_x[46] ? _GEN28182 : _GEN28178;
wire  _GEN28184 = io_x[18] ? _GEN28183 : _GEN28166;
wire  _GEN28185 = io_x[39] ? _GEN22327 : _GEN21910;
wire  _GEN28186 = io_x[46] ? _GEN22145 : _GEN28185;
wire  _GEN28187 = io_x[38] ? _GEN21833 : _GEN21871;
wire  _GEN28188 = io_x[34] ? _GEN28187 : _GEN21927;
wire  _GEN28189 = io_x[34] ? _GEN21927 : _GEN21766;
wire  _GEN28190 = io_x[39] ? _GEN28189 : _GEN28188;
wire  _GEN28191 = io_x[46] ? _GEN27726 : _GEN28190;
wire  _GEN28192 = io_x[18] ? _GEN28191 : _GEN28186;
wire  _GEN28193 = io_x[49] ? _GEN28192 : _GEN28184;
wire  _GEN28194 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28195 = io_x[27] ? _GEN28194 : _GEN21739;
wire  _GEN28196 = io_x[29] ? _GEN28195 : _GEN21744;
wire  _GEN28197 = io_x[75] ? _GEN28196 : _GEN21758;
wire  _GEN28198 = io_x[38] ? _GEN28197 : _GEN21833;
wire  _GEN28199 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28200 = io_x[27] ? _GEN28199 : _GEN21750;
wire  _GEN28201 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28202 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28203 = io_x[27] ? _GEN28202 : _GEN28201;
wire  _GEN28204 = io_x[29] ? _GEN28203 : _GEN28200;
wire  _GEN28205 = io_x[75] ? _GEN21758 : _GEN28204;
wire  _GEN28206 = io_x[38] ? _GEN28205 : _GEN21833;
wire  _GEN28207 = io_x[34] ? _GEN28206 : _GEN28198;
wire  _GEN28208 = io_x[39] ? _GEN21910 : _GEN28207;
wire  _GEN28209 = io_x[39] ? _GEN21910 : _GEN22327;
wire  _GEN28210 = io_x[46] ? _GEN28209 : _GEN28208;
wire  _GEN28211 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28212 = io_x[27] ? _GEN28211 : _GEN21739;
wire  _GEN28213 = io_x[29] ? _GEN28212 : _GEN21743;
wire  _GEN28214 = io_x[75] ? _GEN21758 : _GEN28213;
wire  _GEN28215 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28216 = io_x[27] ? _GEN28215 : _GEN21739;
wire  _GEN28217 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28218 = io_x[27] ? _GEN28217 : _GEN21739;
wire  _GEN28219 = io_x[29] ? _GEN28218 : _GEN28216;
wire  _GEN28220 = io_x[75] ? _GEN21758 : _GEN28219;
wire  _GEN28221 = io_x[38] ? _GEN28220 : _GEN28214;
wire  _GEN28222 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28223 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28224 = io_x[27] ? _GEN28223 : _GEN28222;
wire  _GEN28225 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28226 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28227 = io_x[27] ? _GEN28226 : _GEN28225;
wire  _GEN28228 = io_x[29] ? _GEN28227 : _GEN28224;
wire  _GEN28229 = io_x[75] ? _GEN21758 : _GEN28228;
wire  _GEN28230 = io_x[38] ? _GEN28229 : _GEN21871;
wire  _GEN28231 = io_x[34] ? _GEN28230 : _GEN28221;
wire  _GEN28232 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28233 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28234 = io_x[27] ? _GEN28233 : _GEN28232;
wire  _GEN28235 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28236 = io_x[27] ? _GEN28235 : _GEN21750;
wire  _GEN28237 = io_x[29] ? _GEN28236 : _GEN28234;
wire  _GEN28238 = io_x[75] ? _GEN21758 : _GEN28237;
wire  _GEN28239 = io_x[38] ? _GEN28238 : _GEN21871;
wire  _GEN28240 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28241 = io_x[27] ? _GEN28240 : _GEN21750;
wire  _GEN28242 = io_x[29] ? _GEN28241 : _GEN21744;
wire  _GEN28243 = io_x[75] ? _GEN21772 : _GEN28242;
wire  _GEN28244 = io_x[27] ? _GEN21739 : _GEN21750;
wire  _GEN28245 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28246 = io_x[27] ? _GEN28245 : _GEN21739;
wire  _GEN28247 = io_x[29] ? _GEN28246 : _GEN28244;
wire  _GEN28248 = io_x[75] ? _GEN21758 : _GEN28247;
wire  _GEN28249 = io_x[38] ? _GEN28248 : _GEN28243;
wire  _GEN28250 = io_x[34] ? _GEN28249 : _GEN28239;
wire  _GEN28251 = io_x[39] ? _GEN28250 : _GEN28231;
wire  _GEN28252 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN28253 = io_x[38] ? _GEN28252 : _GEN21871;
wire  _GEN28254 = io_x[75] ? _GEN21772 : _GEN21758;
wire  _GEN28255 = io_x[38] ? _GEN28254 : _GEN21871;
wire  _GEN28256 = io_x[34] ? _GEN28255 : _GEN28253;
wire  _GEN28257 = io_x[39] ? _GEN21910 : _GEN28256;
wire  _GEN28258 = io_x[46] ? _GEN28257 : _GEN28251;
wire  _GEN28259 = io_x[18] ? _GEN28258 : _GEN28210;
wire  _GEN28260 = io_x[34] ? _GEN21766 : _GEN21927;
wire  _GEN28261 = io_x[39] ? _GEN22327 : _GEN28260;
wire  _GEN28262 = io_x[46] ? _GEN27726 : _GEN28261;
wire  _GEN28263 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28264 = io_x[27] ? _GEN28263 : _GEN21739;
wire  _GEN28265 = io_x[29] ? _GEN28264 : _GEN21743;
wire  _GEN28266 = io_x[75] ? _GEN28265 : _GEN21758;
wire  _GEN28267 = io_x[38] ? _GEN28266 : _GEN21833;
wire  _GEN28268 = io_x[34] ? _GEN28267 : _GEN21927;
wire  _GEN28269 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28270 = io_x[27] ? _GEN28269 : _GEN21739;
wire  _GEN28271 = io_x[29] ? _GEN28270 : _GEN21743;
wire  _GEN28272 = io_x[75] ? _GEN28271 : _GEN21772;
wire  _GEN28273 = io_x[38] ? _GEN21833 : _GEN28272;
wire  _GEN28274 = io_x[34] ? _GEN21927 : _GEN28273;
wire  _GEN28275 = io_x[39] ? _GEN28274 : _GEN28268;
wire  _GEN28276 = io_x[46] ? _GEN27726 : _GEN28275;
wire  _GEN28277 = io_x[18] ? _GEN28276 : _GEN28262;
wire  _GEN28278 = io_x[49] ? _GEN28277 : _GEN28259;
wire  _GEN28279 = io_x[24] ? _GEN28278 : _GEN28193;
wire  _GEN28280 = io_x[75] ? _GEN21758 : _GEN21772;
wire  _GEN28281 = io_x[38] ? _GEN21833 : _GEN28280;
wire  _GEN28282 = io_x[34] ? _GEN21927 : _GEN28281;
wire  _GEN28283 = io_x[39] ? _GEN21910 : _GEN28282;
wire  _GEN28284 = io_x[46] ? _GEN22145 : _GEN28283;
wire  _GEN28285 = io_x[29] ? _GEN21743 : _GEN21744;
wire  _GEN28286 = io_x[75] ? _GEN21758 : _GEN28285;
wire  _GEN28287 = io_x[38] ? _GEN28286 : _GEN21871;
wire  _GEN28288 = io_x[37] ? _GEN21735 : _GEN21734;
wire  _GEN28289 = io_x[27] ? _GEN28288 : _GEN21750;
wire  _GEN28290 = io_x[29] ? _GEN28289 : _GEN21743;
wire  _GEN28291 = io_x[75] ? _GEN21758 : _GEN28290;
wire  _GEN28292 = io_x[38] ? _GEN28291 : _GEN21833;
wire  _GEN28293 = io_x[34] ? _GEN28292 : _GEN28287;
wire  _GEN28294 = io_x[39] ? _GEN28293 : _GEN21910;
wire  _GEN28295 = io_x[46] ? _GEN22145 : _GEN28294;
wire  _GEN28296 = io_x[18] ? _GEN28295 : _GEN28284;
wire  _GEN28297 = io_x[49] ? _GEN22268 : _GEN28296;
wire  _GEN28298 = io_x[24] ? _GEN28297 : _GEN27801;
wire  _GEN28299 = io_x[80] ? _GEN28298 : _GEN28279;
wire  _GEN28300 = io_x[16] ? _GEN28299 : _GEN28159;
wire  _GEN28301 = io_x[22] ? _GEN28300 : _GEN28111;
wire  _GEN28302 = io_x[20] ? _GEN28301 : _GEN27957;
wire  _GEN28303 = io_x[33] ? _GEN28302 : _GEN27713;
assign io_y[1] = _GEN28303;
wire  _GEN28304 = 1'b0;
wire  _GEN28305 = 1'b1;
wire  _GEN28306 = io_x[34] ? _GEN28305 : _GEN28304;
wire  _GEN28307 = io_x[34] ? _GEN28305 : _GEN28304;
wire  _GEN28308 = io_x[38] ? _GEN28307 : _GEN28306;
wire  _GEN28309 = io_x[34] ? _GEN28305 : _GEN28304;
wire  _GEN28310 = io_x[34] ? _GEN28305 : _GEN28304;
wire  _GEN28311 = io_x[38] ? _GEN28310 : _GEN28309;
wire  _GEN28312 = io_x[44] ? _GEN28311 : _GEN28308;
wire  _GEN28313 = io_x[34] ? _GEN28305 : _GEN28304;
wire  _GEN28314 = io_x[34] ? _GEN28305 : _GEN28304;
wire  _GEN28315 = io_x[38] ? _GEN28314 : _GEN28313;
wire  _GEN28316 = io_x[34] ? _GEN28305 : _GEN28304;
wire  _GEN28317 = io_x[34] ? _GEN28305 : _GEN28304;
wire  _GEN28318 = io_x[38] ? _GEN28317 : _GEN28316;
wire  _GEN28319 = io_x[44] ? _GEN28318 : _GEN28315;
wire  _GEN28320 = io_x[4] ? _GEN28319 : _GEN28312;
assign io_y[0] = _GEN28320;
endmodule