module BBGSharePredictorImp_BSD_sim(
    input [31:0] pc,
    input [31:0] train_pc,
    input  train_taken,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    input [15:0] train_ghr_rdata,
    output  taken,
    output  pht_wdata,
    output [8:0] pht_raddr,
    output [8:0] pht_waddr,
    output  ghr_wdata
);
wire [98:0] io_x;
wire [20:0] io_y;
assign io_x = { pc, train_pc, train_taken, pht_rdata, ghr_rdata, train_ghr_rdata };
assign { taken, pht_wdata, pht_raddr, pht_waddr, ghr_wdata } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN3 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN4 = io_x[34] ? _GEN3 : _GEN2;
assign io_y[20] = _GEN4;
wire  _GEN5 = 1'b0;
wire  _GEN6 = 1'b1;
wire  _GEN7 = io_x[34] ? _GEN6 : _GEN5;
assign io_y[19] = _GEN7;
wire  _GEN8 = 1'b0;
wire  _GEN9 = 1'b1;
wire  _GEN10 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN11 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN12 = io_x[27] ? _GEN11 : _GEN10;
wire  _GEN13 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN14 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN15 = io_x[27] ? _GEN14 : _GEN13;
wire  _GEN16 = io_x[31] ? _GEN15 : _GEN12;
wire  _GEN17 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN18 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN19 = io_x[27] ? _GEN18 : _GEN17;
wire  _GEN20 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN21 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN22 = io_x[27] ? _GEN21 : _GEN20;
wire  _GEN23 = io_x[31] ? _GEN22 : _GEN19;
wire  _GEN24 = io_x[19] ? _GEN23 : _GEN16;
wire  _GEN25 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN26 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN27 = io_x[27] ? _GEN26 : _GEN25;
wire  _GEN28 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN29 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN30 = io_x[27] ? _GEN29 : _GEN28;
wire  _GEN31 = io_x[31] ? _GEN30 : _GEN27;
wire  _GEN32 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN33 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN34 = io_x[27] ? _GEN33 : _GEN32;
wire  _GEN35 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN36 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN37 = io_x[27] ? _GEN36 : _GEN35;
wire  _GEN38 = io_x[31] ? _GEN37 : _GEN34;
wire  _GEN39 = io_x[19] ? _GEN38 : _GEN31;
wire  _GEN40 = io_x[77] ? _GEN39 : _GEN24;
wire  _GEN41 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN42 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN43 = io_x[27] ? _GEN42 : _GEN41;
wire  _GEN44 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN45 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN46 = io_x[27] ? _GEN45 : _GEN44;
wire  _GEN47 = io_x[31] ? _GEN46 : _GEN43;
wire  _GEN48 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN49 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN50 = io_x[27] ? _GEN49 : _GEN48;
wire  _GEN51 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN52 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN53 = io_x[27] ? _GEN52 : _GEN51;
wire  _GEN54 = io_x[31] ? _GEN53 : _GEN50;
wire  _GEN55 = io_x[19] ? _GEN54 : _GEN47;
wire  _GEN56 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN57 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN58 = io_x[27] ? _GEN57 : _GEN56;
wire  _GEN59 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN60 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN61 = io_x[27] ? _GEN60 : _GEN59;
wire  _GEN62 = io_x[31] ? _GEN61 : _GEN58;
wire  _GEN63 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN64 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN65 = io_x[27] ? _GEN64 : _GEN63;
wire  _GEN66 = io_x[23] ? _GEN8 : _GEN9;
wire  _GEN67 = io_x[23] ? _GEN9 : _GEN8;
wire  _GEN68 = io_x[27] ? _GEN67 : _GEN66;
wire  _GEN69 = io_x[31] ? _GEN68 : _GEN65;
wire  _GEN70 = io_x[19] ? _GEN69 : _GEN62;
wire  _GEN71 = io_x[77] ? _GEN70 : _GEN55;
wire  _GEN72 = io_x[69] ? _GEN71 : _GEN40;
assign io_y[18] = _GEN72;
wire  _GEN73 = 1'b0;
wire  _GEN74 = 1'b1;
wire  _GEN75 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN76 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN77 = io_x[26] ? _GEN76 : _GEN75;
wire  _GEN78 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN79 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN80 = io_x[26] ? _GEN79 : _GEN78;
wire  _GEN81 = io_x[18] ? _GEN80 : _GEN77;
wire  _GEN82 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN83 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN84 = io_x[26] ? _GEN83 : _GEN82;
wire  _GEN85 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN86 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN87 = io_x[26] ? _GEN86 : _GEN85;
wire  _GEN88 = io_x[18] ? _GEN87 : _GEN84;
wire  _GEN89 = io_x[30] ? _GEN88 : _GEN81;
wire  _GEN90 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN91 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN92 = io_x[26] ? _GEN91 : _GEN90;
wire  _GEN93 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN94 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN95 = io_x[26] ? _GEN94 : _GEN93;
wire  _GEN96 = io_x[18] ? _GEN95 : _GEN92;
wire  _GEN97 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN98 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN99 = io_x[26] ? _GEN98 : _GEN97;
wire  _GEN100 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN101 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN102 = io_x[26] ? _GEN101 : _GEN100;
wire  _GEN103 = io_x[18] ? _GEN102 : _GEN99;
wire  _GEN104 = io_x[30] ? _GEN103 : _GEN96;
wire  _GEN105 = io_x[76] ? _GEN104 : _GEN89;
wire  _GEN106 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN107 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN108 = io_x[26] ? _GEN107 : _GEN106;
wire  _GEN109 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN110 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN111 = io_x[26] ? _GEN110 : _GEN109;
wire  _GEN112 = io_x[18] ? _GEN111 : _GEN108;
wire  _GEN113 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN114 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN115 = io_x[26] ? _GEN114 : _GEN113;
wire  _GEN116 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN117 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN118 = io_x[26] ? _GEN117 : _GEN116;
wire  _GEN119 = io_x[18] ? _GEN118 : _GEN115;
wire  _GEN120 = io_x[30] ? _GEN119 : _GEN112;
wire  _GEN121 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN122 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN123 = io_x[26] ? _GEN122 : _GEN121;
wire  _GEN124 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN125 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN126 = io_x[26] ? _GEN125 : _GEN124;
wire  _GEN127 = io_x[18] ? _GEN126 : _GEN123;
wire  _GEN128 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN129 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN130 = io_x[26] ? _GEN129 : _GEN128;
wire  _GEN131 = io_x[22] ? _GEN73 : _GEN74;
wire  _GEN132 = io_x[22] ? _GEN74 : _GEN73;
wire  _GEN133 = io_x[26] ? _GEN132 : _GEN131;
wire  _GEN134 = io_x[18] ? _GEN133 : _GEN130;
wire  _GEN135 = io_x[30] ? _GEN134 : _GEN127;
wire  _GEN136 = io_x[76] ? _GEN135 : _GEN120;
wire  _GEN137 = io_x[74] ? _GEN136 : _GEN105;
assign io_y[17] = _GEN137;
wire  _GEN138 = 1'b0;
wire  _GEN139 = 1'b1;
wire  _GEN140 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN141 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN142 = io_x[25] ? _GEN141 : _GEN140;
wire  _GEN143 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN144 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN145 = io_x[25] ? _GEN144 : _GEN143;
wire  _GEN146 = io_x[17] ? _GEN145 : _GEN142;
wire  _GEN147 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN148 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN149 = io_x[25] ? _GEN148 : _GEN147;
wire  _GEN150 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN151 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN152 = io_x[25] ? _GEN151 : _GEN150;
wire  _GEN153 = io_x[17] ? _GEN152 : _GEN149;
wire  _GEN154 = io_x[29] ? _GEN153 : _GEN146;
wire  _GEN155 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN156 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN157 = io_x[25] ? _GEN156 : _GEN155;
wire  _GEN158 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN159 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN160 = io_x[25] ? _GEN159 : _GEN158;
wire  _GEN161 = io_x[17] ? _GEN160 : _GEN157;
wire  _GEN162 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN163 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN164 = io_x[25] ? _GEN163 : _GEN162;
wire  _GEN165 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN166 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN167 = io_x[25] ? _GEN166 : _GEN165;
wire  _GEN168 = io_x[17] ? _GEN167 : _GEN164;
wire  _GEN169 = io_x[29] ? _GEN168 : _GEN161;
wire  _GEN170 = io_x[75] ? _GEN169 : _GEN154;
wire  _GEN171 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN172 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN173 = io_x[25] ? _GEN172 : _GEN171;
wire  _GEN174 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN175 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN176 = io_x[25] ? _GEN175 : _GEN174;
wire  _GEN177 = io_x[17] ? _GEN176 : _GEN173;
wire  _GEN178 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN179 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN180 = io_x[25] ? _GEN179 : _GEN178;
wire  _GEN181 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN182 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN183 = io_x[25] ? _GEN182 : _GEN181;
wire  _GEN184 = io_x[17] ? _GEN183 : _GEN180;
wire  _GEN185 = io_x[29] ? _GEN184 : _GEN177;
wire  _GEN186 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN187 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN188 = io_x[25] ? _GEN187 : _GEN186;
wire  _GEN189 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN190 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN191 = io_x[25] ? _GEN190 : _GEN189;
wire  _GEN192 = io_x[17] ? _GEN191 : _GEN188;
wire  _GEN193 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN194 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN195 = io_x[25] ? _GEN194 : _GEN193;
wire  _GEN196 = io_x[21] ? _GEN138 : _GEN139;
wire  _GEN197 = io_x[21] ? _GEN139 : _GEN138;
wire  _GEN198 = io_x[25] ? _GEN197 : _GEN196;
wire  _GEN199 = io_x[17] ? _GEN198 : _GEN195;
wire  _GEN200 = io_x[29] ? _GEN199 : _GEN192;
wire  _GEN201 = io_x[75] ? _GEN200 : _GEN185;
wire  _GEN202 = io_x[27] ? _GEN201 : _GEN170;
assign io_y[16] = _GEN202;
wire  _GEN203 = 1'b0;
wire  _GEN204 = 1'b1;
wire  _GEN205 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN206 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN207 = io_x[28] ? _GEN206 : _GEN205;
wire  _GEN208 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN209 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN210 = io_x[28] ? _GEN209 : _GEN208;
wire  _GEN211 = io_x[20] ? _GEN210 : _GEN207;
wire  _GEN212 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN213 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN214 = io_x[28] ? _GEN213 : _GEN212;
wire  _GEN215 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN216 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN217 = io_x[28] ? _GEN216 : _GEN215;
wire  _GEN218 = io_x[20] ? _GEN217 : _GEN214;
wire  _GEN219 = io_x[16] ? _GEN218 : _GEN211;
wire  _GEN220 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN221 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN222 = io_x[28] ? _GEN221 : _GEN220;
wire  _GEN223 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN224 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN225 = io_x[28] ? _GEN224 : _GEN223;
wire  _GEN226 = io_x[20] ? _GEN225 : _GEN222;
wire  _GEN227 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN228 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN229 = io_x[28] ? _GEN228 : _GEN227;
wire  _GEN230 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN231 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN232 = io_x[28] ? _GEN231 : _GEN230;
wire  _GEN233 = io_x[20] ? _GEN232 : _GEN229;
wire  _GEN234 = io_x[16] ? _GEN233 : _GEN226;
wire  _GEN235 = io_x[74] ? _GEN234 : _GEN219;
wire  _GEN236 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN237 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN238 = io_x[28] ? _GEN237 : _GEN236;
wire  _GEN239 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN240 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN241 = io_x[28] ? _GEN240 : _GEN239;
wire  _GEN242 = io_x[20] ? _GEN241 : _GEN238;
wire  _GEN243 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN244 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN245 = io_x[28] ? _GEN244 : _GEN243;
wire  _GEN246 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN247 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN248 = io_x[28] ? _GEN247 : _GEN246;
wire  _GEN249 = io_x[20] ? _GEN248 : _GEN245;
wire  _GEN250 = io_x[16] ? _GEN249 : _GEN242;
wire  _GEN251 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN252 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN253 = io_x[28] ? _GEN252 : _GEN251;
wire  _GEN254 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN255 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN256 = io_x[28] ? _GEN255 : _GEN254;
wire  _GEN257 = io_x[20] ? _GEN256 : _GEN253;
wire  _GEN258 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN259 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN260 = io_x[28] ? _GEN259 : _GEN258;
wire  _GEN261 = io_x[24] ? _GEN203 : _GEN204;
wire  _GEN262 = io_x[24] ? _GEN204 : _GEN203;
wire  _GEN263 = io_x[28] ? _GEN262 : _GEN261;
wire  _GEN264 = io_x[20] ? _GEN263 : _GEN260;
wire  _GEN265 = io_x[16] ? _GEN264 : _GEN257;
wire  _GEN266 = io_x[74] ? _GEN265 : _GEN250;
wire  _GEN267 = io_x[72] ? _GEN266 : _GEN235;
assign io_y[15] = _GEN267;
wire  _GEN268 = 1'b0;
wire  _GEN269 = 1'b1;
wire  _GEN270 = io_x[73] ? _GEN269 : _GEN268;
wire  _GEN271 = io_x[73] ? _GEN269 : _GEN268;
wire  _GEN272 = io_x[69] ? _GEN271 : _GEN270;
assign io_y[14] = _GEN272;
wire  _GEN273 = 1'b0;
wire  _GEN274 = 1'b1;
wire  _GEN275 = io_x[72] ? _GEN274 : _GEN273;
wire  _GEN276 = io_x[72] ? _GEN274 : _GEN273;
wire  _GEN277 = io_x[78] ? _GEN276 : _GEN275;
assign io_y[13] = _GEN277;
wire  _GEN278 = 1'b0;
wire  _GEN279 = 1'b1;
wire  _GEN280 = io_x[71] ? _GEN279 : _GEN278;
assign io_y[12] = _GEN280;
wire  _GEN281 = 1'b0;
wire  _GEN282 = 1'b1;
wire  _GEN283 = io_x[70] ? _GEN282 : _GEN281;
wire  _GEN284 = io_x[70] ? _GEN282 : _GEN281;
wire  _GEN285 = io_x[73] ? _GEN284 : _GEN283;
wire  _GEN286 = io_x[70] ? _GEN282 : _GEN281;
wire  _GEN287 = io_x[70] ? _GEN282 : _GEN281;
wire  _GEN288 = io_x[73] ? _GEN287 : _GEN286;
wire  _GEN289 = io_x[74] ? _GEN288 : _GEN285;
assign io_y[11] = _GEN289;
wire  _GEN290 = 1'b0;
wire  _GEN291 = 1'b1;
wire  _GEN292 = io_x[69] ? _GEN291 : _GEN290;
wire  _GEN293 = io_x[69] ? _GEN291 : _GEN290;
wire  _GEN294 = io_x[73] ? _GEN293 : _GEN292;
wire  _GEN295 = io_x[69] ? _GEN291 : _GEN290;
wire  _GEN296 = io_x[69] ? _GEN291 : _GEN290;
wire  _GEN297 = io_x[73] ? _GEN296 : _GEN295;
wire  _GEN298 = io_x[78] ? _GEN297 : _GEN294;
assign io_y[10] = _GEN298;
wire  _GEN299 = 1'b0;
wire  _GEN300 = 1'b1;
wire  _GEN301 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN302 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN303 = io_x[27] ? _GEN302 : _GEN301;
wire  _GEN304 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN305 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN306 = io_x[27] ? _GEN305 : _GEN304;
wire  _GEN307 = io_x[31] ? _GEN306 : _GEN303;
wire  _GEN308 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN309 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN310 = io_x[27] ? _GEN309 : _GEN308;
wire  _GEN311 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN312 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN313 = io_x[27] ? _GEN312 : _GEN311;
wire  _GEN314 = io_x[31] ? _GEN313 : _GEN310;
wire  _GEN315 = io_x[19] ? _GEN314 : _GEN307;
wire  _GEN316 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN317 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN318 = io_x[27] ? _GEN317 : _GEN316;
wire  _GEN319 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN320 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN321 = io_x[27] ? _GEN320 : _GEN319;
wire  _GEN322 = io_x[31] ? _GEN321 : _GEN318;
wire  _GEN323 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN324 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN325 = io_x[27] ? _GEN324 : _GEN323;
wire  _GEN326 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN327 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN328 = io_x[27] ? _GEN327 : _GEN326;
wire  _GEN329 = io_x[31] ? _GEN328 : _GEN325;
wire  _GEN330 = io_x[19] ? _GEN329 : _GEN322;
wire  _GEN331 = io_x[77] ? _GEN330 : _GEN315;
wire  _GEN332 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN333 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN334 = io_x[27] ? _GEN333 : _GEN332;
wire  _GEN335 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN336 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN337 = io_x[27] ? _GEN336 : _GEN335;
wire  _GEN338 = io_x[31] ? _GEN337 : _GEN334;
wire  _GEN339 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN340 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN341 = io_x[27] ? _GEN340 : _GEN339;
wire  _GEN342 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN343 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN344 = io_x[27] ? _GEN343 : _GEN342;
wire  _GEN345 = io_x[31] ? _GEN344 : _GEN341;
wire  _GEN346 = io_x[19] ? _GEN345 : _GEN338;
wire  _GEN347 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN348 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN349 = io_x[27] ? _GEN348 : _GEN347;
wire  _GEN350 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN351 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN352 = io_x[27] ? _GEN351 : _GEN350;
wire  _GEN353 = io_x[31] ? _GEN352 : _GEN349;
wire  _GEN354 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN355 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN356 = io_x[27] ? _GEN355 : _GEN354;
wire  _GEN357 = io_x[23] ? _GEN299 : _GEN300;
wire  _GEN358 = io_x[23] ? _GEN300 : _GEN299;
wire  _GEN359 = io_x[27] ? _GEN358 : _GEN357;
wire  _GEN360 = io_x[31] ? _GEN359 : _GEN356;
wire  _GEN361 = io_x[19] ? _GEN360 : _GEN353;
wire  _GEN362 = io_x[77] ? _GEN361 : _GEN346;
wire  _GEN363 = io_x[69] ? _GEN362 : _GEN331;
assign io_y[9] = _GEN363;
wire  _GEN364 = 1'b0;
wire  _GEN365 = 1'b1;
wire  _GEN366 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN367 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN368 = io_x[26] ? _GEN367 : _GEN366;
wire  _GEN369 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN370 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN371 = io_x[26] ? _GEN370 : _GEN369;
wire  _GEN372 = io_x[18] ? _GEN371 : _GEN368;
wire  _GEN373 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN374 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN375 = io_x[26] ? _GEN374 : _GEN373;
wire  _GEN376 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN377 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN378 = io_x[26] ? _GEN377 : _GEN376;
wire  _GEN379 = io_x[18] ? _GEN378 : _GEN375;
wire  _GEN380 = io_x[30] ? _GEN379 : _GEN372;
wire  _GEN381 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN382 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN383 = io_x[26] ? _GEN382 : _GEN381;
wire  _GEN384 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN385 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN386 = io_x[26] ? _GEN385 : _GEN384;
wire  _GEN387 = io_x[18] ? _GEN386 : _GEN383;
wire  _GEN388 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN389 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN390 = io_x[26] ? _GEN389 : _GEN388;
wire  _GEN391 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN392 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN393 = io_x[26] ? _GEN392 : _GEN391;
wire  _GEN394 = io_x[18] ? _GEN393 : _GEN390;
wire  _GEN395 = io_x[30] ? _GEN394 : _GEN387;
wire  _GEN396 = io_x[76] ? _GEN395 : _GEN380;
wire  _GEN397 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN398 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN399 = io_x[26] ? _GEN398 : _GEN397;
wire  _GEN400 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN401 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN402 = io_x[26] ? _GEN401 : _GEN400;
wire  _GEN403 = io_x[18] ? _GEN402 : _GEN399;
wire  _GEN404 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN405 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN406 = io_x[26] ? _GEN405 : _GEN404;
wire  _GEN407 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN408 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN409 = io_x[26] ? _GEN408 : _GEN407;
wire  _GEN410 = io_x[18] ? _GEN409 : _GEN406;
wire  _GEN411 = io_x[30] ? _GEN410 : _GEN403;
wire  _GEN412 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN413 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN414 = io_x[26] ? _GEN413 : _GEN412;
wire  _GEN415 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN416 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN417 = io_x[26] ? _GEN416 : _GEN415;
wire  _GEN418 = io_x[18] ? _GEN417 : _GEN414;
wire  _GEN419 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN420 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN421 = io_x[26] ? _GEN420 : _GEN419;
wire  _GEN422 = io_x[22] ? _GEN364 : _GEN365;
wire  _GEN423 = io_x[22] ? _GEN365 : _GEN364;
wire  _GEN424 = io_x[26] ? _GEN423 : _GEN422;
wire  _GEN425 = io_x[18] ? _GEN424 : _GEN421;
wire  _GEN426 = io_x[30] ? _GEN425 : _GEN418;
wire  _GEN427 = io_x[76] ? _GEN426 : _GEN411;
wire  _GEN428 = io_x[74] ? _GEN427 : _GEN396;
assign io_y[8] = _GEN428;
wire  _GEN429 = 1'b0;
wire  _GEN430 = 1'b1;
wire  _GEN431 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN432 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN433 = io_x[25] ? _GEN432 : _GEN431;
wire  _GEN434 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN435 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN436 = io_x[25] ? _GEN435 : _GEN434;
wire  _GEN437 = io_x[17] ? _GEN436 : _GEN433;
wire  _GEN438 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN439 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN440 = io_x[25] ? _GEN439 : _GEN438;
wire  _GEN441 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN442 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN443 = io_x[25] ? _GEN442 : _GEN441;
wire  _GEN444 = io_x[17] ? _GEN443 : _GEN440;
wire  _GEN445 = io_x[29] ? _GEN444 : _GEN437;
wire  _GEN446 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN447 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN448 = io_x[25] ? _GEN447 : _GEN446;
wire  _GEN449 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN450 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN451 = io_x[25] ? _GEN450 : _GEN449;
wire  _GEN452 = io_x[17] ? _GEN451 : _GEN448;
wire  _GEN453 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN454 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN455 = io_x[25] ? _GEN454 : _GEN453;
wire  _GEN456 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN457 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN458 = io_x[25] ? _GEN457 : _GEN456;
wire  _GEN459 = io_x[17] ? _GEN458 : _GEN455;
wire  _GEN460 = io_x[29] ? _GEN459 : _GEN452;
wire  _GEN461 = io_x[75] ? _GEN460 : _GEN445;
wire  _GEN462 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN463 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN464 = io_x[25] ? _GEN463 : _GEN462;
wire  _GEN465 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN466 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN467 = io_x[25] ? _GEN466 : _GEN465;
wire  _GEN468 = io_x[17] ? _GEN467 : _GEN464;
wire  _GEN469 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN470 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN471 = io_x[25] ? _GEN470 : _GEN469;
wire  _GEN472 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN473 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN474 = io_x[25] ? _GEN473 : _GEN472;
wire  _GEN475 = io_x[17] ? _GEN474 : _GEN471;
wire  _GEN476 = io_x[29] ? _GEN475 : _GEN468;
wire  _GEN477 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN478 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN479 = io_x[25] ? _GEN478 : _GEN477;
wire  _GEN480 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN481 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN482 = io_x[25] ? _GEN481 : _GEN480;
wire  _GEN483 = io_x[17] ? _GEN482 : _GEN479;
wire  _GEN484 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN485 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN486 = io_x[25] ? _GEN485 : _GEN484;
wire  _GEN487 = io_x[21] ? _GEN429 : _GEN430;
wire  _GEN488 = io_x[21] ? _GEN430 : _GEN429;
wire  _GEN489 = io_x[25] ? _GEN488 : _GEN487;
wire  _GEN490 = io_x[17] ? _GEN489 : _GEN486;
wire  _GEN491 = io_x[29] ? _GEN490 : _GEN483;
wire  _GEN492 = io_x[75] ? _GEN491 : _GEN476;
wire  _GEN493 = io_x[27] ? _GEN492 : _GEN461;
assign io_y[7] = _GEN493;
wire  _GEN494 = 1'b0;
wire  _GEN495 = 1'b1;
wire  _GEN496 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN497 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN498 = io_x[28] ? _GEN497 : _GEN496;
wire  _GEN499 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN500 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN501 = io_x[28] ? _GEN500 : _GEN499;
wire  _GEN502 = io_x[20] ? _GEN501 : _GEN498;
wire  _GEN503 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN504 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN505 = io_x[28] ? _GEN504 : _GEN503;
wire  _GEN506 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN507 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN508 = io_x[28] ? _GEN507 : _GEN506;
wire  _GEN509 = io_x[20] ? _GEN508 : _GEN505;
wire  _GEN510 = io_x[16] ? _GEN509 : _GEN502;
wire  _GEN511 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN512 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN513 = io_x[28] ? _GEN512 : _GEN511;
wire  _GEN514 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN515 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN516 = io_x[28] ? _GEN515 : _GEN514;
wire  _GEN517 = io_x[20] ? _GEN516 : _GEN513;
wire  _GEN518 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN519 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN520 = io_x[28] ? _GEN519 : _GEN518;
wire  _GEN521 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN522 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN523 = io_x[28] ? _GEN522 : _GEN521;
wire  _GEN524 = io_x[20] ? _GEN523 : _GEN520;
wire  _GEN525 = io_x[16] ? _GEN524 : _GEN517;
wire  _GEN526 = io_x[74] ? _GEN525 : _GEN510;
wire  _GEN527 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN528 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN529 = io_x[28] ? _GEN528 : _GEN527;
wire  _GEN530 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN531 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN532 = io_x[28] ? _GEN531 : _GEN530;
wire  _GEN533 = io_x[20] ? _GEN532 : _GEN529;
wire  _GEN534 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN535 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN536 = io_x[28] ? _GEN535 : _GEN534;
wire  _GEN537 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN538 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN539 = io_x[28] ? _GEN538 : _GEN537;
wire  _GEN540 = io_x[20] ? _GEN539 : _GEN536;
wire  _GEN541 = io_x[16] ? _GEN540 : _GEN533;
wire  _GEN542 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN543 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN544 = io_x[28] ? _GEN543 : _GEN542;
wire  _GEN545 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN546 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN547 = io_x[28] ? _GEN546 : _GEN545;
wire  _GEN548 = io_x[20] ? _GEN547 : _GEN544;
wire  _GEN549 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN550 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN551 = io_x[28] ? _GEN550 : _GEN549;
wire  _GEN552 = io_x[24] ? _GEN494 : _GEN495;
wire  _GEN553 = io_x[24] ? _GEN495 : _GEN494;
wire  _GEN554 = io_x[28] ? _GEN553 : _GEN552;
wire  _GEN555 = io_x[20] ? _GEN554 : _GEN551;
wire  _GEN556 = io_x[16] ? _GEN555 : _GEN548;
wire  _GEN557 = io_x[74] ? _GEN556 : _GEN541;
wire  _GEN558 = io_x[72] ? _GEN557 : _GEN526;
assign io_y[6] = _GEN558;
wire  _GEN559 = 1'b0;
wire  _GEN560 = 1'b1;
wire  _GEN561 = io_x[73] ? _GEN560 : _GEN559;
wire  _GEN562 = io_x[73] ? _GEN560 : _GEN559;
wire  _GEN563 = io_x[69] ? _GEN562 : _GEN561;
assign io_y[5] = _GEN563;
wire  _GEN564 = 1'b0;
wire  _GEN565 = 1'b1;
wire  _GEN566 = io_x[72] ? _GEN565 : _GEN564;
wire  _GEN567 = io_x[72] ? _GEN565 : _GEN564;
wire  _GEN568 = io_x[78] ? _GEN567 : _GEN566;
assign io_y[4] = _GEN568;
wire  _GEN569 = 1'b0;
wire  _GEN570 = 1'b1;
wire  _GEN571 = io_x[71] ? _GEN570 : _GEN569;
assign io_y[3] = _GEN571;
wire  _GEN572 = 1'b0;
wire  _GEN573 = 1'b1;
wire  _GEN574 = io_x[70] ? _GEN573 : _GEN572;
wire  _GEN575 = io_x[70] ? _GEN573 : _GEN572;
wire  _GEN576 = io_x[73] ? _GEN575 : _GEN574;
wire  _GEN577 = io_x[70] ? _GEN573 : _GEN572;
wire  _GEN578 = io_x[70] ? _GEN573 : _GEN572;
wire  _GEN579 = io_x[73] ? _GEN578 : _GEN577;
wire  _GEN580 = io_x[74] ? _GEN579 : _GEN576;
assign io_y[2] = _GEN580;
wire  _GEN581 = 1'b0;
wire  _GEN582 = 1'b1;
wire  _GEN583 = io_x[69] ? _GEN582 : _GEN581;
wire  _GEN584 = io_x[69] ? _GEN582 : _GEN581;
wire  _GEN585 = io_x[73] ? _GEN584 : _GEN583;
wire  _GEN586 = io_x[69] ? _GEN582 : _GEN581;
wire  _GEN587 = io_x[69] ? _GEN582 : _GEN581;
wire  _GEN588 = io_x[73] ? _GEN587 : _GEN586;
wire  _GEN589 = io_x[78] ? _GEN588 : _GEN585;
assign io_y[1] = _GEN589;
wire  _GEN590 = 1'b0;
wire  _GEN591 = 1'b1;
wire  _GEN592 = io_x[34] ? _GEN591 : _GEN590;
assign io_y[0] = _GEN592;
endmodule
