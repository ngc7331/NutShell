module BBGSharePredictorImp_BSD_b_NutShell_split(
    input [31:0] pc,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    output  taken,
    output [8:0] pht_raddr,
    input [31:0] train_pc,
    input  train_taken,
    input [15:0] train_ghr_rdata,
    output  pht_wdata,
    output [8:0] pht_waddr,
    output  ghr_wdata
);

BBGSharePredictorImp_BSD_NutShell_pred _pred(
    .pc        (pc),
    .pht_rdata (pht_rdata),
    .ghr_rdata (ghr_rdata),
    .taken     (taken),
    .pht_raddr (pht_raddr)
);

BBGSharePredictorImp_BSD_NutShell_train _train(
    .train_pc        (train_pc),
    .train_taken     (train_taken),
    .train_ghr_rdata (train_ghr_rdata),
    .pht_wdata       (pht_wdata),
    .pht_waddr       (pht_waddr),
    .ghr_wdata       (ghr_wdata)
);
endmodule
module BBGSharePredictorImp_BSD_NutShell_pred(
    input [31:0] pc,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    output  taken,
    output [8:0] pht_raddr
);
wire [49:0] io_x;
wire [9:0] io_y;
assign io_x = { pc, pht_rdata, ghr_rdata };
assign { taken, pht_raddr } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN3 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN4 = io_x[16] ? _GEN3 : _GEN2;
wire  _GEN5 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN6 = io_x[17] ? _GEN1 : _GEN0;
wire  _GEN7 = io_x[16] ? _GEN6 : _GEN5;
wire  _GEN8 = io_x[2] ? _GEN7 : _GEN4;
assign io_y[9] = _GEN8;
wire  _GEN9 = 1'b0;
wire  _GEN10 = 1'b1;
wire  _GEN11 = io_x[28] ? _GEN10 : _GEN9;
wire  _GEN12 = io_x[28] ? _GEN9 : _GEN10;
wire  _GEN13 = io_x[15] ? _GEN12 : _GEN11;
wire  _GEN14 = io_x[28] ? _GEN9 : _GEN10;
wire  _GEN15 = io_x[28] ? _GEN10 : _GEN9;
wire  _GEN16 = io_x[15] ? _GEN15 : _GEN14;
wire  _GEN17 = io_x[7] ? _GEN16 : _GEN13;
wire  _GEN18 = io_x[28] ? _GEN9 : _GEN10;
wire  _GEN19 = io_x[28] ? _GEN10 : _GEN9;
wire  _GEN20 = io_x[15] ? _GEN19 : _GEN18;
wire  _GEN21 = io_x[28] ? _GEN10 : _GEN9;
wire  _GEN22 = io_x[28] ? _GEN9 : _GEN10;
wire  _GEN23 = io_x[15] ? _GEN22 : _GEN21;
wire  _GEN24 = io_x[7] ? _GEN23 : _GEN20;
wire  _GEN25 = io_x[11] ? _GEN24 : _GEN17;
wire  _GEN26 = io_x[28] ? _GEN9 : _GEN10;
wire  _GEN27 = io_x[28] ? _GEN10 : _GEN9;
wire  _GEN28 = io_x[15] ? _GEN27 : _GEN26;
wire  _GEN29 = io_x[28] ? _GEN10 : _GEN9;
wire  _GEN30 = io_x[28] ? _GEN9 : _GEN10;
wire  _GEN31 = io_x[15] ? _GEN30 : _GEN29;
wire  _GEN32 = io_x[7] ? _GEN31 : _GEN28;
wire  _GEN33 = io_x[28] ? _GEN10 : _GEN9;
wire  _GEN34 = io_x[28] ? _GEN9 : _GEN10;
wire  _GEN35 = io_x[15] ? _GEN34 : _GEN33;
wire  _GEN36 = io_x[28] ? _GEN9 : _GEN10;
wire  _GEN37 = io_x[28] ? _GEN10 : _GEN9;
wire  _GEN38 = io_x[15] ? _GEN37 : _GEN36;
wire  _GEN39 = io_x[7] ? _GEN38 : _GEN35;
wire  _GEN40 = io_x[11] ? _GEN39 : _GEN32;
wire  _GEN41 = io_x[3] ? _GEN40 : _GEN25;
assign io_y[8] = _GEN41;
wire  _GEN42 = 1'b0;
wire  _GEN43 = 1'b1;
wire  _GEN44 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN45 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN46 = io_x[6] ? _GEN45 : _GEN44;
wire  _GEN47 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN48 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN49 = io_x[6] ? _GEN48 : _GEN47;
wire  _GEN50 = io_x[2] ? _GEN49 : _GEN46;
wire  _GEN51 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN52 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN53 = io_x[6] ? _GEN52 : _GEN51;
wire  _GEN54 = 1'b1;
wire  _GEN55 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN56 = io_x[6] ? _GEN55 : _GEN54;
wire  _GEN57 = io_x[2] ? _GEN56 : _GEN53;
wire  _GEN58 = io_x[14] ? _GEN57 : _GEN50;
wire  _GEN59 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN60 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN61 = io_x[6] ? _GEN60 : _GEN59;
wire  _GEN62 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN63 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN64 = io_x[6] ? _GEN63 : _GEN62;
wire  _GEN65 = io_x[2] ? _GEN64 : _GEN61;
wire  _GEN66 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN67 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN68 = io_x[6] ? _GEN67 : _GEN66;
wire  _GEN69 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN70 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN71 = io_x[6] ? _GEN70 : _GEN69;
wire  _GEN72 = io_x[2] ? _GEN71 : _GEN68;
wire  _GEN73 = io_x[14] ? _GEN72 : _GEN65;
wire  _GEN74 = io_x[10] ? _GEN73 : _GEN58;
wire  _GEN75 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN76 = io_x[6] ? _GEN75 : _GEN54;
wire  _GEN77 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN78 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN79 = io_x[6] ? _GEN78 : _GEN77;
wire  _GEN80 = io_x[2] ? _GEN79 : _GEN76;
wire  _GEN81 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN82 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN83 = io_x[6] ? _GEN82 : _GEN81;
wire  _GEN84 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN85 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN86 = io_x[6] ? _GEN85 : _GEN84;
wire  _GEN87 = io_x[2] ? _GEN86 : _GEN83;
wire  _GEN88 = io_x[14] ? _GEN87 : _GEN80;
wire  _GEN89 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN90 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN91 = io_x[6] ? _GEN90 : _GEN89;
wire  _GEN92 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN93 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN94 = io_x[6] ? _GEN93 : _GEN92;
wire  _GEN95 = io_x[2] ? _GEN94 : _GEN91;
wire  _GEN96 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN97 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN98 = io_x[6] ? _GEN97 : _GEN96;
wire  _GEN99 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN100 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN101 = io_x[6] ? _GEN100 : _GEN99;
wire  _GEN102 = io_x[2] ? _GEN101 : _GEN98;
wire  _GEN103 = io_x[14] ? _GEN102 : _GEN95;
wire  _GEN104 = io_x[10] ? _GEN103 : _GEN88;
wire  _GEN105 = io_x[17] ? _GEN104 : _GEN74;
wire  _GEN106 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN107 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN108 = io_x[6] ? _GEN107 : _GEN106;
wire  _GEN109 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN110 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN111 = io_x[6] ? _GEN110 : _GEN109;
wire  _GEN112 = io_x[2] ? _GEN111 : _GEN108;
wire  _GEN113 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN114 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN115 = io_x[6] ? _GEN114 : _GEN113;
wire  _GEN116 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN117 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN118 = io_x[6] ? _GEN117 : _GEN116;
wire  _GEN119 = io_x[2] ? _GEN118 : _GEN115;
wire  _GEN120 = io_x[14] ? _GEN119 : _GEN112;
wire  _GEN121 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN122 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN123 = io_x[6] ? _GEN122 : _GEN121;
wire  _GEN124 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN125 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN126 = io_x[6] ? _GEN125 : _GEN124;
wire  _GEN127 = io_x[2] ? _GEN126 : _GEN123;
wire  _GEN128 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN129 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN130 = io_x[6] ? _GEN129 : _GEN128;
wire  _GEN131 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN132 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN133 = io_x[6] ? _GEN132 : _GEN131;
wire  _GEN134 = io_x[2] ? _GEN133 : _GEN130;
wire  _GEN135 = io_x[14] ? _GEN134 : _GEN127;
wire  _GEN136 = io_x[10] ? _GEN135 : _GEN120;
wire  _GEN137 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN138 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN139 = io_x[6] ? _GEN138 : _GEN137;
wire  _GEN140 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN141 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN142 = io_x[6] ? _GEN141 : _GEN140;
wire  _GEN143 = io_x[2] ? _GEN142 : _GEN139;
wire  _GEN144 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN145 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN146 = io_x[6] ? _GEN145 : _GEN144;
wire  _GEN147 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN148 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN149 = io_x[6] ? _GEN148 : _GEN147;
wire  _GEN150 = io_x[2] ? _GEN149 : _GEN146;
wire  _GEN151 = io_x[14] ? _GEN150 : _GEN143;
wire  _GEN152 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN153 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN154 = io_x[6] ? _GEN153 : _GEN152;
wire  _GEN155 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN156 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN157 = io_x[6] ? _GEN156 : _GEN155;
wire  _GEN158 = io_x[2] ? _GEN157 : _GEN154;
wire  _GEN159 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN160 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN161 = io_x[6] ? _GEN160 : _GEN159;
wire  _GEN162 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN163 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN164 = io_x[6] ? _GEN163 : _GEN162;
wire  _GEN165 = io_x[2] ? _GEN164 : _GEN161;
wire  _GEN166 = io_x[14] ? _GEN165 : _GEN158;
wire  _GEN167 = io_x[10] ? _GEN166 : _GEN151;
wire  _GEN168 = io_x[17] ? _GEN167 : _GEN136;
wire  _GEN169 = io_x[25] ? _GEN168 : _GEN105;
wire  _GEN170 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN171 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN172 = io_x[6] ? _GEN171 : _GEN170;
wire  _GEN173 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN174 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN175 = io_x[6] ? _GEN174 : _GEN173;
wire  _GEN176 = io_x[2] ? _GEN175 : _GEN172;
wire  _GEN177 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN178 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN179 = io_x[6] ? _GEN178 : _GEN177;
wire  _GEN180 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN181 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN182 = io_x[6] ? _GEN181 : _GEN180;
wire  _GEN183 = io_x[2] ? _GEN182 : _GEN179;
wire  _GEN184 = io_x[14] ? _GEN183 : _GEN176;
wire  _GEN185 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN186 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN187 = io_x[6] ? _GEN186 : _GEN185;
wire  _GEN188 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN189 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN190 = io_x[6] ? _GEN189 : _GEN188;
wire  _GEN191 = io_x[2] ? _GEN190 : _GEN187;
wire  _GEN192 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN193 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN194 = io_x[6] ? _GEN193 : _GEN192;
wire  _GEN195 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN196 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN197 = io_x[6] ? _GEN196 : _GEN195;
wire  _GEN198 = io_x[2] ? _GEN197 : _GEN194;
wire  _GEN199 = io_x[14] ? _GEN198 : _GEN191;
wire  _GEN200 = io_x[10] ? _GEN199 : _GEN184;
wire  _GEN201 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN202 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN203 = io_x[6] ? _GEN202 : _GEN201;
wire  _GEN204 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN205 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN206 = io_x[6] ? _GEN205 : _GEN204;
wire  _GEN207 = io_x[2] ? _GEN206 : _GEN203;
wire  _GEN208 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN209 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN210 = io_x[6] ? _GEN209 : _GEN208;
wire  _GEN211 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN212 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN213 = io_x[6] ? _GEN212 : _GEN211;
wire  _GEN214 = io_x[2] ? _GEN213 : _GEN210;
wire  _GEN215 = io_x[14] ? _GEN214 : _GEN207;
wire  _GEN216 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN217 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN218 = io_x[6] ? _GEN217 : _GEN216;
wire  _GEN219 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN220 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN221 = io_x[6] ? _GEN220 : _GEN219;
wire  _GEN222 = io_x[2] ? _GEN221 : _GEN218;
wire  _GEN223 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN224 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN225 = io_x[6] ? _GEN224 : _GEN223;
wire  _GEN226 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN227 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN228 = io_x[6] ? _GEN227 : _GEN226;
wire  _GEN229 = io_x[2] ? _GEN228 : _GEN225;
wire  _GEN230 = io_x[14] ? _GEN229 : _GEN222;
wire  _GEN231 = io_x[10] ? _GEN230 : _GEN215;
wire  _GEN232 = io_x[17] ? _GEN231 : _GEN200;
wire  _GEN233 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN234 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN235 = io_x[6] ? _GEN234 : _GEN233;
wire  _GEN236 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN237 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN238 = io_x[6] ? _GEN237 : _GEN236;
wire  _GEN239 = io_x[2] ? _GEN238 : _GEN235;
wire  _GEN240 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN241 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN242 = io_x[6] ? _GEN241 : _GEN240;
wire  _GEN243 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN244 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN245 = io_x[6] ? _GEN244 : _GEN243;
wire  _GEN246 = io_x[2] ? _GEN245 : _GEN242;
wire  _GEN247 = io_x[14] ? _GEN246 : _GEN239;
wire  _GEN248 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN249 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN250 = io_x[6] ? _GEN249 : _GEN248;
wire  _GEN251 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN252 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN253 = io_x[6] ? _GEN252 : _GEN251;
wire  _GEN254 = io_x[2] ? _GEN253 : _GEN250;
wire  _GEN255 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN256 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN257 = io_x[6] ? _GEN256 : _GEN255;
wire  _GEN258 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN259 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN260 = io_x[6] ? _GEN259 : _GEN258;
wire  _GEN261 = io_x[2] ? _GEN260 : _GEN257;
wire  _GEN262 = io_x[14] ? _GEN261 : _GEN254;
wire  _GEN263 = io_x[10] ? _GEN262 : _GEN247;
wire  _GEN264 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN265 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN266 = io_x[6] ? _GEN265 : _GEN264;
wire  _GEN267 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN268 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN269 = io_x[6] ? _GEN268 : _GEN267;
wire  _GEN270 = io_x[2] ? _GEN269 : _GEN266;
wire  _GEN271 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN272 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN273 = io_x[6] ? _GEN272 : _GEN271;
wire  _GEN274 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN275 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN276 = io_x[6] ? _GEN275 : _GEN274;
wire  _GEN277 = io_x[2] ? _GEN276 : _GEN273;
wire  _GEN278 = io_x[14] ? _GEN277 : _GEN270;
wire  _GEN279 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN280 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN281 = io_x[6] ? _GEN280 : _GEN279;
wire  _GEN282 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN283 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN284 = io_x[6] ? _GEN283 : _GEN282;
wire  _GEN285 = io_x[2] ? _GEN284 : _GEN281;
wire  _GEN286 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN287 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN288 = io_x[6] ? _GEN287 : _GEN286;
wire  _GEN289 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN290 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN291 = io_x[6] ? _GEN290 : _GEN289;
wire  _GEN292 = io_x[2] ? _GEN291 : _GEN288;
wire  _GEN293 = io_x[14] ? _GEN292 : _GEN285;
wire  _GEN294 = io_x[10] ? _GEN293 : _GEN278;
wire  _GEN295 = io_x[17] ? _GEN294 : _GEN263;
wire  _GEN296 = io_x[25] ? _GEN295 : _GEN232;
wire  _GEN297 = io_x[24] ? _GEN296 : _GEN169;
wire  _GEN298 = 1'b0;
wire  _GEN299 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN300 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN301 = io_x[6] ? _GEN300 : _GEN298;
wire  _GEN302 = io_x[2] ? _GEN301 : _GEN299;
wire  _GEN303 = 1'b1;
wire  _GEN304 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN305 = io_x[6] ? _GEN304 : _GEN54;
wire  _GEN306 = io_x[2] ? _GEN305 : _GEN303;
wire  _GEN307 = io_x[14] ? _GEN306 : _GEN302;
wire  _GEN308 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN309 = io_x[6] ? _GEN308 : _GEN298;
wire  _GEN310 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN311 = io_x[6] ? _GEN310 : _GEN54;
wire  _GEN312 = io_x[2] ? _GEN311 : _GEN309;
wire  _GEN313 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN314 = io_x[6] ? _GEN313 : _GEN54;
wire  _GEN315 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN316 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN317 = io_x[6] ? _GEN316 : _GEN315;
wire  _GEN318 = io_x[2] ? _GEN317 : _GEN314;
wire  _GEN319 = io_x[14] ? _GEN318 : _GEN312;
wire  _GEN320 = io_x[10] ? _GEN319 : _GEN307;
wire  _GEN321 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN322 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN323 = io_x[6] ? _GEN322 : _GEN298;
wire  _GEN324 = io_x[2] ? _GEN323 : _GEN321;
wire  _GEN325 = io_x[6] ? _GEN54 : _GEN298;
wire  _GEN326 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN327 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN328 = io_x[6] ? _GEN327 : _GEN326;
wire  _GEN329 = io_x[2] ? _GEN328 : _GEN325;
wire  _GEN330 = io_x[14] ? _GEN329 : _GEN324;
wire  _GEN331 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN332 = io_x[6] ? _GEN331 : _GEN298;
wire  _GEN333 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN334 = io_x[6] ? _GEN333 : _GEN54;
wire  _GEN335 = io_x[2] ? _GEN334 : _GEN332;
wire  _GEN336 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN337 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN338 = io_x[6] ? _GEN337 : _GEN336;
wire  _GEN339 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN340 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN341 = io_x[6] ? _GEN340 : _GEN339;
wire  _GEN342 = io_x[2] ? _GEN341 : _GEN338;
wire  _GEN343 = io_x[14] ? _GEN342 : _GEN335;
wire  _GEN344 = io_x[10] ? _GEN343 : _GEN330;
wire  _GEN345 = io_x[17] ? _GEN344 : _GEN320;
wire  _GEN346 = 1'b1;
wire  _GEN347 = 1'b1;
wire  _GEN348 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN349 = io_x[6] ? _GEN348 : _GEN54;
wire  _GEN350 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN351 = io_x[2] ? _GEN350 : _GEN349;
wire  _GEN352 = io_x[14] ? _GEN351 : _GEN347;
wire  _GEN353 = io_x[10] ? _GEN352 : _GEN346;
wire  _GEN354 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN355 = io_x[6] ? _GEN354 : _GEN54;
wire  _GEN356 = io_x[2] ? _GEN355 : _GEN303;
wire  _GEN357 = io_x[14] ? _GEN356 : _GEN347;
wire  _GEN358 = 1'b0;
wire  _GEN359 = io_x[2] ? _GEN303 : _GEN358;
wire  _GEN360 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN361 = io_x[2] ? _GEN360 : _GEN303;
wire  _GEN362 = io_x[14] ? _GEN361 : _GEN359;
wire  _GEN363 = io_x[10] ? _GEN362 : _GEN357;
wire  _GEN364 = io_x[17] ? _GEN363 : _GEN353;
wire  _GEN365 = io_x[25] ? _GEN364 : _GEN345;
wire  _GEN366 = 1'b0;
wire  _GEN367 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN368 = io_x[6] ? _GEN367 : _GEN54;
wire  _GEN369 = io_x[2] ? _GEN368 : _GEN303;
wire  _GEN370 = io_x[14] ? _GEN369 : _GEN366;
wire  _GEN371 = io_x[2] ? _GEN303 : _GEN358;
wire  _GEN372 = io_x[14] ? _GEN371 : _GEN347;
wire  _GEN373 = io_x[10] ? _GEN372 : _GEN370;
wire  _GEN374 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN375 = io_x[6] ? _GEN374 : _GEN54;
wire  _GEN376 = io_x[2] ? _GEN375 : _GEN303;
wire  _GEN377 = io_x[14] ? _GEN376 : _GEN366;
wire  _GEN378 = io_x[10] ? _GEN377 : _GEN346;
wire  _GEN379 = io_x[17] ? _GEN378 : _GEN373;
wire  _GEN380 = io_x[6] ? _GEN54 : _GEN298;
wire  _GEN381 = io_x[2] ? _GEN380 : _GEN303;
wire  _GEN382 = io_x[14] ? _GEN347 : _GEN381;
wire  _GEN383 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN384 = io_x[6] ? _GEN383 : _GEN54;
wire  _GEN385 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN386 = io_x[6] ? _GEN385 : _GEN54;
wire  _GEN387 = io_x[2] ? _GEN386 : _GEN384;
wire  _GEN388 = io_x[14] ? _GEN387 : _GEN347;
wire  _GEN389 = io_x[10] ? _GEN388 : _GEN382;
wire  _GEN390 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN391 = io_x[6] ? _GEN390 : _GEN54;
wire  _GEN392 = io_x[2] ? _GEN391 : _GEN303;
wire  _GEN393 = io_x[14] ? _GEN392 : _GEN347;
wire  _GEN394 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN395 = io_x[6] ? _GEN394 : _GEN54;
wire  _GEN396 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN397 = io_x[2] ? _GEN396 : _GEN395;
wire  _GEN398 = io_x[14] ? _GEN397 : _GEN347;
wire  _GEN399 = io_x[10] ? _GEN398 : _GEN393;
wire  _GEN400 = io_x[17] ? _GEN399 : _GEN389;
wire  _GEN401 = io_x[25] ? _GEN400 : _GEN379;
wire  _GEN402 = io_x[24] ? _GEN401 : _GEN365;
wire  _GEN403 = io_x[32] ? _GEN402 : _GEN297;
wire  _GEN404 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN405 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN406 = io_x[6] ? _GEN405 : _GEN404;
wire  _GEN407 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN408 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN409 = io_x[6] ? _GEN408 : _GEN407;
wire  _GEN410 = io_x[2] ? _GEN409 : _GEN406;
wire  _GEN411 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN412 = io_x[6] ? _GEN411 : _GEN298;
wire  _GEN413 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN414 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN415 = io_x[6] ? _GEN414 : _GEN413;
wire  _GEN416 = io_x[2] ? _GEN415 : _GEN412;
wire  _GEN417 = io_x[14] ? _GEN416 : _GEN410;
wire  _GEN418 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN419 = io_x[6] ? _GEN418 : _GEN54;
wire  _GEN420 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN421 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN422 = io_x[6] ? _GEN421 : _GEN420;
wire  _GEN423 = io_x[2] ? _GEN422 : _GEN419;
wire  _GEN424 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN425 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN426 = io_x[6] ? _GEN425 : _GEN424;
wire  _GEN427 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN428 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN429 = io_x[6] ? _GEN428 : _GEN427;
wire  _GEN430 = io_x[2] ? _GEN429 : _GEN426;
wire  _GEN431 = io_x[14] ? _GEN430 : _GEN423;
wire  _GEN432 = io_x[10] ? _GEN431 : _GEN417;
wire  _GEN433 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN434 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN435 = io_x[6] ? _GEN434 : _GEN433;
wire  _GEN436 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN437 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN438 = io_x[6] ? _GEN437 : _GEN436;
wire  _GEN439 = io_x[2] ? _GEN438 : _GEN435;
wire  _GEN440 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN441 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN442 = io_x[6] ? _GEN441 : _GEN440;
wire  _GEN443 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN444 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN445 = io_x[6] ? _GEN444 : _GEN443;
wire  _GEN446 = io_x[2] ? _GEN445 : _GEN442;
wire  _GEN447 = io_x[14] ? _GEN446 : _GEN439;
wire  _GEN448 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN449 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN450 = io_x[6] ? _GEN449 : _GEN448;
wire  _GEN451 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN452 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN453 = io_x[6] ? _GEN452 : _GEN451;
wire  _GEN454 = io_x[2] ? _GEN453 : _GEN450;
wire  _GEN455 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN456 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN457 = io_x[6] ? _GEN456 : _GEN455;
wire  _GEN458 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN459 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN460 = io_x[6] ? _GEN459 : _GEN458;
wire  _GEN461 = io_x[2] ? _GEN460 : _GEN457;
wire  _GEN462 = io_x[14] ? _GEN461 : _GEN454;
wire  _GEN463 = io_x[10] ? _GEN462 : _GEN447;
wire  _GEN464 = io_x[17] ? _GEN463 : _GEN432;
wire  _GEN465 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN466 = io_x[6] ? _GEN54 : _GEN465;
wire  _GEN467 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN468 = io_x[6] ? _GEN298 : _GEN467;
wire  _GEN469 = io_x[2] ? _GEN468 : _GEN466;
wire  _GEN470 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN471 = io_x[6] ? _GEN470 : _GEN54;
wire  _GEN472 = io_x[2] ? _GEN358 : _GEN471;
wire  _GEN473 = io_x[14] ? _GEN472 : _GEN469;
wire  _GEN474 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN475 = io_x[6] ? _GEN474 : _GEN298;
wire  _GEN476 = io_x[2] ? _GEN475 : _GEN358;
wire  _GEN477 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN478 = io_x[6] ? _GEN477 : _GEN298;
wire  _GEN479 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN480 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN481 = io_x[6] ? _GEN480 : _GEN479;
wire  _GEN482 = io_x[2] ? _GEN481 : _GEN478;
wire  _GEN483 = io_x[14] ? _GEN482 : _GEN476;
wire  _GEN484 = io_x[10] ? _GEN483 : _GEN473;
wire  _GEN485 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN486 = io_x[6] ? _GEN485 : _GEN298;
wire  _GEN487 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN488 = io_x[2] ? _GEN487 : _GEN486;
wire  _GEN489 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN490 = io_x[6] ? _GEN489 : _GEN298;
wire  _GEN491 = io_x[2] ? _GEN490 : _GEN303;
wire  _GEN492 = io_x[14] ? _GEN491 : _GEN488;
wire  _GEN493 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN494 = io_x[6] ? _GEN493 : _GEN298;
wire  _GEN495 = io_x[2] ? _GEN494 : _GEN358;
wire  _GEN496 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN497 = io_x[6] ? _GEN496 : _GEN54;
wire  _GEN498 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN499 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN500 = io_x[6] ? _GEN499 : _GEN498;
wire  _GEN501 = io_x[2] ? _GEN500 : _GEN497;
wire  _GEN502 = io_x[14] ? _GEN501 : _GEN495;
wire  _GEN503 = io_x[10] ? _GEN502 : _GEN492;
wire  _GEN504 = io_x[17] ? _GEN503 : _GEN484;
wire  _GEN505 = io_x[25] ? _GEN504 : _GEN464;
wire  _GEN506 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN507 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN508 = io_x[6] ? _GEN507 : _GEN506;
wire  _GEN509 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN510 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN511 = io_x[6] ? _GEN510 : _GEN509;
wire  _GEN512 = io_x[2] ? _GEN511 : _GEN508;
wire  _GEN513 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN514 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN515 = io_x[6] ? _GEN514 : _GEN513;
wire  _GEN516 = io_x[2] ? _GEN515 : _GEN303;
wire  _GEN517 = io_x[14] ? _GEN516 : _GEN512;
wire  _GEN518 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN519 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN520 = io_x[6] ? _GEN519 : _GEN518;
wire  _GEN521 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN522 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN523 = io_x[6] ? _GEN522 : _GEN521;
wire  _GEN524 = io_x[2] ? _GEN523 : _GEN520;
wire  _GEN525 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN526 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN527 = io_x[6] ? _GEN526 : _GEN525;
wire  _GEN528 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN529 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN530 = io_x[6] ? _GEN529 : _GEN528;
wire  _GEN531 = io_x[2] ? _GEN530 : _GEN527;
wire  _GEN532 = io_x[14] ? _GEN531 : _GEN524;
wire  _GEN533 = io_x[10] ? _GEN532 : _GEN517;
wire  _GEN534 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN535 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN536 = io_x[6] ? _GEN535 : _GEN534;
wire  _GEN537 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN538 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN539 = io_x[6] ? _GEN538 : _GEN537;
wire  _GEN540 = io_x[2] ? _GEN539 : _GEN536;
wire  _GEN541 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN542 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN543 = io_x[6] ? _GEN542 : _GEN541;
wire  _GEN544 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN545 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN546 = io_x[6] ? _GEN545 : _GEN544;
wire  _GEN547 = io_x[2] ? _GEN546 : _GEN543;
wire  _GEN548 = io_x[14] ? _GEN547 : _GEN540;
wire  _GEN549 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN550 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN551 = io_x[6] ? _GEN550 : _GEN549;
wire  _GEN552 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN553 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN554 = io_x[6] ? _GEN553 : _GEN552;
wire  _GEN555 = io_x[2] ? _GEN554 : _GEN551;
wire  _GEN556 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN557 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN558 = io_x[6] ? _GEN557 : _GEN556;
wire  _GEN559 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN560 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN561 = io_x[6] ? _GEN560 : _GEN559;
wire  _GEN562 = io_x[2] ? _GEN561 : _GEN558;
wire  _GEN563 = io_x[14] ? _GEN562 : _GEN555;
wire  _GEN564 = io_x[10] ? _GEN563 : _GEN548;
wire  _GEN565 = io_x[17] ? _GEN564 : _GEN533;
wire  _GEN566 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN567 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN568 = io_x[6] ? _GEN567 : _GEN566;
wire  _GEN569 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN570 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN571 = io_x[6] ? _GEN570 : _GEN569;
wire  _GEN572 = io_x[2] ? _GEN571 : _GEN568;
wire  _GEN573 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN574 = io_x[6] ? _GEN573 : _GEN54;
wire  _GEN575 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN576 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN577 = io_x[6] ? _GEN576 : _GEN575;
wire  _GEN578 = io_x[2] ? _GEN577 : _GEN574;
wire  _GEN579 = io_x[14] ? _GEN578 : _GEN572;
wire  _GEN580 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN581 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN582 = io_x[6] ? _GEN581 : _GEN580;
wire  _GEN583 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN584 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN585 = io_x[6] ? _GEN584 : _GEN583;
wire  _GEN586 = io_x[2] ? _GEN585 : _GEN582;
wire  _GEN587 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN588 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN589 = io_x[6] ? _GEN588 : _GEN587;
wire  _GEN590 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN591 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN592 = io_x[6] ? _GEN591 : _GEN590;
wire  _GEN593 = io_x[2] ? _GEN592 : _GEN589;
wire  _GEN594 = io_x[14] ? _GEN593 : _GEN586;
wire  _GEN595 = io_x[10] ? _GEN594 : _GEN579;
wire  _GEN596 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN597 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN598 = io_x[6] ? _GEN597 : _GEN596;
wire  _GEN599 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN600 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN601 = io_x[6] ? _GEN600 : _GEN599;
wire  _GEN602 = io_x[2] ? _GEN601 : _GEN598;
wire  _GEN603 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN604 = io_x[6] ? _GEN603 : _GEN54;
wire  _GEN605 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN606 = io_x[6] ? _GEN605 : _GEN298;
wire  _GEN607 = io_x[2] ? _GEN606 : _GEN604;
wire  _GEN608 = io_x[14] ? _GEN607 : _GEN602;
wire  _GEN609 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN610 = io_x[6] ? _GEN609 : _GEN54;
wire  _GEN611 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN612 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN613 = io_x[6] ? _GEN612 : _GEN611;
wire  _GEN614 = io_x[2] ? _GEN613 : _GEN610;
wire  _GEN615 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN616 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN617 = io_x[6] ? _GEN616 : _GEN615;
wire  _GEN618 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN619 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN620 = io_x[6] ? _GEN619 : _GEN618;
wire  _GEN621 = io_x[2] ? _GEN620 : _GEN617;
wire  _GEN622 = io_x[14] ? _GEN621 : _GEN614;
wire  _GEN623 = io_x[10] ? _GEN622 : _GEN608;
wire  _GEN624 = io_x[17] ? _GEN623 : _GEN595;
wire  _GEN625 = io_x[25] ? _GEN624 : _GEN565;
wire  _GEN626 = io_x[24] ? _GEN625 : _GEN505;
wire  _GEN627 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN628 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN629 = io_x[6] ? _GEN628 : _GEN627;
wire  _GEN630 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN631 = io_x[6] ? _GEN54 : _GEN630;
wire  _GEN632 = io_x[2] ? _GEN631 : _GEN629;
wire  _GEN633 = io_x[14] ? _GEN366 : _GEN632;
wire  _GEN634 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN635 = io_x[6] ? _GEN634 : _GEN298;
wire  _GEN636 = io_x[2] ? _GEN635 : _GEN358;
wire  _GEN637 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN638 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN639 = io_x[6] ? _GEN638 : _GEN637;
wire  _GEN640 = io_x[2] ? _GEN639 : _GEN303;
wire  _GEN641 = io_x[14] ? _GEN640 : _GEN636;
wire  _GEN642 = io_x[10] ? _GEN641 : _GEN633;
wire  _GEN643 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN644 = io_x[6] ? _GEN54 : _GEN643;
wire  _GEN645 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN646 = io_x[6] ? _GEN54 : _GEN645;
wire  _GEN647 = io_x[2] ? _GEN646 : _GEN644;
wire  _GEN648 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN649 = io_x[6] ? _GEN648 : _GEN54;
wire  _GEN650 = io_x[2] ? _GEN649 : _GEN358;
wire  _GEN651 = io_x[14] ? _GEN650 : _GEN647;
wire  _GEN652 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN653 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN654 = io_x[6] ? _GEN653 : _GEN298;
wire  _GEN655 = io_x[2] ? _GEN654 : _GEN652;
wire  _GEN656 = io_x[6] ? _GEN54 : _GEN298;
wire  _GEN657 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN658 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN659 = io_x[6] ? _GEN658 : _GEN657;
wire  _GEN660 = io_x[2] ? _GEN659 : _GEN656;
wire  _GEN661 = io_x[14] ? _GEN660 : _GEN655;
wire  _GEN662 = io_x[10] ? _GEN661 : _GEN651;
wire  _GEN663 = io_x[17] ? _GEN662 : _GEN642;
wire  _GEN664 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN665 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN666 = io_x[6] ? _GEN665 : _GEN664;
wire  _GEN667 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN668 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN669 = io_x[6] ? _GEN668 : _GEN667;
wire  _GEN670 = io_x[2] ? _GEN669 : _GEN666;
wire  _GEN671 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN672 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN673 = io_x[6] ? _GEN672 : _GEN671;
wire  _GEN674 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN675 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN676 = io_x[6] ? _GEN675 : _GEN674;
wire  _GEN677 = io_x[2] ? _GEN676 : _GEN673;
wire  _GEN678 = io_x[14] ? _GEN677 : _GEN670;
wire  _GEN679 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN680 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN681 = io_x[6] ? _GEN680 : _GEN679;
wire  _GEN682 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN683 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN684 = io_x[6] ? _GEN683 : _GEN682;
wire  _GEN685 = io_x[2] ? _GEN684 : _GEN681;
wire  _GEN686 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN687 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN688 = io_x[6] ? _GEN687 : _GEN686;
wire  _GEN689 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN690 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN691 = io_x[6] ? _GEN690 : _GEN689;
wire  _GEN692 = io_x[2] ? _GEN691 : _GEN688;
wire  _GEN693 = io_x[14] ? _GEN692 : _GEN685;
wire  _GEN694 = io_x[10] ? _GEN693 : _GEN678;
wire  _GEN695 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN696 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN697 = io_x[6] ? _GEN696 : _GEN695;
wire  _GEN698 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN699 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN700 = io_x[6] ? _GEN699 : _GEN698;
wire  _GEN701 = io_x[2] ? _GEN700 : _GEN697;
wire  _GEN702 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN703 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN704 = io_x[6] ? _GEN703 : _GEN702;
wire  _GEN705 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN706 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN707 = io_x[6] ? _GEN706 : _GEN705;
wire  _GEN708 = io_x[2] ? _GEN707 : _GEN704;
wire  _GEN709 = io_x[14] ? _GEN708 : _GEN701;
wire  _GEN710 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN711 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN712 = io_x[6] ? _GEN711 : _GEN710;
wire  _GEN713 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN714 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN715 = io_x[6] ? _GEN714 : _GEN713;
wire  _GEN716 = io_x[2] ? _GEN715 : _GEN712;
wire  _GEN717 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN718 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN719 = io_x[6] ? _GEN718 : _GEN717;
wire  _GEN720 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN721 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN722 = io_x[6] ? _GEN721 : _GEN720;
wire  _GEN723 = io_x[2] ? _GEN722 : _GEN719;
wire  _GEN724 = io_x[14] ? _GEN723 : _GEN716;
wire  _GEN725 = io_x[10] ? _GEN724 : _GEN709;
wire  _GEN726 = io_x[17] ? _GEN725 : _GEN694;
wire  _GEN727 = io_x[25] ? _GEN726 : _GEN663;
wire  _GEN728 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN729 = io_x[6] ? _GEN54 : _GEN728;
wire  _GEN730 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN731 = io_x[6] ? _GEN298 : _GEN730;
wire  _GEN732 = io_x[2] ? _GEN731 : _GEN729;
wire  _GEN733 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN734 = io_x[6] ? _GEN298 : _GEN733;
wire  _GEN735 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN736 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN737 = io_x[6] ? _GEN736 : _GEN735;
wire  _GEN738 = io_x[2] ? _GEN737 : _GEN734;
wire  _GEN739 = io_x[14] ? _GEN738 : _GEN732;
wire  _GEN740 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN741 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN742 = io_x[6] ? _GEN54 : _GEN741;
wire  _GEN743 = io_x[2] ? _GEN742 : _GEN740;
wire  _GEN744 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN745 = io_x[6] ? _GEN54 : _GEN744;
wire  _GEN746 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN747 = io_x[6] ? _GEN298 : _GEN746;
wire  _GEN748 = io_x[2] ? _GEN747 : _GEN745;
wire  _GEN749 = io_x[14] ? _GEN748 : _GEN743;
wire  _GEN750 = io_x[10] ? _GEN749 : _GEN739;
wire  _GEN751 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN752 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN753 = io_x[6] ? _GEN752 : _GEN751;
wire  _GEN754 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN755 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN756 = io_x[6] ? _GEN755 : _GEN754;
wire  _GEN757 = io_x[2] ? _GEN756 : _GEN753;
wire  _GEN758 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN759 = io_x[6] ? _GEN298 : _GEN758;
wire  _GEN760 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN761 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN762 = io_x[6] ? _GEN761 : _GEN760;
wire  _GEN763 = io_x[2] ? _GEN762 : _GEN759;
wire  _GEN764 = io_x[14] ? _GEN763 : _GEN757;
wire  _GEN765 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN766 = io_x[6] ? _GEN298 : _GEN765;
wire  _GEN767 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN768 = io_x[6] ? _GEN54 : _GEN767;
wire  _GEN769 = io_x[2] ? _GEN768 : _GEN766;
wire  _GEN770 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN771 = io_x[6] ? _GEN54 : _GEN770;
wire  _GEN772 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN773 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN774 = io_x[6] ? _GEN773 : _GEN772;
wire  _GEN775 = io_x[2] ? _GEN774 : _GEN771;
wire  _GEN776 = io_x[14] ? _GEN775 : _GEN769;
wire  _GEN777 = io_x[10] ? _GEN776 : _GEN764;
wire  _GEN778 = io_x[17] ? _GEN777 : _GEN750;
wire  _GEN779 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN780 = io_x[6] ? _GEN298 : _GEN779;
wire  _GEN781 = io_x[2] ? _GEN303 : _GEN780;
wire  _GEN782 = io_x[14] ? _GEN347 : _GEN781;
wire  _GEN783 = io_x[10] ? _GEN346 : _GEN782;
wire  _GEN784 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN785 = io_x[2] ? _GEN303 : _GEN784;
wire  _GEN786 = io_x[14] ? _GEN347 : _GEN785;
wire  _GEN787 = io_x[10] ? _GEN346 : _GEN786;
wire  _GEN788 = io_x[17] ? _GEN787 : _GEN783;
wire  _GEN789 = io_x[25] ? _GEN788 : _GEN778;
wire  _GEN790 = io_x[24] ? _GEN789 : _GEN727;
wire  _GEN791 = io_x[32] ? _GEN790 : _GEN626;
wire  _GEN792 = io_x[28] ? _GEN791 : _GEN403;
wire  _GEN793 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN794 = io_x[6] ? _GEN298 : _GEN793;
wire  _GEN795 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN796 = io_x[6] ? _GEN795 : _GEN298;
wire  _GEN797 = io_x[2] ? _GEN796 : _GEN794;
wire  _GEN798 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN799 = io_x[6] ? _GEN798 : _GEN298;
wire  _GEN800 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN801 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN802 = io_x[6] ? _GEN801 : _GEN800;
wire  _GEN803 = io_x[2] ? _GEN802 : _GEN799;
wire  _GEN804 = io_x[14] ? _GEN803 : _GEN797;
wire  _GEN805 = io_x[6] ? _GEN54 : _GEN298;
wire  _GEN806 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN807 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN808 = io_x[6] ? _GEN807 : _GEN806;
wire  _GEN809 = io_x[2] ? _GEN808 : _GEN805;
wire  _GEN810 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN811 = io_x[6] ? _GEN810 : _GEN54;
wire  _GEN812 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN813 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN814 = io_x[6] ? _GEN813 : _GEN812;
wire  _GEN815 = io_x[2] ? _GEN814 : _GEN811;
wire  _GEN816 = io_x[14] ? _GEN815 : _GEN809;
wire  _GEN817 = io_x[10] ? _GEN816 : _GEN804;
wire  _GEN818 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN819 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN820 = io_x[6] ? _GEN819 : _GEN818;
wire  _GEN821 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN822 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN823 = io_x[6] ? _GEN822 : _GEN821;
wire  _GEN824 = io_x[2] ? _GEN823 : _GEN820;
wire  _GEN825 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN826 = io_x[6] ? _GEN825 : _GEN298;
wire  _GEN827 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN828 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN829 = io_x[6] ? _GEN828 : _GEN827;
wire  _GEN830 = io_x[2] ? _GEN829 : _GEN826;
wire  _GEN831 = io_x[14] ? _GEN830 : _GEN824;
wire  _GEN832 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN833 = io_x[6] ? _GEN832 : _GEN298;
wire  _GEN834 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN835 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN836 = io_x[6] ? _GEN835 : _GEN834;
wire  _GEN837 = io_x[2] ? _GEN836 : _GEN833;
wire  _GEN838 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN839 = io_x[6] ? _GEN838 : _GEN54;
wire  _GEN840 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN841 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN842 = io_x[6] ? _GEN841 : _GEN840;
wire  _GEN843 = io_x[2] ? _GEN842 : _GEN839;
wire  _GEN844 = io_x[14] ? _GEN843 : _GEN837;
wire  _GEN845 = io_x[10] ? _GEN844 : _GEN831;
wire  _GEN846 = io_x[17] ? _GEN845 : _GEN817;
wire  _GEN847 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN848 = io_x[6] ? _GEN54 : _GEN847;
wire  _GEN849 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN850 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN851 = io_x[6] ? _GEN850 : _GEN849;
wire  _GEN852 = io_x[2] ? _GEN851 : _GEN848;
wire  _GEN853 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN854 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN855 = io_x[6] ? _GEN854 : _GEN298;
wire  _GEN856 = io_x[2] ? _GEN855 : _GEN853;
wire  _GEN857 = io_x[14] ? _GEN856 : _GEN852;
wire  _GEN858 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN859 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN860 = io_x[6] ? _GEN859 : _GEN858;
wire  _GEN861 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN862 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN863 = io_x[6] ? _GEN862 : _GEN861;
wire  _GEN864 = io_x[2] ? _GEN863 : _GEN860;
wire  _GEN865 = io_x[6] ? _GEN54 : _GEN298;
wire  _GEN866 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN867 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN868 = io_x[6] ? _GEN867 : _GEN866;
wire  _GEN869 = io_x[2] ? _GEN868 : _GEN865;
wire  _GEN870 = io_x[14] ? _GEN869 : _GEN864;
wire  _GEN871 = io_x[10] ? _GEN870 : _GEN857;
wire  _GEN872 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN873 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN874 = io_x[6] ? _GEN873 : _GEN872;
wire  _GEN875 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN876 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN877 = io_x[6] ? _GEN876 : _GEN875;
wire  _GEN878 = io_x[2] ? _GEN877 : _GEN874;
wire  _GEN879 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN880 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN881 = io_x[6] ? _GEN880 : _GEN879;
wire  _GEN882 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN883 = io_x[6] ? _GEN882 : _GEN298;
wire  _GEN884 = io_x[2] ? _GEN883 : _GEN881;
wire  _GEN885 = io_x[14] ? _GEN884 : _GEN878;
wire  _GEN886 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN887 = io_x[6] ? _GEN886 : _GEN54;
wire  _GEN888 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN889 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN890 = io_x[6] ? _GEN889 : _GEN888;
wire  _GEN891 = io_x[2] ? _GEN890 : _GEN887;
wire  _GEN892 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN893 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN894 = io_x[6] ? _GEN893 : _GEN892;
wire  _GEN895 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN896 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN897 = io_x[6] ? _GEN896 : _GEN895;
wire  _GEN898 = io_x[2] ? _GEN897 : _GEN894;
wire  _GEN899 = io_x[14] ? _GEN898 : _GEN891;
wire  _GEN900 = io_x[10] ? _GEN899 : _GEN885;
wire  _GEN901 = io_x[17] ? _GEN900 : _GEN871;
wire  _GEN902 = io_x[25] ? _GEN901 : _GEN846;
wire  _GEN903 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN904 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN905 = io_x[6] ? _GEN904 : _GEN903;
wire  _GEN906 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN907 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN908 = io_x[6] ? _GEN907 : _GEN906;
wire  _GEN909 = io_x[2] ? _GEN908 : _GEN905;
wire  _GEN910 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN911 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN912 = io_x[6] ? _GEN911 : _GEN910;
wire  _GEN913 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN914 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN915 = io_x[6] ? _GEN914 : _GEN913;
wire  _GEN916 = io_x[2] ? _GEN915 : _GEN912;
wire  _GEN917 = io_x[14] ? _GEN916 : _GEN909;
wire  _GEN918 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN919 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN920 = io_x[6] ? _GEN919 : _GEN918;
wire  _GEN921 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN922 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN923 = io_x[6] ? _GEN922 : _GEN921;
wire  _GEN924 = io_x[2] ? _GEN923 : _GEN920;
wire  _GEN925 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN926 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN927 = io_x[6] ? _GEN926 : _GEN925;
wire  _GEN928 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN929 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN930 = io_x[6] ? _GEN929 : _GEN928;
wire  _GEN931 = io_x[2] ? _GEN930 : _GEN927;
wire  _GEN932 = io_x[14] ? _GEN931 : _GEN924;
wire  _GEN933 = io_x[10] ? _GEN932 : _GEN917;
wire  _GEN934 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN935 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN936 = io_x[6] ? _GEN935 : _GEN934;
wire  _GEN937 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN938 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN939 = io_x[6] ? _GEN938 : _GEN937;
wire  _GEN940 = io_x[2] ? _GEN939 : _GEN936;
wire  _GEN941 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN942 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN943 = io_x[6] ? _GEN942 : _GEN941;
wire  _GEN944 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN945 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN946 = io_x[6] ? _GEN945 : _GEN944;
wire  _GEN947 = io_x[2] ? _GEN946 : _GEN943;
wire  _GEN948 = io_x[14] ? _GEN947 : _GEN940;
wire  _GEN949 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN950 = io_x[6] ? _GEN949 : _GEN298;
wire  _GEN951 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN952 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN953 = io_x[6] ? _GEN952 : _GEN951;
wire  _GEN954 = io_x[2] ? _GEN953 : _GEN950;
wire  _GEN955 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN956 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN957 = io_x[6] ? _GEN956 : _GEN955;
wire  _GEN958 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN959 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN960 = io_x[6] ? _GEN959 : _GEN958;
wire  _GEN961 = io_x[2] ? _GEN960 : _GEN957;
wire  _GEN962 = io_x[14] ? _GEN961 : _GEN954;
wire  _GEN963 = io_x[10] ? _GEN962 : _GEN948;
wire  _GEN964 = io_x[17] ? _GEN963 : _GEN933;
wire  _GEN965 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN966 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN967 = io_x[6] ? _GEN966 : _GEN965;
wire  _GEN968 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN969 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN970 = io_x[6] ? _GEN969 : _GEN968;
wire  _GEN971 = io_x[2] ? _GEN970 : _GEN967;
wire  _GEN972 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN973 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN974 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN975 = io_x[6] ? _GEN974 : _GEN973;
wire  _GEN976 = io_x[2] ? _GEN975 : _GEN972;
wire  _GEN977 = io_x[14] ? _GEN976 : _GEN971;
wire  _GEN978 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN979 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN980 = io_x[6] ? _GEN979 : _GEN298;
wire  _GEN981 = io_x[2] ? _GEN980 : _GEN978;
wire  _GEN982 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN983 = io_x[6] ? _GEN982 : _GEN298;
wire  _GEN984 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN985 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN986 = io_x[6] ? _GEN985 : _GEN984;
wire  _GEN987 = io_x[2] ? _GEN986 : _GEN983;
wire  _GEN988 = io_x[14] ? _GEN987 : _GEN981;
wire  _GEN989 = io_x[10] ? _GEN988 : _GEN977;
wire  _GEN990 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN991 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN992 = io_x[6] ? _GEN991 : _GEN990;
wire  _GEN993 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN994 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN995 = io_x[6] ? _GEN994 : _GEN993;
wire  _GEN996 = io_x[2] ? _GEN995 : _GEN992;
wire  _GEN997 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN998 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN999 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1000 = io_x[6] ? _GEN999 : _GEN998;
wire  _GEN1001 = io_x[2] ? _GEN1000 : _GEN997;
wire  _GEN1002 = io_x[14] ? _GEN1001 : _GEN996;
wire  _GEN1003 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN1004 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1005 = io_x[6] ? _GEN1004 : _GEN298;
wire  _GEN1006 = io_x[2] ? _GEN1005 : _GEN1003;
wire  _GEN1007 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1008 = io_x[6] ? _GEN1007 : _GEN298;
wire  _GEN1009 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1010 = io_x[6] ? _GEN1009 : _GEN54;
wire  _GEN1011 = io_x[2] ? _GEN1010 : _GEN1008;
wire  _GEN1012 = io_x[14] ? _GEN1011 : _GEN1006;
wire  _GEN1013 = io_x[10] ? _GEN1012 : _GEN1002;
wire  _GEN1014 = io_x[17] ? _GEN1013 : _GEN989;
wire  _GEN1015 = io_x[25] ? _GEN1014 : _GEN964;
wire  _GEN1016 = io_x[24] ? _GEN1015 : _GEN902;
wire  _GEN1017 = io_x[2] ? _GEN303 : _GEN358;
wire  _GEN1018 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1019 = io_x[6] ? _GEN1018 : _GEN54;
wire  _GEN1020 = io_x[2] ? _GEN1019 : _GEN303;
wire  _GEN1021 = io_x[14] ? _GEN1020 : _GEN1017;
wire  _GEN1022 = io_x[6] ? _GEN54 : _GEN298;
wire  _GEN1023 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1024 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1025 = io_x[6] ? _GEN1024 : _GEN1023;
wire  _GEN1026 = io_x[2] ? _GEN1025 : _GEN1022;
wire  _GEN1027 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1028 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1029 = io_x[6] ? _GEN1028 : _GEN1027;
wire  _GEN1030 = io_x[2] ? _GEN1029 : _GEN358;
wire  _GEN1031 = io_x[14] ? _GEN1030 : _GEN1026;
wire  _GEN1032 = io_x[10] ? _GEN1031 : _GEN1021;
wire  _GEN1033 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1034 = io_x[6] ? _GEN298 : _GEN1033;
wire  _GEN1035 = io_x[2] ? _GEN303 : _GEN1034;
wire  _GEN1036 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1037 = io_x[6] ? _GEN1036 : _GEN54;
wire  _GEN1038 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1039 = io_x[6] ? _GEN1038 : _GEN54;
wire  _GEN1040 = io_x[2] ? _GEN1039 : _GEN1037;
wire  _GEN1041 = io_x[14] ? _GEN1040 : _GEN1035;
wire  _GEN1042 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1043 = io_x[6] ? _GEN1042 : _GEN54;
wire  _GEN1044 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1045 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1046 = io_x[6] ? _GEN1045 : _GEN1044;
wire  _GEN1047 = io_x[2] ? _GEN1046 : _GEN1043;
wire  _GEN1048 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1049 = io_x[6] ? _GEN1048 : _GEN54;
wire  _GEN1050 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1051 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1052 = io_x[6] ? _GEN1051 : _GEN1050;
wire  _GEN1053 = io_x[2] ? _GEN1052 : _GEN1049;
wire  _GEN1054 = io_x[14] ? _GEN1053 : _GEN1047;
wire  _GEN1055 = io_x[10] ? _GEN1054 : _GEN1041;
wire  _GEN1056 = io_x[17] ? _GEN1055 : _GEN1032;
wire  _GEN1057 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1058 = io_x[6] ? _GEN298 : _GEN1057;
wire  _GEN1059 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1060 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1061 = io_x[6] ? _GEN1060 : _GEN1059;
wire  _GEN1062 = io_x[2] ? _GEN1061 : _GEN1058;
wire  _GEN1063 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1064 = io_x[6] ? _GEN298 : _GEN1063;
wire  _GEN1065 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN1066 = io_x[2] ? _GEN1065 : _GEN1064;
wire  _GEN1067 = io_x[14] ? _GEN1066 : _GEN1062;
wire  _GEN1068 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1069 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1070 = io_x[6] ? _GEN1069 : _GEN1068;
wire  _GEN1071 = io_x[2] ? _GEN1070 : _GEN358;
wire  _GEN1072 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1073 = io_x[6] ? _GEN54 : _GEN1072;
wire  _GEN1074 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1075 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1076 = io_x[6] ? _GEN1075 : _GEN1074;
wire  _GEN1077 = io_x[2] ? _GEN1076 : _GEN1073;
wire  _GEN1078 = io_x[14] ? _GEN1077 : _GEN1071;
wire  _GEN1079 = io_x[10] ? _GEN1078 : _GEN1067;
wire  _GEN1080 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1081 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1082 = io_x[6] ? _GEN1081 : _GEN1080;
wire  _GEN1083 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1084 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1085 = io_x[6] ? _GEN1084 : _GEN1083;
wire  _GEN1086 = io_x[2] ? _GEN1085 : _GEN1082;
wire  _GEN1087 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1088 = io_x[6] ? _GEN54 : _GEN1087;
wire  _GEN1089 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1090 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1091 = io_x[6] ? _GEN1090 : _GEN1089;
wire  _GEN1092 = io_x[2] ? _GEN1091 : _GEN1088;
wire  _GEN1093 = io_x[14] ? _GEN1092 : _GEN1086;
wire  _GEN1094 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1095 = io_x[6] ? _GEN1094 : _GEN298;
wire  _GEN1096 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1097 = io_x[6] ? _GEN1096 : _GEN54;
wire  _GEN1098 = io_x[2] ? _GEN1097 : _GEN1095;
wire  _GEN1099 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1100 = io_x[6] ? _GEN54 : _GEN1099;
wire  _GEN1101 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1102 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1103 = io_x[6] ? _GEN1102 : _GEN1101;
wire  _GEN1104 = io_x[2] ? _GEN1103 : _GEN1100;
wire  _GEN1105 = io_x[14] ? _GEN1104 : _GEN1098;
wire  _GEN1106 = io_x[10] ? _GEN1105 : _GEN1093;
wire  _GEN1107 = io_x[17] ? _GEN1106 : _GEN1079;
wire  _GEN1108 = io_x[25] ? _GEN1107 : _GEN1056;
wire  _GEN1109 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1110 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1111 = io_x[6] ? _GEN1110 : _GEN1109;
wire  _GEN1112 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1113 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1114 = io_x[6] ? _GEN1113 : _GEN1112;
wire  _GEN1115 = io_x[2] ? _GEN1114 : _GEN1111;
wire  _GEN1116 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1117 = io_x[6] ? _GEN1116 : _GEN298;
wire  _GEN1118 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1119 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1120 = io_x[6] ? _GEN1119 : _GEN1118;
wire  _GEN1121 = io_x[2] ? _GEN1120 : _GEN1117;
wire  _GEN1122 = io_x[14] ? _GEN1121 : _GEN1115;
wire  _GEN1123 = io_x[6] ? _GEN54 : _GEN298;
wire  _GEN1124 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1125 = io_x[6] ? _GEN1124 : _GEN54;
wire  _GEN1126 = io_x[2] ? _GEN1125 : _GEN1123;
wire  _GEN1127 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1128 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1129 = io_x[6] ? _GEN1128 : _GEN1127;
wire  _GEN1130 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1131 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1132 = io_x[6] ? _GEN1131 : _GEN1130;
wire  _GEN1133 = io_x[2] ? _GEN1132 : _GEN1129;
wire  _GEN1134 = io_x[14] ? _GEN1133 : _GEN1126;
wire  _GEN1135 = io_x[10] ? _GEN1134 : _GEN1122;
wire  _GEN1136 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1137 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1138 = io_x[6] ? _GEN1137 : _GEN1136;
wire  _GEN1139 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1140 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1141 = io_x[6] ? _GEN1140 : _GEN1139;
wire  _GEN1142 = io_x[2] ? _GEN1141 : _GEN1138;
wire  _GEN1143 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1144 = io_x[6] ? _GEN1143 : _GEN298;
wire  _GEN1145 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1146 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1147 = io_x[6] ? _GEN1146 : _GEN1145;
wire  _GEN1148 = io_x[2] ? _GEN1147 : _GEN1144;
wire  _GEN1149 = io_x[14] ? _GEN1148 : _GEN1142;
wire  _GEN1150 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1151 = io_x[6] ? _GEN1150 : _GEN298;
wire  _GEN1152 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1153 = io_x[6] ? _GEN1152 : _GEN54;
wire  _GEN1154 = io_x[2] ? _GEN1153 : _GEN1151;
wire  _GEN1155 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1156 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1157 = io_x[6] ? _GEN1156 : _GEN1155;
wire  _GEN1158 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1159 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1160 = io_x[6] ? _GEN1159 : _GEN1158;
wire  _GEN1161 = io_x[2] ? _GEN1160 : _GEN1157;
wire  _GEN1162 = io_x[14] ? _GEN1161 : _GEN1154;
wire  _GEN1163 = io_x[10] ? _GEN1162 : _GEN1149;
wire  _GEN1164 = io_x[17] ? _GEN1163 : _GEN1135;
wire  _GEN1165 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1166 = io_x[6] ? _GEN298 : _GEN1165;
wire  _GEN1167 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1168 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1169 = io_x[6] ? _GEN1168 : _GEN1167;
wire  _GEN1170 = io_x[2] ? _GEN1169 : _GEN1166;
wire  _GEN1171 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1172 = io_x[6] ? _GEN54 : _GEN1171;
wire  _GEN1173 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1174 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1175 = io_x[6] ? _GEN1174 : _GEN1173;
wire  _GEN1176 = io_x[2] ? _GEN1175 : _GEN1172;
wire  _GEN1177 = io_x[14] ? _GEN1176 : _GEN1170;
wire  _GEN1178 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1179 = io_x[6] ? _GEN1178 : _GEN298;
wire  _GEN1180 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1181 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1182 = io_x[6] ? _GEN1181 : _GEN1180;
wire  _GEN1183 = io_x[2] ? _GEN1182 : _GEN1179;
wire  _GEN1184 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1185 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1186 = io_x[6] ? _GEN1185 : _GEN1184;
wire  _GEN1187 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1188 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1189 = io_x[6] ? _GEN1188 : _GEN1187;
wire  _GEN1190 = io_x[2] ? _GEN1189 : _GEN1186;
wire  _GEN1191 = io_x[14] ? _GEN1190 : _GEN1183;
wire  _GEN1192 = io_x[10] ? _GEN1191 : _GEN1177;
wire  _GEN1193 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN1194 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1195 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1196 = io_x[6] ? _GEN1195 : _GEN1194;
wire  _GEN1197 = io_x[2] ? _GEN1196 : _GEN1193;
wire  _GEN1198 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1199 = io_x[6] ? _GEN1198 : _GEN298;
wire  _GEN1200 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1201 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1202 = io_x[6] ? _GEN1201 : _GEN1200;
wire  _GEN1203 = io_x[2] ? _GEN1202 : _GEN1199;
wire  _GEN1204 = io_x[14] ? _GEN1203 : _GEN1197;
wire  _GEN1205 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1206 = io_x[6] ? _GEN1205 : _GEN298;
wire  _GEN1207 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1208 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1209 = io_x[6] ? _GEN1208 : _GEN1207;
wire  _GEN1210 = io_x[2] ? _GEN1209 : _GEN1206;
wire  _GEN1211 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1212 = io_x[6] ? _GEN1211 : _GEN54;
wire  _GEN1213 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1214 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1215 = io_x[6] ? _GEN1214 : _GEN1213;
wire  _GEN1216 = io_x[2] ? _GEN1215 : _GEN1212;
wire  _GEN1217 = io_x[14] ? _GEN1216 : _GEN1210;
wire  _GEN1218 = io_x[10] ? _GEN1217 : _GEN1204;
wire  _GEN1219 = io_x[17] ? _GEN1218 : _GEN1192;
wire  _GEN1220 = io_x[25] ? _GEN1219 : _GEN1164;
wire  _GEN1221 = io_x[24] ? _GEN1220 : _GEN1108;
wire  _GEN1222 = io_x[32] ? _GEN1221 : _GEN1016;
wire  _GEN1223 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1224 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1225 = io_x[6] ? _GEN1224 : _GEN1223;
wire  _GEN1226 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1227 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1228 = io_x[6] ? _GEN1227 : _GEN1226;
wire  _GEN1229 = io_x[2] ? _GEN1228 : _GEN1225;
wire  _GEN1230 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1231 = io_x[6] ? _GEN1230 : _GEN54;
wire  _GEN1232 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1233 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1234 = io_x[6] ? _GEN1233 : _GEN1232;
wire  _GEN1235 = io_x[2] ? _GEN1234 : _GEN1231;
wire  _GEN1236 = io_x[14] ? _GEN1235 : _GEN1229;
wire  _GEN1237 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1238 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1239 = io_x[6] ? _GEN1238 : _GEN1237;
wire  _GEN1240 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1241 = io_x[6] ? _GEN1240 : _GEN298;
wire  _GEN1242 = io_x[2] ? _GEN1241 : _GEN1239;
wire  _GEN1243 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1244 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1245 = io_x[6] ? _GEN1244 : _GEN1243;
wire  _GEN1246 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1247 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1248 = io_x[6] ? _GEN1247 : _GEN1246;
wire  _GEN1249 = io_x[2] ? _GEN1248 : _GEN1245;
wire  _GEN1250 = io_x[14] ? _GEN1249 : _GEN1242;
wire  _GEN1251 = io_x[10] ? _GEN1250 : _GEN1236;
wire  _GEN1252 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1253 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1254 = io_x[6] ? _GEN1253 : _GEN1252;
wire  _GEN1255 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1256 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1257 = io_x[6] ? _GEN1256 : _GEN1255;
wire  _GEN1258 = io_x[2] ? _GEN1257 : _GEN1254;
wire  _GEN1259 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1260 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1261 = io_x[6] ? _GEN1260 : _GEN1259;
wire  _GEN1262 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1263 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1264 = io_x[6] ? _GEN1263 : _GEN1262;
wire  _GEN1265 = io_x[2] ? _GEN1264 : _GEN1261;
wire  _GEN1266 = io_x[14] ? _GEN1265 : _GEN1258;
wire  _GEN1267 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1268 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1269 = io_x[6] ? _GEN1268 : _GEN1267;
wire  _GEN1270 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1271 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1272 = io_x[6] ? _GEN1271 : _GEN1270;
wire  _GEN1273 = io_x[2] ? _GEN1272 : _GEN1269;
wire  _GEN1274 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1275 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1276 = io_x[6] ? _GEN1275 : _GEN1274;
wire  _GEN1277 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1278 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1279 = io_x[6] ? _GEN1278 : _GEN1277;
wire  _GEN1280 = io_x[2] ? _GEN1279 : _GEN1276;
wire  _GEN1281 = io_x[14] ? _GEN1280 : _GEN1273;
wire  _GEN1282 = io_x[10] ? _GEN1281 : _GEN1266;
wire  _GEN1283 = io_x[17] ? _GEN1282 : _GEN1251;
wire  _GEN1284 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1285 = io_x[6] ? _GEN1284 : _GEN298;
wire  _GEN1286 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1287 = io_x[6] ? _GEN1286 : _GEN54;
wire  _GEN1288 = io_x[2] ? _GEN1287 : _GEN1285;
wire  _GEN1289 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1290 = io_x[6] ? _GEN1289 : _GEN54;
wire  _GEN1291 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1292 = io_x[6] ? _GEN1291 : _GEN298;
wire  _GEN1293 = io_x[2] ? _GEN1292 : _GEN1290;
wire  _GEN1294 = io_x[14] ? _GEN1293 : _GEN1288;
wire  _GEN1295 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1296 = io_x[6] ? _GEN1295 : _GEN54;
wire  _GEN1297 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1298 = io_x[6] ? _GEN1297 : _GEN298;
wire  _GEN1299 = io_x[2] ? _GEN1298 : _GEN1296;
wire  _GEN1300 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1301 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1302 = io_x[6] ? _GEN1301 : _GEN1300;
wire  _GEN1303 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1304 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1305 = io_x[6] ? _GEN1304 : _GEN1303;
wire  _GEN1306 = io_x[2] ? _GEN1305 : _GEN1302;
wire  _GEN1307 = io_x[14] ? _GEN1306 : _GEN1299;
wire  _GEN1308 = io_x[10] ? _GEN1307 : _GEN1294;
wire  _GEN1309 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1310 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1311 = io_x[6] ? _GEN1310 : _GEN1309;
wire  _GEN1312 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1313 = io_x[6] ? _GEN1312 : _GEN54;
wire  _GEN1314 = io_x[2] ? _GEN1313 : _GEN1311;
wire  _GEN1315 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN1316 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1317 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1318 = io_x[6] ? _GEN1317 : _GEN1316;
wire  _GEN1319 = io_x[2] ? _GEN1318 : _GEN1315;
wire  _GEN1320 = io_x[14] ? _GEN1319 : _GEN1314;
wire  _GEN1321 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1322 = io_x[6] ? _GEN1321 : _GEN54;
wire  _GEN1323 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1324 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1325 = io_x[6] ? _GEN1324 : _GEN1323;
wire  _GEN1326 = io_x[2] ? _GEN1325 : _GEN1322;
wire  _GEN1327 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1328 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1329 = io_x[6] ? _GEN1328 : _GEN1327;
wire  _GEN1330 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1331 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1332 = io_x[6] ? _GEN1331 : _GEN1330;
wire  _GEN1333 = io_x[2] ? _GEN1332 : _GEN1329;
wire  _GEN1334 = io_x[14] ? _GEN1333 : _GEN1326;
wire  _GEN1335 = io_x[10] ? _GEN1334 : _GEN1320;
wire  _GEN1336 = io_x[17] ? _GEN1335 : _GEN1308;
wire  _GEN1337 = io_x[25] ? _GEN1336 : _GEN1283;
wire  _GEN1338 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1339 = io_x[6] ? _GEN54 : _GEN1338;
wire  _GEN1340 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1341 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1342 = io_x[6] ? _GEN1341 : _GEN1340;
wire  _GEN1343 = io_x[2] ? _GEN1342 : _GEN1339;
wire  _GEN1344 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1345 = io_x[6] ? _GEN1344 : _GEN54;
wire  _GEN1346 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1347 = io_x[6] ? _GEN1346 : _GEN54;
wire  _GEN1348 = io_x[2] ? _GEN1347 : _GEN1345;
wire  _GEN1349 = io_x[14] ? _GEN1348 : _GEN1343;
wire  _GEN1350 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1351 = io_x[6] ? _GEN1350 : _GEN54;
wire  _GEN1352 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1353 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1354 = io_x[6] ? _GEN1353 : _GEN1352;
wire  _GEN1355 = io_x[2] ? _GEN1354 : _GEN1351;
wire  _GEN1356 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1357 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1358 = io_x[6] ? _GEN1357 : _GEN1356;
wire  _GEN1359 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1360 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1361 = io_x[6] ? _GEN1360 : _GEN1359;
wire  _GEN1362 = io_x[2] ? _GEN1361 : _GEN1358;
wire  _GEN1363 = io_x[14] ? _GEN1362 : _GEN1355;
wire  _GEN1364 = io_x[10] ? _GEN1363 : _GEN1349;
wire  _GEN1365 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1366 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1367 = io_x[6] ? _GEN1366 : _GEN1365;
wire  _GEN1368 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1369 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1370 = io_x[6] ? _GEN1369 : _GEN1368;
wire  _GEN1371 = io_x[2] ? _GEN1370 : _GEN1367;
wire  _GEN1372 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1373 = io_x[6] ? _GEN1372 : _GEN54;
wire  _GEN1374 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1375 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1376 = io_x[6] ? _GEN1375 : _GEN1374;
wire  _GEN1377 = io_x[2] ? _GEN1376 : _GEN1373;
wire  _GEN1378 = io_x[14] ? _GEN1377 : _GEN1371;
wire  _GEN1379 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1380 = io_x[6] ? _GEN1379 : _GEN54;
wire  _GEN1381 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1382 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1383 = io_x[6] ? _GEN1382 : _GEN1381;
wire  _GEN1384 = io_x[2] ? _GEN1383 : _GEN1380;
wire  _GEN1385 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1386 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1387 = io_x[6] ? _GEN1386 : _GEN1385;
wire  _GEN1388 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1389 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1390 = io_x[6] ? _GEN1389 : _GEN1388;
wire  _GEN1391 = io_x[2] ? _GEN1390 : _GEN1387;
wire  _GEN1392 = io_x[14] ? _GEN1391 : _GEN1384;
wire  _GEN1393 = io_x[10] ? _GEN1392 : _GEN1378;
wire  _GEN1394 = io_x[17] ? _GEN1393 : _GEN1364;
wire  _GEN1395 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1396 = io_x[6] ? _GEN1395 : _GEN298;
wire  _GEN1397 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN1398 = io_x[2] ? _GEN1397 : _GEN1396;
wire  _GEN1399 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1400 = io_x[6] ? _GEN1399 : _GEN54;
wire  _GEN1401 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1402 = io_x[6] ? _GEN1401 : _GEN298;
wire  _GEN1403 = io_x[2] ? _GEN1402 : _GEN1400;
wire  _GEN1404 = io_x[14] ? _GEN1403 : _GEN1398;
wire  _GEN1405 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1406 = io_x[6] ? _GEN1405 : _GEN298;
wire  _GEN1407 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1408 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1409 = io_x[6] ? _GEN1408 : _GEN1407;
wire  _GEN1410 = io_x[2] ? _GEN1409 : _GEN1406;
wire  _GEN1411 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1412 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1413 = io_x[6] ? _GEN1412 : _GEN1411;
wire  _GEN1414 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1415 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1416 = io_x[6] ? _GEN1415 : _GEN1414;
wire  _GEN1417 = io_x[2] ? _GEN1416 : _GEN1413;
wire  _GEN1418 = io_x[14] ? _GEN1417 : _GEN1410;
wire  _GEN1419 = io_x[10] ? _GEN1418 : _GEN1404;
wire  _GEN1420 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1421 = io_x[6] ? _GEN1420 : _GEN298;
wire  _GEN1422 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1423 = io_x[6] ? _GEN1422 : _GEN54;
wire  _GEN1424 = io_x[2] ? _GEN1423 : _GEN1421;
wire  _GEN1425 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1426 = io_x[6] ? _GEN1425 : _GEN54;
wire  _GEN1427 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1428 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1429 = io_x[6] ? _GEN1428 : _GEN1427;
wire  _GEN1430 = io_x[2] ? _GEN1429 : _GEN1426;
wire  _GEN1431 = io_x[14] ? _GEN1430 : _GEN1424;
wire  _GEN1432 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1433 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1434 = io_x[6] ? _GEN1433 : _GEN1432;
wire  _GEN1435 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1436 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1437 = io_x[6] ? _GEN1436 : _GEN1435;
wire  _GEN1438 = io_x[2] ? _GEN1437 : _GEN1434;
wire  _GEN1439 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1440 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1441 = io_x[6] ? _GEN1440 : _GEN1439;
wire  _GEN1442 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1443 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1444 = io_x[6] ? _GEN1443 : _GEN1442;
wire  _GEN1445 = io_x[2] ? _GEN1444 : _GEN1441;
wire  _GEN1446 = io_x[14] ? _GEN1445 : _GEN1438;
wire  _GEN1447 = io_x[10] ? _GEN1446 : _GEN1431;
wire  _GEN1448 = io_x[17] ? _GEN1447 : _GEN1419;
wire  _GEN1449 = io_x[25] ? _GEN1448 : _GEN1394;
wire  _GEN1450 = io_x[24] ? _GEN1449 : _GEN1337;
wire  _GEN1451 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN1452 = io_x[2] ? _GEN303 : _GEN1451;
wire  _GEN1453 = io_x[14] ? _GEN366 : _GEN1452;
wire  _GEN1454 = io_x[10] ? _GEN346 : _GEN1453;
wire  _GEN1455 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN1456 = io_x[2] ? _GEN358 : _GEN1455;
wire  _GEN1457 = io_x[6] ? _GEN54 : _GEN298;
wire  _GEN1458 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN1459 = io_x[2] ? _GEN1458 : _GEN1457;
wire  _GEN1460 = io_x[14] ? _GEN1459 : _GEN1456;
wire  _GEN1461 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1462 = io_x[6] ? _GEN1461 : _GEN298;
wire  _GEN1463 = io_x[2] ? _GEN1462 : _GEN303;
wire  _GEN1464 = io_x[14] ? _GEN1463 : _GEN366;
wire  _GEN1465 = io_x[10] ? _GEN1464 : _GEN1460;
wire  _GEN1466 = io_x[17] ? _GEN1465 : _GEN1454;
wire  _GEN1467 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1468 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1469 = io_x[6] ? _GEN1468 : _GEN1467;
wire  _GEN1470 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1471 = io_x[6] ? _GEN1470 : _GEN298;
wire  _GEN1472 = io_x[2] ? _GEN1471 : _GEN1469;
wire  _GEN1473 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1474 = io_x[6] ? _GEN1473 : _GEN298;
wire  _GEN1475 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1476 = io_x[6] ? _GEN1475 : _GEN54;
wire  _GEN1477 = io_x[2] ? _GEN1476 : _GEN1474;
wire  _GEN1478 = io_x[14] ? _GEN1477 : _GEN1472;
wire  _GEN1479 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1480 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1481 = io_x[6] ? _GEN1480 : _GEN1479;
wire  _GEN1482 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1483 = io_x[6] ? _GEN298 : _GEN1482;
wire  _GEN1484 = io_x[2] ? _GEN1483 : _GEN1481;
wire  _GEN1485 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1486 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1487 = io_x[6] ? _GEN1486 : _GEN1485;
wire  _GEN1488 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1489 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1490 = io_x[6] ? _GEN1489 : _GEN1488;
wire  _GEN1491 = io_x[2] ? _GEN1490 : _GEN1487;
wire  _GEN1492 = io_x[14] ? _GEN1491 : _GEN1484;
wire  _GEN1493 = io_x[10] ? _GEN1492 : _GEN1478;
wire  _GEN1494 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1495 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1496 = io_x[6] ? _GEN1495 : _GEN1494;
wire  _GEN1497 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1498 = io_x[6] ? _GEN1497 : _GEN298;
wire  _GEN1499 = io_x[2] ? _GEN1498 : _GEN1496;
wire  _GEN1500 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1501 = io_x[6] ? _GEN1500 : _GEN298;
wire  _GEN1502 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1503 = io_x[6] ? _GEN1502 : _GEN54;
wire  _GEN1504 = io_x[2] ? _GEN1503 : _GEN1501;
wire  _GEN1505 = io_x[14] ? _GEN1504 : _GEN1499;
wire  _GEN1506 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1507 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1508 = io_x[6] ? _GEN1507 : _GEN1506;
wire  _GEN1509 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1510 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1511 = io_x[6] ? _GEN1510 : _GEN1509;
wire  _GEN1512 = io_x[2] ? _GEN1511 : _GEN1508;
wire  _GEN1513 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1514 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1515 = io_x[6] ? _GEN1514 : _GEN1513;
wire  _GEN1516 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1517 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1518 = io_x[6] ? _GEN1517 : _GEN1516;
wire  _GEN1519 = io_x[2] ? _GEN1518 : _GEN1515;
wire  _GEN1520 = io_x[14] ? _GEN1519 : _GEN1512;
wire  _GEN1521 = io_x[10] ? _GEN1520 : _GEN1505;
wire  _GEN1522 = io_x[17] ? _GEN1521 : _GEN1493;
wire  _GEN1523 = io_x[25] ? _GEN1522 : _GEN1466;
wire  _GEN1524 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1525 = io_x[6] ? _GEN298 : _GEN1524;
wire  _GEN1526 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1527 = io_x[6] ? _GEN54 : _GEN1526;
wire  _GEN1528 = io_x[2] ? _GEN1527 : _GEN1525;
wire  _GEN1529 = io_x[14] ? _GEN366 : _GEN1528;
wire  _GEN1530 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1531 = io_x[6] ? _GEN1530 : _GEN54;
wire  _GEN1532 = io_x[2] ? _GEN358 : _GEN1531;
wire  _GEN1533 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1534 = io_x[6] ? _GEN1533 : _GEN54;
wire  _GEN1535 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1536 = io_x[6] ? _GEN1535 : _GEN54;
wire  _GEN1537 = io_x[2] ? _GEN1536 : _GEN1534;
wire  _GEN1538 = io_x[14] ? _GEN1537 : _GEN1532;
wire  _GEN1539 = io_x[10] ? _GEN1538 : _GEN1529;
wire  _GEN1540 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1541 = io_x[6] ? _GEN54 : _GEN1540;
wire  _GEN1542 = io_x[6] ? _GEN54 : _GEN298;
wire  _GEN1543 = io_x[2] ? _GEN1542 : _GEN1541;
wire  _GEN1544 = io_x[14] ? _GEN366 : _GEN1543;
wire  _GEN1545 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1546 = io_x[6] ? _GEN1545 : _GEN54;
wire  _GEN1547 = io_x[2] ? _GEN358 : _GEN1546;
wire  _GEN1548 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1549 = io_x[6] ? _GEN1548 : _GEN298;
wire  _GEN1550 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1551 = io_x[6] ? _GEN1550 : _GEN54;
wire  _GEN1552 = io_x[2] ? _GEN1551 : _GEN1549;
wire  _GEN1553 = io_x[14] ? _GEN1552 : _GEN1547;
wire  _GEN1554 = io_x[10] ? _GEN1553 : _GEN1544;
wire  _GEN1555 = io_x[17] ? _GEN1554 : _GEN1539;
wire  _GEN1556 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1557 = io_x[6] ? _GEN298 : _GEN1556;
wire  _GEN1558 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN1559 = io_x[2] ? _GEN1558 : _GEN1557;
wire  _GEN1560 = io_x[27] ? _GEN42 : _GEN43;
wire  _GEN1561 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1562 = io_x[6] ? _GEN1561 : _GEN1560;
wire  _GEN1563 = io_x[2] ? _GEN303 : _GEN1562;
wire  _GEN1564 = io_x[14] ? _GEN1563 : _GEN1559;
wire  _GEN1565 = io_x[2] ? _GEN358 : _GEN303;
wire  _GEN1566 = io_x[14] ? _GEN1565 : _GEN347;
wire  _GEN1567 = io_x[10] ? _GEN1566 : _GEN1564;
wire  _GEN1568 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1569 = io_x[6] ? _GEN298 : _GEN1568;
wire  _GEN1570 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1571 = io_x[6] ? _GEN1570 : _GEN54;
wire  _GEN1572 = io_x[2] ? _GEN1571 : _GEN1569;
wire  _GEN1573 = io_x[27] ? _GEN43 : _GEN42;
wire  _GEN1574 = io_x[6] ? _GEN1573 : _GEN298;
wire  _GEN1575 = io_x[2] ? _GEN303 : _GEN1574;
wire  _GEN1576 = io_x[14] ? _GEN1575 : _GEN1572;
wire  _GEN1577 = io_x[2] ? _GEN303 : _GEN358;
wire  _GEN1578 = io_x[6] ? _GEN54 : _GEN298;
wire  _GEN1579 = io_x[6] ? _GEN298 : _GEN54;
wire  _GEN1580 = io_x[2] ? _GEN1579 : _GEN1578;
wire  _GEN1581 = io_x[14] ? _GEN1580 : _GEN1577;
wire  _GEN1582 = io_x[10] ? _GEN1581 : _GEN1576;
wire  _GEN1583 = io_x[17] ? _GEN1582 : _GEN1567;
wire  _GEN1584 = io_x[25] ? _GEN1583 : _GEN1555;
wire  _GEN1585 = io_x[24] ? _GEN1584 : _GEN1523;
wire  _GEN1586 = io_x[32] ? _GEN1585 : _GEN1450;
wire  _GEN1587 = io_x[28] ? _GEN1586 : _GEN1222;
wire  _GEN1588 = io_x[26] ? _GEN1587 : _GEN792;
assign io_y[7] = _GEN1588;
wire  _GEN1589 = 1'b0;
wire  _GEN1590 = 1'b1;
wire  _GEN1591 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1592 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1593 = io_x[13] ? _GEN1592 : _GEN1591;
wire  _GEN1594 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1595 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1596 = io_x[13] ? _GEN1595 : _GEN1594;
wire  _GEN1597 = io_x[5] ? _GEN1596 : _GEN1593;
wire  _GEN1598 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1599 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1600 = io_x[13] ? _GEN1599 : _GEN1598;
wire  _GEN1601 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1602 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1603 = io_x[13] ? _GEN1602 : _GEN1601;
wire  _GEN1604 = io_x[5] ? _GEN1603 : _GEN1600;
wire  _GEN1605 = io_x[1] ? _GEN1604 : _GEN1597;
wire  _GEN1606 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1607 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1608 = io_x[13] ? _GEN1607 : _GEN1606;
wire  _GEN1609 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1610 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1611 = io_x[13] ? _GEN1610 : _GEN1609;
wire  _GEN1612 = io_x[5] ? _GEN1611 : _GEN1608;
wire  _GEN1613 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1614 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1615 = io_x[13] ? _GEN1614 : _GEN1613;
wire  _GEN1616 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1617 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1618 = io_x[13] ? _GEN1617 : _GEN1616;
wire  _GEN1619 = io_x[5] ? _GEN1618 : _GEN1615;
wire  _GEN1620 = io_x[1] ? _GEN1619 : _GEN1612;
wire  _GEN1621 = io_x[11] ? _GEN1620 : _GEN1605;
wire  _GEN1622 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1623 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1624 = io_x[13] ? _GEN1623 : _GEN1622;
wire  _GEN1625 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1626 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1627 = io_x[13] ? _GEN1626 : _GEN1625;
wire  _GEN1628 = io_x[5] ? _GEN1627 : _GEN1624;
wire  _GEN1629 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1630 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1631 = io_x[13] ? _GEN1630 : _GEN1629;
wire  _GEN1632 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1633 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1634 = io_x[13] ? _GEN1633 : _GEN1632;
wire  _GEN1635 = io_x[5] ? _GEN1634 : _GEN1631;
wire  _GEN1636 = io_x[1] ? _GEN1635 : _GEN1628;
wire  _GEN1637 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1638 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1639 = io_x[13] ? _GEN1638 : _GEN1637;
wire  _GEN1640 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1641 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1642 = io_x[13] ? _GEN1641 : _GEN1640;
wire  _GEN1643 = io_x[5] ? _GEN1642 : _GEN1639;
wire  _GEN1644 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1645 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1646 = io_x[13] ? _GEN1645 : _GEN1644;
wire  _GEN1647 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1648 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1649 = io_x[13] ? _GEN1648 : _GEN1647;
wire  _GEN1650 = io_x[5] ? _GEN1649 : _GEN1646;
wire  _GEN1651 = io_x[1] ? _GEN1650 : _GEN1643;
wire  _GEN1652 = io_x[11] ? _GEN1651 : _GEN1636;
wire  _GEN1653 = io_x[26] ? _GEN1652 : _GEN1621;
wire  _GEN1654 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1655 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1656 = io_x[13] ? _GEN1655 : _GEN1654;
wire  _GEN1657 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1658 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1659 = io_x[13] ? _GEN1658 : _GEN1657;
wire  _GEN1660 = io_x[5] ? _GEN1659 : _GEN1656;
wire  _GEN1661 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1662 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1663 = io_x[13] ? _GEN1662 : _GEN1661;
wire  _GEN1664 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1665 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1666 = io_x[13] ? _GEN1665 : _GEN1664;
wire  _GEN1667 = io_x[5] ? _GEN1666 : _GEN1663;
wire  _GEN1668 = io_x[1] ? _GEN1667 : _GEN1660;
wire  _GEN1669 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1670 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1671 = io_x[13] ? _GEN1670 : _GEN1669;
wire  _GEN1672 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1673 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1674 = io_x[13] ? _GEN1673 : _GEN1672;
wire  _GEN1675 = io_x[5] ? _GEN1674 : _GEN1671;
wire  _GEN1676 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1677 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1678 = io_x[13] ? _GEN1677 : _GEN1676;
wire  _GEN1679 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1680 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1681 = io_x[13] ? _GEN1680 : _GEN1679;
wire  _GEN1682 = io_x[5] ? _GEN1681 : _GEN1678;
wire  _GEN1683 = io_x[1] ? _GEN1682 : _GEN1675;
wire  _GEN1684 = io_x[11] ? _GEN1683 : _GEN1668;
wire  _GEN1685 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1686 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1687 = io_x[13] ? _GEN1686 : _GEN1685;
wire  _GEN1688 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1689 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1690 = io_x[13] ? _GEN1689 : _GEN1688;
wire  _GEN1691 = io_x[5] ? _GEN1690 : _GEN1687;
wire  _GEN1692 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1693 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1694 = io_x[13] ? _GEN1693 : _GEN1692;
wire  _GEN1695 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1696 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1697 = io_x[13] ? _GEN1696 : _GEN1695;
wire  _GEN1698 = io_x[5] ? _GEN1697 : _GEN1694;
wire  _GEN1699 = io_x[1] ? _GEN1698 : _GEN1691;
wire  _GEN1700 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1701 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1702 = io_x[13] ? _GEN1701 : _GEN1700;
wire  _GEN1703 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1704 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1705 = io_x[13] ? _GEN1704 : _GEN1703;
wire  _GEN1706 = io_x[5] ? _GEN1705 : _GEN1702;
wire  _GEN1707 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1708 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1709 = io_x[13] ? _GEN1708 : _GEN1707;
wire  _GEN1710 = io_x[9] ? _GEN1589 : _GEN1590;
wire  _GEN1711 = io_x[9] ? _GEN1590 : _GEN1589;
wire  _GEN1712 = io_x[13] ? _GEN1711 : _GEN1710;
wire  _GEN1713 = io_x[5] ? _GEN1712 : _GEN1709;
wire  _GEN1714 = io_x[1] ? _GEN1713 : _GEN1706;
wire  _GEN1715 = io_x[11] ? _GEN1714 : _GEN1699;
wire  _GEN1716 = io_x[26] ? _GEN1715 : _GEN1684;
wire  _GEN1717 = io_x[23] ? _GEN1716 : _GEN1653;
assign io_y[6] = _GEN1717;
wire  _GEN1718 = 1'b0;
wire  _GEN1719 = 1'b1;
wire  _GEN1720 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1721 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1722 = io_x[8] ? _GEN1721 : _GEN1720;
wire  _GEN1723 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1724 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1725 = io_x[8] ? _GEN1724 : _GEN1723;
wire  _GEN1726 = io_x[4] ? _GEN1725 : _GEN1722;
wire  _GEN1727 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1728 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1729 = io_x[8] ? _GEN1728 : _GEN1727;
wire  _GEN1730 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1731 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1732 = io_x[8] ? _GEN1731 : _GEN1730;
wire  _GEN1733 = io_x[4] ? _GEN1732 : _GEN1729;
wire  _GEN1734 = io_x[0] ? _GEN1733 : _GEN1726;
wire  _GEN1735 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1736 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1737 = io_x[8] ? _GEN1736 : _GEN1735;
wire  _GEN1738 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1739 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1740 = io_x[8] ? _GEN1739 : _GEN1738;
wire  _GEN1741 = io_x[4] ? _GEN1740 : _GEN1737;
wire  _GEN1742 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1743 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1744 = io_x[8] ? _GEN1743 : _GEN1742;
wire  _GEN1745 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1746 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1747 = io_x[8] ? _GEN1746 : _GEN1745;
wire  _GEN1748 = io_x[4] ? _GEN1747 : _GEN1744;
wire  _GEN1749 = io_x[0] ? _GEN1748 : _GEN1741;
wire  _GEN1750 = io_x[11] ? _GEN1749 : _GEN1734;
wire  _GEN1751 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1752 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1753 = io_x[8] ? _GEN1752 : _GEN1751;
wire  _GEN1754 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1755 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1756 = io_x[8] ? _GEN1755 : _GEN1754;
wire  _GEN1757 = io_x[4] ? _GEN1756 : _GEN1753;
wire  _GEN1758 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1759 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1760 = io_x[8] ? _GEN1759 : _GEN1758;
wire  _GEN1761 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1762 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1763 = io_x[8] ? _GEN1762 : _GEN1761;
wire  _GEN1764 = io_x[4] ? _GEN1763 : _GEN1760;
wire  _GEN1765 = io_x[0] ? _GEN1764 : _GEN1757;
wire  _GEN1766 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1767 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1768 = io_x[8] ? _GEN1767 : _GEN1766;
wire  _GEN1769 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1770 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1771 = io_x[8] ? _GEN1770 : _GEN1769;
wire  _GEN1772 = io_x[4] ? _GEN1771 : _GEN1768;
wire  _GEN1773 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1774 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1775 = io_x[8] ? _GEN1774 : _GEN1773;
wire  _GEN1776 = io_x[12] ? _GEN1718 : _GEN1719;
wire  _GEN1777 = io_x[12] ? _GEN1719 : _GEN1718;
wire  _GEN1778 = io_x[8] ? _GEN1777 : _GEN1776;
wire  _GEN1779 = io_x[4] ? _GEN1778 : _GEN1775;
wire  _GEN1780 = io_x[0] ? _GEN1779 : _GEN1772;
wire  _GEN1781 = io_x[11] ? _GEN1780 : _GEN1765;
wire  _GEN1782 = io_x[25] ? _GEN1781 : _GEN1750;
assign io_y[5] = _GEN1782;
wire  _GEN1783 = 1'b0;
wire  _GEN1784 = 1'b1;
wire  _GEN1785 = io_x[24] ? _GEN1784 : _GEN1783;
wire  _GEN1786 = io_x[24] ? _GEN1784 : _GEN1783;
wire  _GEN1787 = io_x[25] ? _GEN1786 : _GEN1785;
wire  _GEN1788 = io_x[24] ? _GEN1784 : _GEN1783;
wire  _GEN1789 = io_x[24] ? _GEN1784 : _GEN1783;
wire  _GEN1790 = io_x[25] ? _GEN1789 : _GEN1788;
wire  _GEN1791 = io_x[29] ? _GEN1790 : _GEN1787;
assign io_y[4] = _GEN1791;
wire  _GEN1792 = 1'b0;
wire  _GEN1793 = 1'b1;
wire  _GEN1794 = io_x[23] ? _GEN1793 : _GEN1792;
wire  _GEN1795 = io_x[23] ? _GEN1793 : _GEN1792;
wire  _GEN1796 = io_x[32] ? _GEN1795 : _GEN1794;
wire  _GEN1797 = io_x[23] ? _GEN1793 : _GEN1792;
wire  _GEN1798 = io_x[23] ? _GEN1793 : _GEN1792;
wire  _GEN1799 = io_x[32] ? _GEN1798 : _GEN1797;
wire  _GEN1800 = io_x[3] ? _GEN1799 : _GEN1796;
assign io_y[3] = _GEN1800;
wire  _GEN1801 = 1'b0;
wire  _GEN1802 = 1'b1;
wire  _GEN1803 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1804 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1805 = io_x[25] ? _GEN1804 : _GEN1803;
wire  _GEN1806 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1807 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1808 = io_x[25] ? _GEN1807 : _GEN1806;
wire  _GEN1809 = io_x[21] ? _GEN1808 : _GEN1805;
wire  _GEN1810 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1811 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1812 = io_x[25] ? _GEN1811 : _GEN1810;
wire  _GEN1813 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1814 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1815 = io_x[25] ? _GEN1814 : _GEN1813;
wire  _GEN1816 = io_x[21] ? _GEN1815 : _GEN1812;
wire  _GEN1817 = io_x[29] ? _GEN1816 : _GEN1809;
wire  _GEN1818 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1819 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1820 = io_x[25] ? _GEN1819 : _GEN1818;
wire  _GEN1821 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1822 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1823 = io_x[25] ? _GEN1822 : _GEN1821;
wire  _GEN1824 = io_x[21] ? _GEN1823 : _GEN1820;
wire  _GEN1825 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1826 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1827 = io_x[25] ? _GEN1826 : _GEN1825;
wire  _GEN1828 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1829 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1830 = io_x[25] ? _GEN1829 : _GEN1828;
wire  _GEN1831 = io_x[21] ? _GEN1830 : _GEN1827;
wire  _GEN1832 = io_x[29] ? _GEN1831 : _GEN1824;
wire  _GEN1833 = io_x[31] ? _GEN1832 : _GEN1817;
wire  _GEN1834 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1835 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1836 = io_x[25] ? _GEN1835 : _GEN1834;
wire  _GEN1837 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1838 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1839 = io_x[25] ? _GEN1838 : _GEN1837;
wire  _GEN1840 = io_x[21] ? _GEN1839 : _GEN1836;
wire  _GEN1841 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1842 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1843 = io_x[25] ? _GEN1842 : _GEN1841;
wire  _GEN1844 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1845 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1846 = io_x[25] ? _GEN1845 : _GEN1844;
wire  _GEN1847 = io_x[21] ? _GEN1846 : _GEN1843;
wire  _GEN1848 = io_x[29] ? _GEN1847 : _GEN1840;
wire  _GEN1849 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1850 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1851 = io_x[25] ? _GEN1850 : _GEN1849;
wire  _GEN1852 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1853 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1854 = io_x[25] ? _GEN1853 : _GEN1852;
wire  _GEN1855 = io_x[21] ? _GEN1854 : _GEN1851;
wire  _GEN1856 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1857 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1858 = io_x[25] ? _GEN1857 : _GEN1856;
wire  _GEN1859 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1860 = io_x[22] ? _GEN1802 : _GEN1801;
wire  _GEN1861 = io_x[25] ? _GEN1860 : _GEN1859;
wire  _GEN1862 = io_x[21] ? _GEN1861 : _GEN1858;
wire  _GEN1863 = io_x[29] ? _GEN1862 : _GEN1855;
wire  _GEN1864 = io_x[31] ? _GEN1863 : _GEN1848;
wire  _GEN1865 = io_x[28] ? _GEN1864 : _GEN1833;
assign io_y[2] = _GEN1865;
wire  _GEN1866 = 1'b0;
wire  _GEN1867 = 1'b1;
wire  _GEN1868 = io_x[21] ? _GEN1867 : _GEN1866;
wire  _GEN1869 = io_x[21] ? _GEN1867 : _GEN1866;
wire  _GEN1870 = io_x[20] ? _GEN1869 : _GEN1868;
assign io_y[1] = _GEN1870;
wire  _GEN1871 = 1'b0;
wire  _GEN1872 = 1'b1;
wire  _GEN1873 = io_x[20] ? _GEN1872 : _GEN1871;
wire  _GEN1874 = io_x[20] ? _GEN1872 : _GEN1871;
wire  _GEN1875 = io_x[23] ? _GEN1874 : _GEN1873;
assign io_y[0] = _GEN1875;
endmodule
module BBGSharePredictorImp_BSD_NutShell_train(
    input [31:0] train_pc,
    input  train_taken,
    input [15:0] train_ghr_rdata,
    output  pht_wdata,
    output [8:0] pht_waddr,
    output  ghr_wdata
);
wire [48:0] io_x;
wire [10:0] io_y;
assign io_x = { train_pc, train_taken, train_ghr_rdata };
assign { pht_wdata, pht_waddr, ghr_wdata } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN3 = io_x[16] ? _GEN1 : _GEN0;
wire  _GEN4 = io_x[26] ? _GEN3 : _GEN2;
assign io_y[10] = _GEN4;
wire  _GEN5 = 1'b0;
wire  _GEN6 = 1'b1;
wire  _GEN7 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN8 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN9 = io_x[7] ? _GEN8 : _GEN7;
wire  _GEN10 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN11 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN12 = io_x[7] ? _GEN11 : _GEN10;
wire  _GEN13 = io_x[11] ? _GEN12 : _GEN9;
wire  _GEN14 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN15 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN16 = io_x[7] ? _GEN15 : _GEN14;
wire  _GEN17 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN18 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN19 = io_x[7] ? _GEN18 : _GEN17;
wire  _GEN20 = io_x[11] ? _GEN19 : _GEN16;
wire  _GEN21 = io_x[1] ? _GEN20 : _GEN13;
wire  _GEN22 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN23 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN24 = io_x[7] ? _GEN23 : _GEN22;
wire  _GEN25 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN26 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN27 = io_x[7] ? _GEN26 : _GEN25;
wire  _GEN28 = io_x[11] ? _GEN27 : _GEN24;
wire  _GEN29 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN30 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN31 = io_x[7] ? _GEN30 : _GEN29;
wire  _GEN32 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN33 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN34 = io_x[7] ? _GEN33 : _GEN32;
wire  _GEN35 = io_x[11] ? _GEN34 : _GEN31;
wire  _GEN36 = io_x[1] ? _GEN35 : _GEN28;
wire  _GEN37 = io_x[27] ? _GEN36 : _GEN21;
wire  _GEN38 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN39 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN40 = io_x[7] ? _GEN39 : _GEN38;
wire  _GEN41 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN42 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN43 = io_x[7] ? _GEN42 : _GEN41;
wire  _GEN44 = io_x[11] ? _GEN43 : _GEN40;
wire  _GEN45 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN46 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN47 = io_x[7] ? _GEN46 : _GEN45;
wire  _GEN48 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN49 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN50 = io_x[7] ? _GEN49 : _GEN48;
wire  _GEN51 = io_x[11] ? _GEN50 : _GEN47;
wire  _GEN52 = io_x[1] ? _GEN51 : _GEN44;
wire  _GEN53 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN54 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN55 = io_x[7] ? _GEN54 : _GEN53;
wire  _GEN56 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN57 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN58 = io_x[7] ? _GEN57 : _GEN56;
wire  _GEN59 = io_x[11] ? _GEN58 : _GEN55;
wire  _GEN60 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN61 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN62 = io_x[7] ? _GEN61 : _GEN60;
wire  _GEN63 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN64 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN65 = io_x[7] ? _GEN64 : _GEN63;
wire  _GEN66 = io_x[11] ? _GEN65 : _GEN62;
wire  _GEN67 = io_x[1] ? _GEN66 : _GEN59;
wire  _GEN68 = io_x[27] ? _GEN67 : _GEN52;
wire  _GEN69 = io_x[15] ? _GEN68 : _GEN37;
wire  _GEN70 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN71 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN72 = io_x[7] ? _GEN71 : _GEN70;
wire  _GEN73 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN74 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN75 = io_x[7] ? _GEN74 : _GEN73;
wire  _GEN76 = io_x[11] ? _GEN75 : _GEN72;
wire  _GEN77 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN78 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN79 = io_x[7] ? _GEN78 : _GEN77;
wire  _GEN80 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN81 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN82 = io_x[7] ? _GEN81 : _GEN80;
wire  _GEN83 = io_x[11] ? _GEN82 : _GEN79;
wire  _GEN84 = io_x[1] ? _GEN83 : _GEN76;
wire  _GEN85 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN86 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN87 = io_x[7] ? _GEN86 : _GEN85;
wire  _GEN88 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN89 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN90 = io_x[7] ? _GEN89 : _GEN88;
wire  _GEN91 = io_x[11] ? _GEN90 : _GEN87;
wire  _GEN92 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN93 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN94 = io_x[7] ? _GEN93 : _GEN92;
wire  _GEN95 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN96 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN97 = io_x[7] ? _GEN96 : _GEN95;
wire  _GEN98 = io_x[11] ? _GEN97 : _GEN94;
wire  _GEN99 = io_x[1] ? _GEN98 : _GEN91;
wire  _GEN100 = io_x[27] ? _GEN99 : _GEN84;
wire  _GEN101 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN102 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN103 = io_x[7] ? _GEN102 : _GEN101;
wire  _GEN104 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN105 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN106 = io_x[7] ? _GEN105 : _GEN104;
wire  _GEN107 = io_x[11] ? _GEN106 : _GEN103;
wire  _GEN108 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN109 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN110 = io_x[7] ? _GEN109 : _GEN108;
wire  _GEN111 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN112 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN113 = io_x[7] ? _GEN112 : _GEN111;
wire  _GEN114 = io_x[11] ? _GEN113 : _GEN110;
wire  _GEN115 = io_x[1] ? _GEN114 : _GEN107;
wire  _GEN116 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN117 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN118 = io_x[7] ? _GEN117 : _GEN116;
wire  _GEN119 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN120 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN121 = io_x[7] ? _GEN120 : _GEN119;
wire  _GEN122 = io_x[11] ? _GEN121 : _GEN118;
wire  _GEN123 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN124 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN125 = io_x[7] ? _GEN124 : _GEN123;
wire  _GEN126 = io_x[3] ? _GEN5 : _GEN6;
wire  _GEN127 = io_x[3] ? _GEN6 : _GEN5;
wire  _GEN128 = io_x[7] ? _GEN127 : _GEN126;
wire  _GEN129 = io_x[11] ? _GEN128 : _GEN125;
wire  _GEN130 = io_x[1] ? _GEN129 : _GEN122;
wire  _GEN131 = io_x[27] ? _GEN130 : _GEN115;
wire  _GEN132 = io_x[15] ? _GEN131 : _GEN100;
wire  _GEN133 = io_x[16] ? _GEN132 : _GEN69;
assign io_y[9] = _GEN133;
wire  _GEN134 = 1'b0;
wire  _GEN135 = 1'b1;
wire  _GEN136 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN137 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN138 = io_x[10] ? _GEN137 : _GEN136;
wire  _GEN139 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN140 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN141 = io_x[10] ? _GEN140 : _GEN139;
wire  _GEN142 = io_x[14] ? _GEN141 : _GEN138;
wire  _GEN143 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN144 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN145 = io_x[10] ? _GEN144 : _GEN143;
wire  _GEN146 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN147 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN148 = io_x[10] ? _GEN147 : _GEN146;
wire  _GEN149 = io_x[14] ? _GEN148 : _GEN145;
wire  _GEN150 = io_x[2] ? _GEN149 : _GEN142;
wire  _GEN151 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN152 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN153 = io_x[10] ? _GEN152 : _GEN151;
wire  _GEN154 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN155 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN156 = io_x[10] ? _GEN155 : _GEN154;
wire  _GEN157 = io_x[14] ? _GEN156 : _GEN153;
wire  _GEN158 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN159 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN160 = io_x[10] ? _GEN159 : _GEN158;
wire  _GEN161 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN162 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN163 = io_x[10] ? _GEN162 : _GEN161;
wire  _GEN164 = io_x[14] ? _GEN163 : _GEN160;
wire  _GEN165 = io_x[2] ? _GEN164 : _GEN157;
wire  _GEN166 = io_x[26] ? _GEN165 : _GEN150;
wire  _GEN167 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN168 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN169 = io_x[10] ? _GEN168 : _GEN167;
wire  _GEN170 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN171 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN172 = io_x[10] ? _GEN171 : _GEN170;
wire  _GEN173 = io_x[14] ? _GEN172 : _GEN169;
wire  _GEN174 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN175 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN176 = io_x[10] ? _GEN175 : _GEN174;
wire  _GEN177 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN178 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN179 = io_x[10] ? _GEN178 : _GEN177;
wire  _GEN180 = io_x[14] ? _GEN179 : _GEN176;
wire  _GEN181 = io_x[2] ? _GEN180 : _GEN173;
wire  _GEN182 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN183 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN184 = io_x[10] ? _GEN183 : _GEN182;
wire  _GEN185 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN186 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN187 = io_x[10] ? _GEN186 : _GEN185;
wire  _GEN188 = io_x[14] ? _GEN187 : _GEN184;
wire  _GEN189 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN190 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN191 = io_x[10] ? _GEN190 : _GEN189;
wire  _GEN192 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN193 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN194 = io_x[10] ? _GEN193 : _GEN192;
wire  _GEN195 = io_x[14] ? _GEN194 : _GEN191;
wire  _GEN196 = io_x[2] ? _GEN195 : _GEN188;
wire  _GEN197 = io_x[26] ? _GEN196 : _GEN181;
wire  _GEN198 = io_x[5] ? _GEN197 : _GEN166;
wire  _GEN199 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN200 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN201 = io_x[10] ? _GEN200 : _GEN199;
wire  _GEN202 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN203 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN204 = io_x[10] ? _GEN203 : _GEN202;
wire  _GEN205 = io_x[14] ? _GEN204 : _GEN201;
wire  _GEN206 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN207 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN208 = io_x[10] ? _GEN207 : _GEN206;
wire  _GEN209 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN210 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN211 = io_x[10] ? _GEN210 : _GEN209;
wire  _GEN212 = io_x[14] ? _GEN211 : _GEN208;
wire  _GEN213 = io_x[2] ? _GEN212 : _GEN205;
wire  _GEN214 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN215 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN216 = io_x[10] ? _GEN215 : _GEN214;
wire  _GEN217 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN218 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN219 = io_x[10] ? _GEN218 : _GEN217;
wire  _GEN220 = io_x[14] ? _GEN219 : _GEN216;
wire  _GEN221 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN222 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN223 = io_x[10] ? _GEN222 : _GEN221;
wire  _GEN224 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN225 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN226 = io_x[10] ? _GEN225 : _GEN224;
wire  _GEN227 = io_x[14] ? _GEN226 : _GEN223;
wire  _GEN228 = io_x[2] ? _GEN227 : _GEN220;
wire  _GEN229 = io_x[26] ? _GEN228 : _GEN213;
wire  _GEN230 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN231 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN232 = io_x[10] ? _GEN231 : _GEN230;
wire  _GEN233 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN234 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN235 = io_x[10] ? _GEN234 : _GEN233;
wire  _GEN236 = io_x[14] ? _GEN235 : _GEN232;
wire  _GEN237 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN238 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN239 = io_x[10] ? _GEN238 : _GEN237;
wire  _GEN240 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN241 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN242 = io_x[10] ? _GEN241 : _GEN240;
wire  _GEN243 = io_x[14] ? _GEN242 : _GEN239;
wire  _GEN244 = io_x[2] ? _GEN243 : _GEN236;
wire  _GEN245 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN246 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN247 = io_x[10] ? _GEN246 : _GEN245;
wire  _GEN248 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN249 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN250 = io_x[10] ? _GEN249 : _GEN248;
wire  _GEN251 = io_x[14] ? _GEN250 : _GEN247;
wire  _GEN252 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN253 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN254 = io_x[10] ? _GEN253 : _GEN252;
wire  _GEN255 = io_x[6] ? _GEN134 : _GEN135;
wire  _GEN256 = io_x[6] ? _GEN135 : _GEN134;
wire  _GEN257 = io_x[10] ? _GEN256 : _GEN255;
wire  _GEN258 = io_x[14] ? _GEN257 : _GEN254;
wire  _GEN259 = io_x[2] ? _GEN258 : _GEN251;
wire  _GEN260 = io_x[26] ? _GEN259 : _GEN244;
wire  _GEN261 = io_x[5] ? _GEN260 : _GEN229;
wire  _GEN262 = io_x[16] ? _GEN261 : _GEN198;
assign io_y[8] = _GEN262;
wire  _GEN263 = 1'b1;
wire  _GEN264 = 1'b0;
wire  _GEN265 = 1'b1;
wire  _GEN266 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN267 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN268 = io_x[9] ? _GEN267 : _GEN266;
wire  _GEN269 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN270 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN271 = io_x[9] ? _GEN270 : _GEN269;
wire  _GEN272 = io_x[13] ? _GEN271 : _GEN268;
wire  _GEN273 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN274 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN275 = io_x[9] ? _GEN274 : _GEN273;
wire  _GEN276 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN277 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN278 = io_x[9] ? _GEN277 : _GEN276;
wire  _GEN279 = io_x[13] ? _GEN278 : _GEN275;
wire  _GEN280 = io_x[1] ? _GEN279 : _GEN272;
wire  _GEN281 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN282 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN283 = io_x[9] ? _GEN282 : _GEN281;
wire  _GEN284 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN285 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN286 = io_x[9] ? _GEN285 : _GEN284;
wire  _GEN287 = io_x[13] ? _GEN286 : _GEN283;
wire  _GEN288 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN289 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN290 = io_x[9] ? _GEN289 : _GEN288;
wire  _GEN291 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN292 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN293 = io_x[9] ? _GEN292 : _GEN291;
wire  _GEN294 = io_x[13] ? _GEN293 : _GEN290;
wire  _GEN295 = io_x[1] ? _GEN294 : _GEN287;
wire  _GEN296 = io_x[0] ? _GEN295 : _GEN280;
wire  _GEN297 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN298 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN299 = io_x[9] ? _GEN298 : _GEN297;
wire  _GEN300 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN301 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN302 = io_x[9] ? _GEN301 : _GEN300;
wire  _GEN303 = io_x[13] ? _GEN302 : _GEN299;
wire  _GEN304 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN305 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN306 = io_x[9] ? _GEN305 : _GEN304;
wire  _GEN307 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN308 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN309 = io_x[9] ? _GEN308 : _GEN307;
wire  _GEN310 = io_x[13] ? _GEN309 : _GEN306;
wire  _GEN311 = io_x[1] ? _GEN310 : _GEN303;
wire  _GEN312 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN313 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN314 = io_x[9] ? _GEN313 : _GEN312;
wire  _GEN315 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN316 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN317 = io_x[9] ? _GEN316 : _GEN315;
wire  _GEN318 = io_x[13] ? _GEN317 : _GEN314;
wire  _GEN319 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN320 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN321 = io_x[9] ? _GEN320 : _GEN319;
wire  _GEN322 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN323 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN324 = io_x[9] ? _GEN323 : _GEN322;
wire  _GEN325 = io_x[13] ? _GEN324 : _GEN321;
wire  _GEN326 = io_x[1] ? _GEN325 : _GEN318;
wire  _GEN327 = io_x[0] ? _GEN326 : _GEN311;
wire  _GEN328 = io_x[31] ? _GEN327 : _GEN296;
wire  _GEN329 = 1'b1;
wire  _GEN330 = io_x[32] ? _GEN329 : _GEN328;
wire  _GEN331 = 1'b1;
wire  _GEN332 = io_x[33] ? _GEN331 : _GEN330;
wire  _GEN333 = 1'b1;
wire  _GEN334 = io_x[34] ? _GEN333 : _GEN332;
wire  _GEN335 = 1'b1;
wire  _GEN336 = io_x[35] ? _GEN335 : _GEN334;
wire  _GEN337 = 1'b1;
wire  _GEN338 = io_x[36] ? _GEN337 : _GEN336;
wire  _GEN339 = 1'b1;
wire  _GEN340 = io_x[37] ? _GEN339 : _GEN338;
wire  _GEN341 = 1'b1;
wire  _GEN342 = io_x[38] ? _GEN341 : _GEN340;
wire  _GEN343 = 1'b1;
wire  _GEN344 = io_x[39] ? _GEN343 : _GEN342;
wire  _GEN345 = 1'b1;
wire  _GEN346 = io_x[40] ? _GEN345 : _GEN344;
wire  _GEN347 = 1'b1;
wire  _GEN348 = io_x[41] ? _GEN347 : _GEN346;
wire  _GEN349 = 1'b1;
wire  _GEN350 = io_x[42] ? _GEN349 : _GEN348;
wire  _GEN351 = 1'b1;
wire  _GEN352 = io_x[43] ? _GEN351 : _GEN350;
wire  _GEN353 = 1'b1;
wire  _GEN354 = io_x[44] ? _GEN353 : _GEN352;
wire  _GEN355 = 1'b1;
wire  _GEN356 = io_x[45] ? _GEN355 : _GEN354;
wire  _GEN357 = 1'b1;
wire  _GEN358 = io_x[46] ? _GEN357 : _GEN356;
wire  _GEN359 = 1'b1;
wire  _GEN360 = io_x[47] ? _GEN359 : _GEN358;
wire  _GEN361 = io_x[48] ? _GEN360 : _GEN263;
wire  _GEN362 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN363 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN364 = io_x[9] ? _GEN363 : _GEN362;
wire  _GEN365 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN366 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN367 = io_x[9] ? _GEN366 : _GEN365;
wire  _GEN368 = io_x[13] ? _GEN367 : _GEN364;
wire  _GEN369 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN370 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN371 = io_x[9] ? _GEN370 : _GEN369;
wire  _GEN372 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN373 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN374 = io_x[9] ? _GEN373 : _GEN372;
wire  _GEN375 = io_x[13] ? _GEN374 : _GEN371;
wire  _GEN376 = io_x[1] ? _GEN375 : _GEN368;
wire  _GEN377 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN378 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN379 = io_x[9] ? _GEN378 : _GEN377;
wire  _GEN380 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN381 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN382 = io_x[9] ? _GEN381 : _GEN380;
wire  _GEN383 = io_x[13] ? _GEN382 : _GEN379;
wire  _GEN384 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN385 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN386 = io_x[9] ? _GEN385 : _GEN384;
wire  _GEN387 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN388 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN389 = io_x[9] ? _GEN388 : _GEN387;
wire  _GEN390 = io_x[13] ? _GEN389 : _GEN386;
wire  _GEN391 = io_x[1] ? _GEN390 : _GEN383;
wire  _GEN392 = io_x[0] ? _GEN391 : _GEN376;
wire  _GEN393 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN394 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN395 = io_x[9] ? _GEN394 : _GEN393;
wire  _GEN396 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN397 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN398 = io_x[9] ? _GEN397 : _GEN396;
wire  _GEN399 = io_x[13] ? _GEN398 : _GEN395;
wire  _GEN400 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN401 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN402 = io_x[9] ? _GEN401 : _GEN400;
wire  _GEN403 = 1'b0;
wire  _GEN404 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN405 = io_x[9] ? _GEN404 : _GEN403;
wire  _GEN406 = io_x[13] ? _GEN405 : _GEN402;
wire  _GEN407 = io_x[1] ? _GEN406 : _GEN399;
wire  _GEN408 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN409 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN410 = io_x[9] ? _GEN409 : _GEN408;
wire  _GEN411 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN412 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN413 = io_x[9] ? _GEN412 : _GEN411;
wire  _GEN414 = io_x[13] ? _GEN413 : _GEN410;
wire  _GEN415 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN416 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN417 = io_x[9] ? _GEN416 : _GEN415;
wire  _GEN418 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN419 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN420 = io_x[9] ? _GEN419 : _GEN418;
wire  _GEN421 = io_x[13] ? _GEN420 : _GEN417;
wire  _GEN422 = io_x[1] ? _GEN421 : _GEN414;
wire  _GEN423 = io_x[0] ? _GEN422 : _GEN407;
wire  _GEN424 = io_x[31] ? _GEN423 : _GEN392;
wire  _GEN425 = io_x[32] ? _GEN329 : _GEN424;
wire  _GEN426 = io_x[33] ? _GEN331 : _GEN425;
wire  _GEN427 = io_x[34] ? _GEN333 : _GEN426;
wire  _GEN428 = io_x[35] ? _GEN335 : _GEN427;
wire  _GEN429 = io_x[36] ? _GEN337 : _GEN428;
wire  _GEN430 = io_x[37] ? _GEN339 : _GEN429;
wire  _GEN431 = io_x[38] ? _GEN341 : _GEN430;
wire  _GEN432 = io_x[39] ? _GEN343 : _GEN431;
wire  _GEN433 = io_x[40] ? _GEN345 : _GEN432;
wire  _GEN434 = io_x[41] ? _GEN347 : _GEN433;
wire  _GEN435 = io_x[42] ? _GEN349 : _GEN434;
wire  _GEN436 = io_x[43] ? _GEN351 : _GEN435;
wire  _GEN437 = io_x[44] ? _GEN353 : _GEN436;
wire  _GEN438 = io_x[45] ? _GEN355 : _GEN437;
wire  _GEN439 = io_x[46] ? _GEN357 : _GEN438;
wire  _GEN440 = io_x[47] ? _GEN359 : _GEN439;
wire  _GEN441 = io_x[48] ? _GEN440 : _GEN263;
wire  _GEN442 = io_x[25] ? _GEN441 : _GEN361;
wire  _GEN443 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN444 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN445 = io_x[9] ? _GEN444 : _GEN443;
wire  _GEN446 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN447 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN448 = io_x[9] ? _GEN447 : _GEN446;
wire  _GEN449 = io_x[13] ? _GEN448 : _GEN445;
wire  _GEN450 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN451 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN452 = io_x[9] ? _GEN451 : _GEN450;
wire  _GEN453 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN454 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN455 = io_x[9] ? _GEN454 : _GEN453;
wire  _GEN456 = io_x[13] ? _GEN455 : _GEN452;
wire  _GEN457 = io_x[1] ? _GEN456 : _GEN449;
wire  _GEN458 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN459 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN460 = io_x[9] ? _GEN459 : _GEN458;
wire  _GEN461 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN462 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN463 = io_x[9] ? _GEN462 : _GEN461;
wire  _GEN464 = io_x[13] ? _GEN463 : _GEN460;
wire  _GEN465 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN466 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN467 = io_x[9] ? _GEN466 : _GEN465;
wire  _GEN468 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN469 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN470 = io_x[9] ? _GEN469 : _GEN468;
wire  _GEN471 = io_x[13] ? _GEN470 : _GEN467;
wire  _GEN472 = io_x[1] ? _GEN471 : _GEN464;
wire  _GEN473 = io_x[0] ? _GEN472 : _GEN457;
wire  _GEN474 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN475 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN476 = io_x[9] ? _GEN475 : _GEN474;
wire  _GEN477 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN478 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN479 = io_x[9] ? _GEN478 : _GEN477;
wire  _GEN480 = io_x[13] ? _GEN479 : _GEN476;
wire  _GEN481 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN482 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN483 = io_x[9] ? _GEN482 : _GEN481;
wire  _GEN484 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN485 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN486 = io_x[9] ? _GEN485 : _GEN484;
wire  _GEN487 = io_x[13] ? _GEN486 : _GEN483;
wire  _GEN488 = io_x[1] ? _GEN487 : _GEN480;
wire  _GEN489 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN490 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN491 = io_x[9] ? _GEN490 : _GEN489;
wire  _GEN492 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN493 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN494 = io_x[9] ? _GEN493 : _GEN492;
wire  _GEN495 = io_x[13] ? _GEN494 : _GEN491;
wire  _GEN496 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN497 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN498 = io_x[9] ? _GEN497 : _GEN496;
wire  _GEN499 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN500 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN501 = io_x[9] ? _GEN500 : _GEN499;
wire  _GEN502 = io_x[13] ? _GEN501 : _GEN498;
wire  _GEN503 = io_x[1] ? _GEN502 : _GEN495;
wire  _GEN504 = io_x[0] ? _GEN503 : _GEN488;
wire  _GEN505 = io_x[31] ? _GEN504 : _GEN473;
wire  _GEN506 = io_x[32] ? _GEN329 : _GEN505;
wire  _GEN507 = io_x[33] ? _GEN331 : _GEN506;
wire  _GEN508 = io_x[34] ? _GEN333 : _GEN507;
wire  _GEN509 = io_x[35] ? _GEN335 : _GEN508;
wire  _GEN510 = io_x[36] ? _GEN337 : _GEN509;
wire  _GEN511 = io_x[37] ? _GEN339 : _GEN510;
wire  _GEN512 = io_x[38] ? _GEN341 : _GEN511;
wire  _GEN513 = io_x[39] ? _GEN343 : _GEN512;
wire  _GEN514 = io_x[40] ? _GEN345 : _GEN513;
wire  _GEN515 = io_x[41] ? _GEN347 : _GEN514;
wire  _GEN516 = io_x[42] ? _GEN349 : _GEN515;
wire  _GEN517 = io_x[43] ? _GEN351 : _GEN516;
wire  _GEN518 = io_x[44] ? _GEN353 : _GEN517;
wire  _GEN519 = io_x[45] ? _GEN355 : _GEN518;
wire  _GEN520 = io_x[46] ? _GEN357 : _GEN519;
wire  _GEN521 = io_x[47] ? _GEN359 : _GEN520;
wire  _GEN522 = io_x[48] ? _GEN521 : _GEN263;
wire  _GEN523 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN524 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN525 = io_x[9] ? _GEN524 : _GEN523;
wire  _GEN526 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN527 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN528 = io_x[9] ? _GEN527 : _GEN526;
wire  _GEN529 = io_x[13] ? _GEN528 : _GEN525;
wire  _GEN530 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN531 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN532 = io_x[9] ? _GEN531 : _GEN530;
wire  _GEN533 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN534 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN535 = io_x[9] ? _GEN534 : _GEN533;
wire  _GEN536 = io_x[13] ? _GEN535 : _GEN532;
wire  _GEN537 = io_x[1] ? _GEN536 : _GEN529;
wire  _GEN538 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN539 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN540 = io_x[9] ? _GEN539 : _GEN538;
wire  _GEN541 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN542 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN543 = io_x[9] ? _GEN542 : _GEN541;
wire  _GEN544 = io_x[13] ? _GEN543 : _GEN540;
wire  _GEN545 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN546 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN547 = io_x[9] ? _GEN546 : _GEN545;
wire  _GEN548 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN549 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN550 = io_x[9] ? _GEN549 : _GEN548;
wire  _GEN551 = io_x[13] ? _GEN550 : _GEN547;
wire  _GEN552 = io_x[1] ? _GEN551 : _GEN544;
wire  _GEN553 = io_x[0] ? _GEN552 : _GEN537;
wire  _GEN554 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN555 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN556 = io_x[9] ? _GEN555 : _GEN554;
wire  _GEN557 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN558 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN559 = io_x[9] ? _GEN558 : _GEN557;
wire  _GEN560 = io_x[13] ? _GEN559 : _GEN556;
wire  _GEN561 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN562 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN563 = io_x[9] ? _GEN562 : _GEN561;
wire  _GEN564 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN565 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN566 = io_x[9] ? _GEN565 : _GEN564;
wire  _GEN567 = io_x[13] ? _GEN566 : _GEN563;
wire  _GEN568 = io_x[1] ? _GEN567 : _GEN560;
wire  _GEN569 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN570 = 1'b1;
wire  _GEN571 = io_x[9] ? _GEN570 : _GEN569;
wire  _GEN572 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN573 = io_x[9] ? _GEN572 : _GEN570;
wire  _GEN574 = io_x[13] ? _GEN573 : _GEN571;
wire  _GEN575 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN576 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN577 = io_x[9] ? _GEN576 : _GEN575;
wire  _GEN578 = io_x[5] ? _GEN264 : _GEN265;
wire  _GEN579 = io_x[5] ? _GEN265 : _GEN264;
wire  _GEN580 = io_x[9] ? _GEN579 : _GEN578;
wire  _GEN581 = io_x[13] ? _GEN580 : _GEN577;
wire  _GEN582 = io_x[1] ? _GEN581 : _GEN574;
wire  _GEN583 = io_x[0] ? _GEN582 : _GEN568;
wire  _GEN584 = io_x[31] ? _GEN583 : _GEN553;
wire  _GEN585 = io_x[32] ? _GEN329 : _GEN584;
wire  _GEN586 = io_x[33] ? _GEN331 : _GEN585;
wire  _GEN587 = io_x[34] ? _GEN333 : _GEN586;
wire  _GEN588 = io_x[35] ? _GEN335 : _GEN587;
wire  _GEN589 = io_x[36] ? _GEN337 : _GEN588;
wire  _GEN590 = io_x[37] ? _GEN339 : _GEN589;
wire  _GEN591 = io_x[38] ? _GEN341 : _GEN590;
wire  _GEN592 = io_x[39] ? _GEN343 : _GEN591;
wire  _GEN593 = io_x[40] ? _GEN345 : _GEN592;
wire  _GEN594 = io_x[41] ? _GEN347 : _GEN593;
wire  _GEN595 = io_x[42] ? _GEN349 : _GEN594;
wire  _GEN596 = io_x[43] ? _GEN351 : _GEN595;
wire  _GEN597 = io_x[44] ? _GEN353 : _GEN596;
wire  _GEN598 = io_x[45] ? _GEN355 : _GEN597;
wire  _GEN599 = io_x[46] ? _GEN357 : _GEN598;
wire  _GEN600 = io_x[47] ? _GEN359 : _GEN599;
wire  _GEN601 = io_x[48] ? _GEN600 : _GEN263;
wire  _GEN602 = io_x[25] ? _GEN601 : _GEN522;
wire  _GEN603 = io_x[22] ? _GEN602 : _GEN442;
assign io_y[7] = _GEN603;
wire  _GEN604 = 1'b0;
wire  _GEN605 = 1'b1;
wire  _GEN606 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN607 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN608 = io_x[24] ? _GEN607 : _GEN606;
wire  _GEN609 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN610 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN611 = io_x[24] ? _GEN610 : _GEN609;
wire  _GEN612 = io_x[26] ? _GEN611 : _GEN608;
wire  _GEN613 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN614 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN615 = io_x[24] ? _GEN614 : _GEN613;
wire  _GEN616 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN617 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN618 = io_x[24] ? _GEN617 : _GEN616;
wire  _GEN619 = io_x[26] ? _GEN618 : _GEN615;
wire  _GEN620 = io_x[3] ? _GEN619 : _GEN612;
wire  _GEN621 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN622 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN623 = io_x[24] ? _GEN622 : _GEN621;
wire  _GEN624 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN625 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN626 = io_x[24] ? _GEN625 : _GEN624;
wire  _GEN627 = io_x[26] ? _GEN626 : _GEN623;
wire  _GEN628 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN629 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN630 = io_x[24] ? _GEN629 : _GEN628;
wire  _GEN631 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN632 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN633 = io_x[24] ? _GEN632 : _GEN631;
wire  _GEN634 = io_x[26] ? _GEN633 : _GEN630;
wire  _GEN635 = io_x[3] ? _GEN634 : _GEN627;
wire  _GEN636 = io_x[8] ? _GEN635 : _GEN620;
wire  _GEN637 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN638 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN639 = io_x[24] ? _GEN638 : _GEN637;
wire  _GEN640 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN641 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN642 = io_x[24] ? _GEN641 : _GEN640;
wire  _GEN643 = io_x[26] ? _GEN642 : _GEN639;
wire  _GEN644 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN645 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN646 = io_x[24] ? _GEN645 : _GEN644;
wire  _GEN647 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN648 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN649 = io_x[24] ? _GEN648 : _GEN647;
wire  _GEN650 = io_x[26] ? _GEN649 : _GEN646;
wire  _GEN651 = io_x[3] ? _GEN650 : _GEN643;
wire  _GEN652 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN653 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN654 = io_x[24] ? _GEN653 : _GEN652;
wire  _GEN655 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN656 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN657 = io_x[24] ? _GEN656 : _GEN655;
wire  _GEN658 = io_x[26] ? _GEN657 : _GEN654;
wire  _GEN659 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN660 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN661 = io_x[24] ? _GEN660 : _GEN659;
wire  _GEN662 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN663 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN664 = io_x[24] ? _GEN663 : _GEN662;
wire  _GEN665 = io_x[26] ? _GEN664 : _GEN661;
wire  _GEN666 = io_x[3] ? _GEN665 : _GEN658;
wire  _GEN667 = io_x[8] ? _GEN666 : _GEN651;
wire  _GEN668 = io_x[4] ? _GEN667 : _GEN636;
wire  _GEN669 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN670 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN671 = io_x[24] ? _GEN670 : _GEN669;
wire  _GEN672 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN673 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN674 = io_x[24] ? _GEN673 : _GEN672;
wire  _GEN675 = io_x[26] ? _GEN674 : _GEN671;
wire  _GEN676 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN677 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN678 = io_x[24] ? _GEN677 : _GEN676;
wire  _GEN679 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN680 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN681 = io_x[24] ? _GEN680 : _GEN679;
wire  _GEN682 = io_x[26] ? _GEN681 : _GEN678;
wire  _GEN683 = io_x[3] ? _GEN682 : _GEN675;
wire  _GEN684 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN685 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN686 = io_x[24] ? _GEN685 : _GEN684;
wire  _GEN687 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN688 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN689 = io_x[24] ? _GEN688 : _GEN687;
wire  _GEN690 = io_x[26] ? _GEN689 : _GEN686;
wire  _GEN691 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN692 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN693 = io_x[24] ? _GEN692 : _GEN691;
wire  _GEN694 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN695 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN696 = io_x[24] ? _GEN695 : _GEN694;
wire  _GEN697 = io_x[26] ? _GEN696 : _GEN693;
wire  _GEN698 = io_x[3] ? _GEN697 : _GEN690;
wire  _GEN699 = io_x[8] ? _GEN698 : _GEN683;
wire  _GEN700 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN701 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN702 = io_x[24] ? _GEN701 : _GEN700;
wire  _GEN703 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN704 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN705 = io_x[24] ? _GEN704 : _GEN703;
wire  _GEN706 = io_x[26] ? _GEN705 : _GEN702;
wire  _GEN707 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN708 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN709 = io_x[24] ? _GEN708 : _GEN707;
wire  _GEN710 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN711 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN712 = io_x[24] ? _GEN711 : _GEN710;
wire  _GEN713 = io_x[26] ? _GEN712 : _GEN709;
wire  _GEN714 = io_x[3] ? _GEN713 : _GEN706;
wire  _GEN715 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN716 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN717 = io_x[24] ? _GEN716 : _GEN715;
wire  _GEN718 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN719 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN720 = io_x[24] ? _GEN719 : _GEN718;
wire  _GEN721 = io_x[26] ? _GEN720 : _GEN717;
wire  _GEN722 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN723 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN724 = io_x[24] ? _GEN723 : _GEN722;
wire  _GEN725 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN726 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN727 = io_x[24] ? _GEN726 : _GEN725;
wire  _GEN728 = io_x[26] ? _GEN727 : _GEN724;
wire  _GEN729 = io_x[3] ? _GEN728 : _GEN721;
wire  _GEN730 = io_x[8] ? _GEN729 : _GEN714;
wire  _GEN731 = io_x[4] ? _GEN730 : _GEN699;
wire  _GEN732 = io_x[12] ? _GEN731 : _GEN668;
wire  _GEN733 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN734 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN735 = io_x[24] ? _GEN734 : _GEN733;
wire  _GEN736 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN737 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN738 = io_x[24] ? _GEN737 : _GEN736;
wire  _GEN739 = io_x[26] ? _GEN738 : _GEN735;
wire  _GEN740 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN741 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN742 = io_x[24] ? _GEN741 : _GEN740;
wire  _GEN743 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN744 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN745 = io_x[24] ? _GEN744 : _GEN743;
wire  _GEN746 = io_x[26] ? _GEN745 : _GEN742;
wire  _GEN747 = io_x[3] ? _GEN746 : _GEN739;
wire  _GEN748 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN749 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN750 = io_x[24] ? _GEN749 : _GEN748;
wire  _GEN751 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN752 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN753 = io_x[24] ? _GEN752 : _GEN751;
wire  _GEN754 = io_x[26] ? _GEN753 : _GEN750;
wire  _GEN755 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN756 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN757 = io_x[24] ? _GEN756 : _GEN755;
wire  _GEN758 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN759 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN760 = io_x[24] ? _GEN759 : _GEN758;
wire  _GEN761 = io_x[26] ? _GEN760 : _GEN757;
wire  _GEN762 = io_x[3] ? _GEN761 : _GEN754;
wire  _GEN763 = io_x[8] ? _GEN762 : _GEN747;
wire  _GEN764 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN765 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN766 = io_x[24] ? _GEN765 : _GEN764;
wire  _GEN767 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN768 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN769 = io_x[24] ? _GEN768 : _GEN767;
wire  _GEN770 = io_x[26] ? _GEN769 : _GEN766;
wire  _GEN771 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN772 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN773 = io_x[24] ? _GEN772 : _GEN771;
wire  _GEN774 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN775 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN776 = io_x[24] ? _GEN775 : _GEN774;
wire  _GEN777 = io_x[26] ? _GEN776 : _GEN773;
wire  _GEN778 = io_x[3] ? _GEN777 : _GEN770;
wire  _GEN779 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN780 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN781 = io_x[24] ? _GEN780 : _GEN779;
wire  _GEN782 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN783 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN784 = io_x[24] ? _GEN783 : _GEN782;
wire  _GEN785 = io_x[26] ? _GEN784 : _GEN781;
wire  _GEN786 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN787 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN788 = io_x[24] ? _GEN787 : _GEN786;
wire  _GEN789 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN790 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN791 = io_x[24] ? _GEN790 : _GEN789;
wire  _GEN792 = io_x[26] ? _GEN791 : _GEN788;
wire  _GEN793 = io_x[3] ? _GEN792 : _GEN785;
wire  _GEN794 = io_x[8] ? _GEN793 : _GEN778;
wire  _GEN795 = io_x[4] ? _GEN794 : _GEN763;
wire  _GEN796 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN797 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN798 = io_x[24] ? _GEN797 : _GEN796;
wire  _GEN799 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN800 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN801 = io_x[24] ? _GEN800 : _GEN799;
wire  _GEN802 = io_x[26] ? _GEN801 : _GEN798;
wire  _GEN803 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN804 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN805 = io_x[24] ? _GEN804 : _GEN803;
wire  _GEN806 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN807 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN808 = io_x[24] ? _GEN807 : _GEN806;
wire  _GEN809 = io_x[26] ? _GEN808 : _GEN805;
wire  _GEN810 = io_x[3] ? _GEN809 : _GEN802;
wire  _GEN811 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN812 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN813 = io_x[24] ? _GEN812 : _GEN811;
wire  _GEN814 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN815 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN816 = io_x[24] ? _GEN815 : _GEN814;
wire  _GEN817 = io_x[26] ? _GEN816 : _GEN813;
wire  _GEN818 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN819 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN820 = io_x[24] ? _GEN819 : _GEN818;
wire  _GEN821 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN822 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN823 = io_x[24] ? _GEN822 : _GEN821;
wire  _GEN824 = io_x[26] ? _GEN823 : _GEN820;
wire  _GEN825 = io_x[3] ? _GEN824 : _GEN817;
wire  _GEN826 = io_x[8] ? _GEN825 : _GEN810;
wire  _GEN827 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN828 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN829 = io_x[24] ? _GEN828 : _GEN827;
wire  _GEN830 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN831 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN832 = io_x[24] ? _GEN831 : _GEN830;
wire  _GEN833 = io_x[26] ? _GEN832 : _GEN829;
wire  _GEN834 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN835 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN836 = io_x[24] ? _GEN835 : _GEN834;
wire  _GEN837 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN838 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN839 = io_x[24] ? _GEN838 : _GEN837;
wire  _GEN840 = io_x[26] ? _GEN839 : _GEN836;
wire  _GEN841 = io_x[3] ? _GEN840 : _GEN833;
wire  _GEN842 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN843 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN844 = io_x[24] ? _GEN843 : _GEN842;
wire  _GEN845 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN846 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN847 = io_x[24] ? _GEN846 : _GEN845;
wire  _GEN848 = io_x[26] ? _GEN847 : _GEN844;
wire  _GEN849 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN850 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN851 = io_x[24] ? _GEN850 : _GEN849;
wire  _GEN852 = io_x[0] ? _GEN604 : _GEN605;
wire  _GEN853 = io_x[0] ? _GEN605 : _GEN604;
wire  _GEN854 = io_x[24] ? _GEN853 : _GEN852;
wire  _GEN855 = io_x[26] ? _GEN854 : _GEN851;
wire  _GEN856 = io_x[3] ? _GEN855 : _GEN848;
wire  _GEN857 = io_x[8] ? _GEN856 : _GEN841;
wire  _GEN858 = io_x[4] ? _GEN857 : _GEN826;
wire  _GEN859 = io_x[12] ? _GEN858 : _GEN795;
wire  _GEN860 = io_x[16] ? _GEN859 : _GEN732;
assign io_y[6] = _GEN860;
wire  _GEN861 = 1'b0;
wire  _GEN862 = 1'b1;
wire  _GEN863 = io_x[23] ? _GEN862 : _GEN861;
wire  _GEN864 = io_x[23] ? _GEN862 : _GEN861;
wire  _GEN865 = io_x[24] ? _GEN864 : _GEN863;
wire  _GEN866 = io_x[23] ? _GEN862 : _GEN861;
wire  _GEN867 = io_x[23] ? _GEN862 : _GEN861;
wire  _GEN868 = io_x[24] ? _GEN867 : _GEN866;
wire  _GEN869 = io_x[15] ? _GEN868 : _GEN865;
assign io_y[5] = _GEN869;
wire  _GEN870 = 1'b0;
wire  _GEN871 = 1'b1;
wire  _GEN872 = io_x[22] ? _GEN871 : _GEN870;
wire  _GEN873 = io_x[22] ? _GEN871 : _GEN870;
wire  _GEN874 = io_x[19] ? _GEN873 : _GEN872;
wire  _GEN875 = io_x[22] ? _GEN871 : _GEN870;
wire  _GEN876 = io_x[22] ? _GEN871 : _GEN870;
wire  _GEN877 = io_x[19] ? _GEN876 : _GEN875;
wire  _GEN878 = io_x[28] ? _GEN877 : _GEN874;
wire  _GEN879 = io_x[22] ? _GEN871 : _GEN870;
wire  _GEN880 = io_x[22] ? _GEN871 : _GEN870;
wire  _GEN881 = io_x[19] ? _GEN880 : _GEN879;
wire  _GEN882 = io_x[22] ? _GEN871 : _GEN870;
wire  _GEN883 = io_x[22] ? _GEN871 : _GEN870;
wire  _GEN884 = io_x[19] ? _GEN883 : _GEN882;
wire  _GEN885 = io_x[28] ? _GEN884 : _GEN881;
wire  _GEN886 = io_x[21] ? _GEN885 : _GEN878;
assign io_y[4] = _GEN886;
wire  _GEN887 = 1'b0;
wire  _GEN888 = 1'b1;
wire  _GEN889 = io_x[21] ? _GEN888 : _GEN887;
assign io_y[3] = _GEN889;
wire  _GEN890 = 1'b0;
wire  _GEN891 = 1'b1;
wire  _GEN892 = io_x[20] ? _GEN891 : _GEN890;
wire  _GEN893 = io_x[20] ? _GEN891 : _GEN890;
wire  _GEN894 = io_x[1] ? _GEN893 : _GEN892;
wire  _GEN895 = io_x[20] ? _GEN891 : _GEN890;
wire  _GEN896 = io_x[20] ? _GEN891 : _GEN890;
wire  _GEN897 = io_x[1] ? _GEN896 : _GEN895;
wire  _GEN898 = io_x[25] ? _GEN897 : _GEN894;
wire  _GEN899 = io_x[20] ? _GEN891 : _GEN890;
wire  _GEN900 = io_x[20] ? _GEN891 : _GEN890;
wire  _GEN901 = io_x[1] ? _GEN900 : _GEN899;
wire  _GEN902 = io_x[20] ? _GEN891 : _GEN890;
wire  _GEN903 = io_x[20] ? _GEN891 : _GEN890;
wire  _GEN904 = io_x[1] ? _GEN903 : _GEN902;
wire  _GEN905 = io_x[25] ? _GEN904 : _GEN901;
wire  _GEN906 = io_x[27] ? _GEN905 : _GEN898;
assign io_y[2] = _GEN906;
wire  _GEN907 = 1'b0;
wire  _GEN908 = 1'b1;
wire  _GEN909 = io_x[19] ? _GEN908 : _GEN907;
wire  _GEN910 = io_x[19] ? _GEN908 : _GEN907;
wire  _GEN911 = io_x[23] ? _GEN910 : _GEN909;
assign io_y[1] = _GEN911;
wire  _GEN912 = 1'b0;
wire  _GEN913 = 1'b1;
wire  _GEN914 = io_x[16] ? _GEN913 : _GEN912;
wire  _GEN915 = io_x[16] ? _GEN913 : _GEN912;
wire  _GEN916 = io_x[26] ? _GEN915 : _GEN914;
assign io_y[0] = _GEN916;
endmodule
