module BBGSharePredictorImp_BSD_b_NutShell_less(
    input [31:0] pc,
    input [31:0] train_pc,
    input  train_taken,
    input [1:0] pht_rdata,
    input [15:0] ghr_rdata,
    input [15:0] train_ghr_rdata,
    output  taken,
    output  pht_wdata,
    output [8:0] pht_raddr,
    output [8:0] pht_waddr,
    output  ghr_wdata
);
wire [98:0] io_x;
wire [20:0] io_y;
assign io_x = { pc, train_pc, train_taken, pht_rdata, ghr_rdata, train_ghr_rdata };
assign { taken, pht_wdata, pht_raddr, pht_waddr, ghr_wdata } = io_y;
wire  _GEN0 = 1'b0;
wire  _GEN1 = 1'b1;
wire  _GEN2 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN3 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN4 = io_x[32] ? _GEN3 : _GEN2;
wire  _GEN5 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN6 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN7 = io_x[32] ? _GEN6 : _GEN5;
wire  _GEN8 = io_x[20] ? _GEN7 : _GEN4;
wire  _GEN9 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN10 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN11 = io_x[32] ? _GEN10 : _GEN9;
wire  _GEN12 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN13 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN14 = io_x[32] ? _GEN13 : _GEN12;
wire  _GEN15 = io_x[20] ? _GEN14 : _GEN11;
wire  _GEN16 = io_x[49] ? _GEN15 : _GEN8;
wire  _GEN17 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN18 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN19 = io_x[32] ? _GEN18 : _GEN17;
wire  _GEN20 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN21 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN22 = io_x[32] ? _GEN21 : _GEN20;
wire  _GEN23 = io_x[20] ? _GEN22 : _GEN19;
wire  _GEN24 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN25 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN26 = io_x[32] ? _GEN25 : _GEN24;
wire  _GEN27 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN28 = io_x[33] ? _GEN1 : _GEN0;
wire  _GEN29 = io_x[32] ? _GEN28 : _GEN27;
wire  _GEN30 = io_x[20] ? _GEN29 : _GEN26;
wire  _GEN31 = io_x[49] ? _GEN30 : _GEN23;
wire  _GEN32 = io_x[80] ? _GEN31 : _GEN16;
assign io_y[20] = _GEN32;
wire  _GEN33 = 1'b0;
wire  _GEN34 = 1'b1;
wire  _GEN35 = io_x[34] ? _GEN34 : _GEN33;
wire  _GEN36 = io_x[34] ? _GEN34 : _GEN33;
wire  _GEN37 = io_x[45] ? _GEN36 : _GEN35;
assign io_y[19] = _GEN37;
wire  _GEN38 = 1'b0;
wire  _GEN39 = 1'b1;
wire  _GEN40 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN41 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN42 = io_x[27] ? _GEN41 : _GEN40;
wire  _GEN43 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN44 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN45 = io_x[27] ? _GEN44 : _GEN43;
wire  _GEN46 = io_x[31] ? _GEN45 : _GEN42;
wire  _GEN47 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN48 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN49 = io_x[27] ? _GEN48 : _GEN47;
wire  _GEN50 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN51 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN52 = io_x[27] ? _GEN51 : _GEN50;
wire  _GEN53 = io_x[31] ? _GEN52 : _GEN49;
wire  _GEN54 = io_x[23] ? _GEN53 : _GEN46;
wire  _GEN55 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN56 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN57 = io_x[27] ? _GEN56 : _GEN55;
wire  _GEN58 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN59 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN60 = io_x[27] ? _GEN59 : _GEN58;
wire  _GEN61 = io_x[31] ? _GEN60 : _GEN57;
wire  _GEN62 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN63 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN64 = io_x[27] ? _GEN63 : _GEN62;
wire  _GEN65 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN66 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN67 = io_x[27] ? _GEN66 : _GEN65;
wire  _GEN68 = io_x[31] ? _GEN67 : _GEN64;
wire  _GEN69 = io_x[23] ? _GEN68 : _GEN61;
wire  _GEN70 = io_x[77] ? _GEN69 : _GEN54;
wire  _GEN71 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN72 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN73 = io_x[27] ? _GEN72 : _GEN71;
wire  _GEN74 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN75 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN76 = io_x[27] ? _GEN75 : _GEN74;
wire  _GEN77 = io_x[31] ? _GEN76 : _GEN73;
wire  _GEN78 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN79 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN80 = io_x[27] ? _GEN79 : _GEN78;
wire  _GEN81 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN82 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN83 = io_x[27] ? _GEN82 : _GEN81;
wire  _GEN84 = io_x[31] ? _GEN83 : _GEN80;
wire  _GEN85 = io_x[23] ? _GEN84 : _GEN77;
wire  _GEN86 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN87 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN88 = io_x[27] ? _GEN87 : _GEN86;
wire  _GEN89 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN90 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN91 = io_x[27] ? _GEN90 : _GEN89;
wire  _GEN92 = io_x[31] ? _GEN91 : _GEN88;
wire  _GEN93 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN94 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN95 = io_x[27] ? _GEN94 : _GEN93;
wire  _GEN96 = io_x[19] ? _GEN38 : _GEN39;
wire  _GEN97 = io_x[19] ? _GEN39 : _GEN38;
wire  _GEN98 = io_x[27] ? _GEN97 : _GEN96;
wire  _GEN99 = io_x[31] ? _GEN98 : _GEN95;
wire  _GEN100 = io_x[23] ? _GEN99 : _GEN92;
wire  _GEN101 = io_x[77] ? _GEN100 : _GEN85;
wire  _GEN102 = io_x[49] ? _GEN101 : _GEN70;
assign io_y[18] = _GEN102;
wire  _GEN103 = 1'b0;
wire  _GEN104 = 1'b1;
wire  _GEN105 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN106 = 1'b0;
wire  _GEN107 = io_x[30] ? _GEN106 : _GEN105;
wire  _GEN108 = 1'b0;
wire  _GEN109 = io_x[26] ? _GEN108 : _GEN107;
wire  _GEN110 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN111 = io_x[30] ? _GEN106 : _GEN110;
wire  _GEN112 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN113 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN114 = io_x[30] ? _GEN113 : _GEN112;
wire  _GEN115 = io_x[26] ? _GEN114 : _GEN111;
wire  _GEN116 = io_x[22] ? _GEN115 : _GEN109;
wire  _GEN117 = 1'b1;
wire  _GEN118 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN119 = 1'b1;
wire  _GEN120 = io_x[26] ? _GEN119 : _GEN118;
wire  _GEN121 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN122 = io_x[30] ? _GEN121 : _GEN117;
wire  _GEN123 = io_x[26] ? _GEN122 : _GEN119;
wire  _GEN124 = io_x[22] ? _GEN123 : _GEN120;
wire  _GEN125 = io_x[13] ? _GEN124 : _GEN116;
wire  _GEN126 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN127 = io_x[30] ? _GEN106 : _GEN126;
wire  _GEN128 = io_x[26] ? _GEN108 : _GEN127;
wire  _GEN129 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN130 = io_x[30] ? _GEN129 : _GEN106;
wire  _GEN131 = io_x[26] ? _GEN119 : _GEN130;
wire  _GEN132 = io_x[22] ? _GEN131 : _GEN128;
wire  _GEN133 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN134 = io_x[30] ? _GEN133 : _GEN117;
wire  _GEN135 = io_x[26] ? _GEN134 : _GEN108;
wire  _GEN136 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN137 = io_x[30] ? _GEN136 : _GEN106;
wire  _GEN138 = io_x[26] ? _GEN137 : _GEN119;
wire  _GEN139 = io_x[22] ? _GEN138 : _GEN135;
wire  _GEN140 = io_x[13] ? _GEN139 : _GEN132;
wire  _GEN141 = io_x[33] ? _GEN140 : _GEN125;
wire  _GEN142 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN143 = io_x[30] ? _GEN106 : _GEN142;
wire  _GEN144 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN145 = io_x[30] ? _GEN144 : _GEN106;
wire  _GEN146 = io_x[26] ? _GEN145 : _GEN143;
wire  _GEN147 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN148 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN149 = io_x[30] ? _GEN148 : _GEN147;
wire  _GEN150 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN151 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN152 = io_x[30] ? _GEN151 : _GEN150;
wire  _GEN153 = io_x[26] ? _GEN152 : _GEN149;
wire  _GEN154 = io_x[22] ? _GEN153 : _GEN146;
wire  _GEN155 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN156 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN157 = io_x[30] ? _GEN156 : _GEN155;
wire  _GEN158 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN159 = io_x[30] ? _GEN158 : _GEN117;
wire  _GEN160 = io_x[26] ? _GEN159 : _GEN157;
wire  _GEN161 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN162 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN163 = io_x[30] ? _GEN162 : _GEN106;
wire  _GEN164 = io_x[26] ? _GEN163 : _GEN161;
wire  _GEN165 = io_x[22] ? _GEN164 : _GEN160;
wire  _GEN166 = io_x[13] ? _GEN165 : _GEN154;
wire  _GEN167 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN168 = io_x[30] ? _GEN117 : _GEN167;
wire  _GEN169 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN170 = io_x[30] ? _GEN106 : _GEN169;
wire  _GEN171 = io_x[26] ? _GEN170 : _GEN168;
wire  _GEN172 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN173 = io_x[30] ? _GEN106 : _GEN172;
wire  _GEN174 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN175 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN176 = io_x[30] ? _GEN175 : _GEN174;
wire  _GEN177 = io_x[26] ? _GEN176 : _GEN173;
wire  _GEN178 = io_x[22] ? _GEN177 : _GEN171;
wire  _GEN179 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN180 = io_x[30] ? _GEN106 : _GEN179;
wire  _GEN181 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN182 = io_x[30] ? _GEN181 : _GEN106;
wire  _GEN183 = io_x[26] ? _GEN182 : _GEN180;
wire  _GEN184 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN185 = io_x[30] ? _GEN117 : _GEN184;
wire  _GEN186 = io_x[26] ? _GEN185 : _GEN119;
wire  _GEN187 = io_x[22] ? _GEN186 : _GEN183;
wire  _GEN188 = io_x[13] ? _GEN187 : _GEN178;
wire  _GEN189 = io_x[33] ? _GEN188 : _GEN166;
wire  _GEN190 = io_x[69] ? _GEN189 : _GEN141;
wire  _GEN191 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN192 = io_x[30] ? _GEN106 : _GEN191;
wire  _GEN193 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN194 = io_x[30] ? _GEN193 : _GEN106;
wire  _GEN195 = io_x[26] ? _GEN194 : _GEN192;
wire  _GEN196 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN197 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN198 = io_x[30] ? _GEN197 : _GEN196;
wire  _GEN199 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN200 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN201 = io_x[30] ? _GEN200 : _GEN199;
wire  _GEN202 = io_x[26] ? _GEN201 : _GEN198;
wire  _GEN203 = io_x[22] ? _GEN202 : _GEN195;
wire  _GEN204 = 1'b0;
wire  _GEN205 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN206 = io_x[30] ? _GEN205 : _GEN106;
wire  _GEN207 = io_x[26] ? _GEN206 : _GEN108;
wire  _GEN208 = io_x[22] ? _GEN207 : _GEN204;
wire  _GEN209 = io_x[13] ? _GEN208 : _GEN203;
wire  _GEN210 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN211 = io_x[30] ? _GEN106 : _GEN210;
wire  _GEN212 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN213 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN214 = io_x[30] ? _GEN213 : _GEN212;
wire  _GEN215 = io_x[26] ? _GEN214 : _GEN211;
wire  _GEN216 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN217 = io_x[30] ? _GEN216 : _GEN106;
wire  _GEN218 = io_x[26] ? _GEN217 : _GEN108;
wire  _GEN219 = io_x[22] ? _GEN218 : _GEN215;
wire  _GEN220 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN221 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN222 = io_x[30] ? _GEN221 : _GEN117;
wire  _GEN223 = io_x[26] ? _GEN222 : _GEN220;
wire  _GEN224 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN225 = io_x[30] ? _GEN224 : _GEN117;
wire  _GEN226 = io_x[26] ? _GEN225 : _GEN108;
wire  _GEN227 = io_x[22] ? _GEN226 : _GEN223;
wire  _GEN228 = io_x[13] ? _GEN227 : _GEN219;
wire  _GEN229 = io_x[33] ? _GEN228 : _GEN209;
wire  _GEN230 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN231 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN232 = io_x[30] ? _GEN231 : _GEN230;
wire  _GEN233 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN234 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN235 = io_x[30] ? _GEN234 : _GEN233;
wire  _GEN236 = io_x[26] ? _GEN235 : _GEN232;
wire  _GEN237 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN238 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN239 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN240 = io_x[30] ? _GEN239 : _GEN238;
wire  _GEN241 = io_x[26] ? _GEN240 : _GEN237;
wire  _GEN242 = io_x[22] ? _GEN241 : _GEN236;
wire  _GEN243 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN244 = io_x[26] ? _GEN119 : _GEN243;
wire  _GEN245 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN246 = io_x[26] ? _GEN245 : _GEN108;
wire  _GEN247 = io_x[22] ? _GEN246 : _GEN244;
wire  _GEN248 = io_x[13] ? _GEN247 : _GEN242;
wire  _GEN249 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN250 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN251 = io_x[30] ? _GEN250 : _GEN249;
wire  _GEN252 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN253 = io_x[26] ? _GEN252 : _GEN251;
wire  _GEN254 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN255 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN256 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN257 = io_x[30] ? _GEN256 : _GEN255;
wire  _GEN258 = io_x[26] ? _GEN257 : _GEN254;
wire  _GEN259 = io_x[22] ? _GEN258 : _GEN253;
wire  _GEN260 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN261 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN262 = io_x[30] ? _GEN261 : _GEN117;
wire  _GEN263 = io_x[26] ? _GEN262 : _GEN260;
wire  _GEN264 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN265 = io_x[30] ? _GEN264 : _GEN117;
wire  _GEN266 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN267 = io_x[30] ? _GEN266 : _GEN117;
wire  _GEN268 = io_x[26] ? _GEN267 : _GEN265;
wire  _GEN269 = io_x[22] ? _GEN268 : _GEN263;
wire  _GEN270 = io_x[13] ? _GEN269 : _GEN259;
wire  _GEN271 = io_x[33] ? _GEN270 : _GEN248;
wire  _GEN272 = io_x[69] ? _GEN271 : _GEN229;
wire  _GEN273 = io_x[71] ? _GEN272 : _GEN190;
wire  _GEN274 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN275 = io_x[30] ? _GEN106 : _GEN274;
wire  _GEN276 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN277 = io_x[30] ? _GEN276 : _GEN106;
wire  _GEN278 = io_x[26] ? _GEN277 : _GEN275;
wire  _GEN279 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN280 = io_x[30] ? _GEN117 : _GEN279;
wire  _GEN281 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN282 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN283 = io_x[30] ? _GEN282 : _GEN281;
wire  _GEN284 = io_x[26] ? _GEN283 : _GEN280;
wire  _GEN285 = io_x[22] ? _GEN284 : _GEN278;
wire  _GEN286 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN287 = io_x[30] ? _GEN286 : _GEN117;
wire  _GEN288 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN289 = io_x[26] ? _GEN288 : _GEN287;
wire  _GEN290 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN291 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN292 = io_x[30] ? _GEN117 : _GEN291;
wire  _GEN293 = io_x[26] ? _GEN292 : _GEN290;
wire  _GEN294 = io_x[22] ? _GEN293 : _GEN289;
wire  _GEN295 = io_x[13] ? _GEN294 : _GEN285;
wire  _GEN296 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN297 = io_x[30] ? _GEN106 : _GEN296;
wire  _GEN298 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN299 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN300 = io_x[30] ? _GEN299 : _GEN298;
wire  _GEN301 = io_x[26] ? _GEN300 : _GEN297;
wire  _GEN302 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN303 = io_x[30] ? _GEN117 : _GEN302;
wire  _GEN304 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN305 = io_x[30] ? _GEN106 : _GEN304;
wire  _GEN306 = io_x[26] ? _GEN305 : _GEN303;
wire  _GEN307 = io_x[22] ? _GEN306 : _GEN301;
wire  _GEN308 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN309 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN310 = io_x[30] ? _GEN309 : _GEN308;
wire  _GEN311 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN312 = io_x[30] ? _GEN311 : _GEN117;
wire  _GEN313 = io_x[26] ? _GEN312 : _GEN310;
wire  _GEN314 = 1'b1;
wire  _GEN315 = io_x[22] ? _GEN314 : _GEN313;
wire  _GEN316 = io_x[13] ? _GEN315 : _GEN307;
wire  _GEN317 = io_x[33] ? _GEN316 : _GEN295;
wire  _GEN318 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN319 = io_x[30] ? _GEN106 : _GEN318;
wire  _GEN320 = io_x[26] ? _GEN119 : _GEN319;
wire  _GEN321 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN322 = io_x[30] ? _GEN321 : _GEN117;
wire  _GEN323 = io_x[26] ? _GEN108 : _GEN322;
wire  _GEN324 = io_x[22] ? _GEN323 : _GEN320;
wire  _GEN325 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN326 = io_x[26] ? _GEN325 : _GEN108;
wire  _GEN327 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN328 = io_x[30] ? _GEN327 : _GEN117;
wire  _GEN329 = io_x[26] ? _GEN328 : _GEN119;
wire  _GEN330 = io_x[22] ? _GEN329 : _GEN326;
wire  _GEN331 = io_x[13] ? _GEN330 : _GEN324;
wire  _GEN332 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN333 = io_x[30] ? _GEN332 : _GEN117;
wire  _GEN334 = io_x[26] ? _GEN333 : _GEN108;
wire  _GEN335 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN336 = io_x[30] ? _GEN117 : _GEN335;
wire  _GEN337 = io_x[26] ? _GEN108 : _GEN336;
wire  _GEN338 = io_x[22] ? _GEN337 : _GEN334;
wire  _GEN339 = io_x[26] ? _GEN108 : _GEN119;
wire  _GEN340 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN341 = io_x[30] ? _GEN340 : _GEN117;
wire  _GEN342 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN343 = io_x[30] ? _GEN342 : _GEN117;
wire  _GEN344 = io_x[26] ? _GEN343 : _GEN341;
wire  _GEN345 = io_x[22] ? _GEN344 : _GEN339;
wire  _GEN346 = io_x[13] ? _GEN345 : _GEN338;
wire  _GEN347 = io_x[33] ? _GEN346 : _GEN331;
wire  _GEN348 = io_x[69] ? _GEN347 : _GEN317;
wire  _GEN349 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN350 = io_x[30] ? _GEN117 : _GEN349;
wire  _GEN351 = io_x[26] ? _GEN108 : _GEN350;
wire  _GEN352 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN353 = io_x[30] ? _GEN106 : _GEN352;
wire  _GEN354 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN355 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN356 = io_x[30] ? _GEN355 : _GEN354;
wire  _GEN357 = io_x[26] ? _GEN356 : _GEN353;
wire  _GEN358 = io_x[22] ? _GEN357 : _GEN351;
wire  _GEN359 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN360 = io_x[30] ? _GEN359 : _GEN117;
wire  _GEN361 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN362 = io_x[30] ? _GEN361 : _GEN117;
wire  _GEN363 = io_x[26] ? _GEN362 : _GEN360;
wire  _GEN364 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN365 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN366 = io_x[30] ? _GEN365 : _GEN117;
wire  _GEN367 = io_x[26] ? _GEN366 : _GEN364;
wire  _GEN368 = io_x[22] ? _GEN367 : _GEN363;
wire  _GEN369 = io_x[13] ? _GEN368 : _GEN358;
wire  _GEN370 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN371 = io_x[30] ? _GEN117 : _GEN370;
wire  _GEN372 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN373 = io_x[30] ? _GEN117 : _GEN372;
wire  _GEN374 = io_x[26] ? _GEN373 : _GEN371;
wire  _GEN375 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN376 = io_x[30] ? _GEN106 : _GEN375;
wire  _GEN377 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN378 = io_x[26] ? _GEN377 : _GEN376;
wire  _GEN379 = io_x[22] ? _GEN378 : _GEN374;
wire  _GEN380 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN381 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN382 = io_x[30] ? _GEN381 : _GEN380;
wire  _GEN383 = io_x[26] ? _GEN108 : _GEN382;
wire  _GEN384 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN385 = io_x[30] ? _GEN384 : _GEN117;
wire  _GEN386 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN387 = io_x[30] ? _GEN386 : _GEN117;
wire  _GEN388 = io_x[26] ? _GEN387 : _GEN385;
wire  _GEN389 = io_x[22] ? _GEN388 : _GEN383;
wire  _GEN390 = io_x[13] ? _GEN389 : _GEN379;
wire  _GEN391 = io_x[33] ? _GEN390 : _GEN369;
wire  _GEN392 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN393 = io_x[30] ? _GEN106 : _GEN392;
wire  _GEN394 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN395 = io_x[26] ? _GEN394 : _GEN393;
wire  _GEN396 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN397 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN398 = io_x[30] ? _GEN397 : _GEN117;
wire  _GEN399 = io_x[26] ? _GEN398 : _GEN396;
wire  _GEN400 = io_x[22] ? _GEN399 : _GEN395;
wire  _GEN401 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN402 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN403 = io_x[26] ? _GEN402 : _GEN401;
wire  _GEN404 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN405 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN406 = io_x[30] ? _GEN405 : _GEN404;
wire  _GEN407 = io_x[26] ? _GEN119 : _GEN406;
wire  _GEN408 = io_x[22] ? _GEN407 : _GEN403;
wire  _GEN409 = io_x[13] ? _GEN408 : _GEN400;
wire  _GEN410 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN411 = io_x[30] ? _GEN106 : _GEN410;
wire  _GEN412 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN413 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN414 = io_x[30] ? _GEN413 : _GEN412;
wire  _GEN415 = io_x[26] ? _GEN414 : _GEN411;
wire  _GEN416 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN417 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN418 = io_x[30] ? _GEN417 : _GEN416;
wire  _GEN419 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN420 = io_x[30] ? _GEN106 : _GEN419;
wire  _GEN421 = io_x[26] ? _GEN420 : _GEN418;
wire  _GEN422 = io_x[22] ? _GEN421 : _GEN415;
wire  _GEN423 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN424 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN425 = io_x[30] ? _GEN106 : _GEN424;
wire  _GEN426 = io_x[26] ? _GEN425 : _GEN423;
wire  _GEN427 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN428 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN429 = io_x[30] ? _GEN428 : _GEN117;
wire  _GEN430 = io_x[26] ? _GEN429 : _GEN427;
wire  _GEN431 = io_x[22] ? _GEN430 : _GEN426;
wire  _GEN432 = io_x[13] ? _GEN431 : _GEN422;
wire  _GEN433 = io_x[33] ? _GEN432 : _GEN409;
wire  _GEN434 = io_x[69] ? _GEN433 : _GEN391;
wire  _GEN435 = io_x[71] ? _GEN434 : _GEN348;
wire  _GEN436 = io_x[72] ? _GEN435 : _GEN273;
wire  _GEN437 = io_x[26] ? _GEN108 : _GEN119;
wire  _GEN438 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN439 = io_x[30] ? _GEN117 : _GEN438;
wire  _GEN440 = io_x[26] ? _GEN119 : _GEN439;
wire  _GEN441 = io_x[22] ? _GEN440 : _GEN437;
wire  _GEN442 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN443 = io_x[22] ? _GEN204 : _GEN442;
wire  _GEN444 = io_x[13] ? _GEN443 : _GEN441;
wire  _GEN445 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN446 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN447 = io_x[26] ? _GEN446 : _GEN445;
wire  _GEN448 = io_x[22] ? _GEN204 : _GEN447;
wire  _GEN449 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN450 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN451 = io_x[26] ? _GEN108 : _GEN450;
wire  _GEN452 = io_x[22] ? _GEN451 : _GEN449;
wire  _GEN453 = io_x[13] ? _GEN452 : _GEN448;
wire  _GEN454 = io_x[33] ? _GEN453 : _GEN444;
wire  _GEN455 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN456 = io_x[30] ? _GEN106 : _GEN455;
wire  _GEN457 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN458 = io_x[26] ? _GEN457 : _GEN456;
wire  _GEN459 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN460 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN461 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN462 = io_x[30] ? _GEN461 : _GEN460;
wire  _GEN463 = io_x[26] ? _GEN462 : _GEN459;
wire  _GEN464 = io_x[22] ? _GEN463 : _GEN458;
wire  _GEN465 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN466 = io_x[30] ? _GEN465 : _GEN117;
wire  _GEN467 = io_x[26] ? _GEN466 : _GEN119;
wire  _GEN468 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN469 = io_x[26] ? _GEN468 : _GEN119;
wire  _GEN470 = io_x[22] ? _GEN469 : _GEN467;
wire  _GEN471 = io_x[13] ? _GEN470 : _GEN464;
wire  _GEN472 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN473 = io_x[30] ? _GEN472 : _GEN117;
wire  _GEN474 = io_x[26] ? _GEN473 : _GEN108;
wire  _GEN475 = io_x[22] ? _GEN474 : _GEN204;
wire  _GEN476 = io_x[22] ? _GEN314 : _GEN204;
wire  _GEN477 = io_x[13] ? _GEN476 : _GEN475;
wire  _GEN478 = io_x[33] ? _GEN477 : _GEN471;
wire  _GEN479 = io_x[69] ? _GEN478 : _GEN454;
wire  _GEN480 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN481 = io_x[30] ? _GEN106 : _GEN480;
wire  _GEN482 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN483 = io_x[26] ? _GEN482 : _GEN481;
wire  _GEN484 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN485 = io_x[30] ? _GEN117 : _GEN484;
wire  _GEN486 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN487 = io_x[30] ? _GEN486 : _GEN117;
wire  _GEN488 = io_x[26] ? _GEN487 : _GEN485;
wire  _GEN489 = io_x[22] ? _GEN488 : _GEN483;
wire  _GEN490 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN491 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN492 = io_x[30] ? _GEN491 : _GEN117;
wire  _GEN493 = io_x[26] ? _GEN492 : _GEN108;
wire  _GEN494 = io_x[22] ? _GEN493 : _GEN490;
wire  _GEN495 = io_x[13] ? _GEN494 : _GEN489;
wire  _GEN496 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN497 = io_x[30] ? _GEN117 : _GEN496;
wire  _GEN498 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN499 = io_x[30] ? _GEN117 : _GEN498;
wire  _GEN500 = io_x[26] ? _GEN499 : _GEN497;
wire  _GEN501 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN502 = io_x[30] ? _GEN117 : _GEN501;
wire  _GEN503 = io_x[26] ? _GEN108 : _GEN502;
wire  _GEN504 = io_x[22] ? _GEN503 : _GEN500;
wire  _GEN505 = io_x[22] ? _GEN314 : _GEN204;
wire  _GEN506 = io_x[13] ? _GEN505 : _GEN504;
wire  _GEN507 = io_x[33] ? _GEN506 : _GEN495;
wire  _GEN508 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN509 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN510 = io_x[26] ? _GEN509 : _GEN508;
wire  _GEN511 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN512 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN513 = io_x[26] ? _GEN512 : _GEN511;
wire  _GEN514 = io_x[22] ? _GEN513 : _GEN510;
wire  _GEN515 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN516 = io_x[30] ? _GEN515 : _GEN117;
wire  _GEN517 = io_x[26] ? _GEN516 : _GEN119;
wire  _GEN518 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN519 = io_x[30] ? _GEN518 : _GEN117;
wire  _GEN520 = io_x[26] ? _GEN119 : _GEN519;
wire  _GEN521 = io_x[22] ? _GEN520 : _GEN517;
wire  _GEN522 = io_x[13] ? _GEN521 : _GEN514;
wire  _GEN523 = 1'b0;
wire  _GEN524 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN525 = io_x[22] ? _GEN524 : _GEN314;
wire  _GEN526 = io_x[13] ? _GEN525 : _GEN523;
wire  _GEN527 = io_x[33] ? _GEN526 : _GEN522;
wire  _GEN528 = io_x[69] ? _GEN527 : _GEN507;
wire  _GEN529 = io_x[71] ? _GEN528 : _GEN479;
wire  _GEN530 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN531 = io_x[30] ? _GEN117 : _GEN530;
wire  _GEN532 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN533 = io_x[26] ? _GEN532 : _GEN531;
wire  _GEN534 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN535 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN536 = io_x[30] ? _GEN535 : _GEN117;
wire  _GEN537 = io_x[26] ? _GEN536 : _GEN534;
wire  _GEN538 = io_x[22] ? _GEN537 : _GEN533;
wire  _GEN539 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN540 = io_x[30] ? _GEN539 : _GEN117;
wire  _GEN541 = io_x[26] ? _GEN108 : _GEN540;
wire  _GEN542 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN543 = io_x[26] ? _GEN542 : _GEN108;
wire  _GEN544 = io_x[22] ? _GEN543 : _GEN541;
wire  _GEN545 = io_x[13] ? _GEN544 : _GEN538;
wire  _GEN546 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN547 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN548 = io_x[26] ? _GEN547 : _GEN546;
wire  _GEN549 = io_x[22] ? _GEN204 : _GEN548;
wire  _GEN550 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN551 = io_x[26] ? _GEN550 : _GEN119;
wire  _GEN552 = io_x[22] ? _GEN314 : _GEN551;
wire  _GEN553 = io_x[13] ? _GEN552 : _GEN549;
wire  _GEN554 = io_x[33] ? _GEN553 : _GEN545;
wire  _GEN555 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN556 = io_x[26] ? _GEN555 : _GEN108;
wire  _GEN557 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN558 = io_x[30] ? _GEN106 : _GEN557;
wire  _GEN559 = io_x[26] ? _GEN119 : _GEN558;
wire  _GEN560 = io_x[22] ? _GEN559 : _GEN556;
wire  _GEN561 = io_x[22] ? _GEN204 : _GEN314;
wire  _GEN562 = io_x[13] ? _GEN561 : _GEN560;
wire  _GEN563 = 1'b1;
wire  _GEN564 = io_x[13] ? _GEN563 : _GEN523;
wire  _GEN565 = io_x[33] ? _GEN564 : _GEN562;
wire  _GEN566 = io_x[69] ? _GEN565 : _GEN554;
wire  _GEN567 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN568 = io_x[26] ? _GEN567 : _GEN119;
wire  _GEN569 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN570 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN571 = io_x[30] ? _GEN117 : _GEN570;
wire  _GEN572 = io_x[26] ? _GEN571 : _GEN569;
wire  _GEN573 = io_x[22] ? _GEN572 : _GEN568;
wire  _GEN574 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN575 = io_x[26] ? _GEN108 : _GEN574;
wire  _GEN576 = io_x[22] ? _GEN204 : _GEN575;
wire  _GEN577 = io_x[13] ? _GEN576 : _GEN573;
wire  _GEN578 = io_x[26] ? _GEN108 : _GEN119;
wire  _GEN579 = io_x[22] ? _GEN578 : _GEN204;
wire  _GEN580 = io_x[13] ? _GEN563 : _GEN579;
wire  _GEN581 = io_x[33] ? _GEN580 : _GEN577;
wire  _GEN582 = io_x[13] ? _GEN523 : _GEN563;
wire  _GEN583 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN584 = io_x[30] ? _GEN583 : _GEN117;
wire  _GEN585 = io_x[26] ? _GEN584 : _GEN119;
wire  _GEN586 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN587 = io_x[30] ? _GEN117 : _GEN586;
wire  _GEN588 = io_x[26] ? _GEN587 : _GEN108;
wire  _GEN589 = io_x[22] ? _GEN588 : _GEN585;
wire  _GEN590 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN591 = io_x[30] ? _GEN590 : _GEN117;
wire  _GEN592 = io_x[26] ? _GEN591 : _GEN108;
wire  _GEN593 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN594 = io_x[30] ? _GEN117 : _GEN593;
wire  _GEN595 = io_x[26] ? _GEN119 : _GEN594;
wire  _GEN596 = io_x[22] ? _GEN595 : _GEN592;
wire  _GEN597 = io_x[13] ? _GEN596 : _GEN589;
wire  _GEN598 = io_x[33] ? _GEN597 : _GEN582;
wire  _GEN599 = io_x[69] ? _GEN598 : _GEN581;
wire  _GEN600 = io_x[71] ? _GEN599 : _GEN566;
wire  _GEN601 = io_x[72] ? _GEN600 : _GEN529;
wire  _GEN602 = io_x[48] ? _GEN601 : _GEN436;
wire  _GEN603 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN604 = io_x[30] ? _GEN106 : _GEN603;
wire  _GEN605 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN606 = io_x[30] ? _GEN117 : _GEN605;
wire  _GEN607 = io_x[26] ? _GEN606 : _GEN604;
wire  _GEN608 = io_x[22] ? _GEN314 : _GEN607;
wire  _GEN609 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN610 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN611 = io_x[30] ? _GEN610 : _GEN609;
wire  _GEN612 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN613 = io_x[26] ? _GEN612 : _GEN611;
wire  _GEN614 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN615 = io_x[30] ? _GEN614 : _GEN117;
wire  _GEN616 = io_x[26] ? _GEN615 : _GEN108;
wire  _GEN617 = io_x[22] ? _GEN616 : _GEN613;
wire  _GEN618 = io_x[13] ? _GEN617 : _GEN608;
wire  _GEN619 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN620 = io_x[30] ? _GEN106 : _GEN619;
wire  _GEN621 = io_x[26] ? _GEN108 : _GEN620;
wire  _GEN622 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN623 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN624 = io_x[30] ? _GEN623 : _GEN622;
wire  _GEN625 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN626 = io_x[30] ? _GEN625 : _GEN106;
wire  _GEN627 = io_x[26] ? _GEN626 : _GEN624;
wire  _GEN628 = io_x[22] ? _GEN627 : _GEN621;
wire  _GEN629 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN630 = io_x[26] ? _GEN119 : _GEN629;
wire  _GEN631 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN632 = io_x[30] ? _GEN631 : _GEN106;
wire  _GEN633 = io_x[26] ? _GEN632 : _GEN108;
wire  _GEN634 = io_x[22] ? _GEN633 : _GEN630;
wire  _GEN635 = io_x[13] ? _GEN634 : _GEN628;
wire  _GEN636 = io_x[33] ? _GEN635 : _GEN618;
wire  _GEN637 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN638 = io_x[30] ? _GEN117 : _GEN637;
wire  _GEN639 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN640 = io_x[30] ? _GEN117 : _GEN639;
wire  _GEN641 = io_x[26] ? _GEN640 : _GEN638;
wire  _GEN642 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN643 = io_x[30] ? _GEN117 : _GEN642;
wire  _GEN644 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN645 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN646 = io_x[30] ? _GEN645 : _GEN644;
wire  _GEN647 = io_x[26] ? _GEN646 : _GEN643;
wire  _GEN648 = io_x[22] ? _GEN647 : _GEN641;
wire  _GEN649 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN650 = io_x[30] ? _GEN649 : _GEN106;
wire  _GEN651 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN652 = io_x[30] ? _GEN651 : _GEN117;
wire  _GEN653 = io_x[26] ? _GEN652 : _GEN650;
wire  _GEN654 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN655 = io_x[30] ? _GEN654 : _GEN106;
wire  _GEN656 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN657 = io_x[30] ? _GEN656 : _GEN117;
wire  _GEN658 = io_x[26] ? _GEN657 : _GEN655;
wire  _GEN659 = io_x[22] ? _GEN658 : _GEN653;
wire  _GEN660 = io_x[13] ? _GEN659 : _GEN648;
wire  _GEN661 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN662 = io_x[30] ? _GEN117 : _GEN661;
wire  _GEN663 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN664 = io_x[30] ? _GEN106 : _GEN663;
wire  _GEN665 = io_x[26] ? _GEN664 : _GEN662;
wire  _GEN666 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN667 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN668 = io_x[30] ? _GEN667 : _GEN666;
wire  _GEN669 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN670 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN671 = io_x[30] ? _GEN670 : _GEN669;
wire  _GEN672 = io_x[26] ? _GEN671 : _GEN668;
wire  _GEN673 = io_x[22] ? _GEN672 : _GEN665;
wire  _GEN674 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN675 = io_x[30] ? _GEN674 : _GEN106;
wire  _GEN676 = io_x[26] ? _GEN675 : _GEN108;
wire  _GEN677 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN678 = io_x[30] ? _GEN677 : _GEN117;
wire  _GEN679 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN680 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN681 = io_x[30] ? _GEN680 : _GEN679;
wire  _GEN682 = io_x[26] ? _GEN681 : _GEN678;
wire  _GEN683 = io_x[22] ? _GEN682 : _GEN676;
wire  _GEN684 = io_x[13] ? _GEN683 : _GEN673;
wire  _GEN685 = io_x[33] ? _GEN684 : _GEN660;
wire  _GEN686 = io_x[69] ? _GEN685 : _GEN636;
wire  _GEN687 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN688 = io_x[30] ? _GEN117 : _GEN687;
wire  _GEN689 = io_x[26] ? _GEN119 : _GEN688;
wire  _GEN690 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN691 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN692 = io_x[30] ? _GEN691 : _GEN690;
wire  _GEN693 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN694 = io_x[30] ? _GEN117 : _GEN693;
wire  _GEN695 = io_x[26] ? _GEN694 : _GEN692;
wire  _GEN696 = io_x[22] ? _GEN695 : _GEN689;
wire  _GEN697 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN698 = io_x[26] ? _GEN697 : _GEN119;
wire  _GEN699 = io_x[22] ? _GEN698 : _GEN314;
wire  _GEN700 = io_x[13] ? _GEN699 : _GEN696;
wire  _GEN701 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN702 = io_x[30] ? _GEN117 : _GEN701;
wire  _GEN703 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN704 = io_x[30] ? _GEN703 : _GEN106;
wire  _GEN705 = io_x[26] ? _GEN704 : _GEN702;
wire  _GEN706 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN707 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN708 = io_x[30] ? _GEN707 : _GEN706;
wire  _GEN709 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN710 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN711 = io_x[30] ? _GEN710 : _GEN709;
wire  _GEN712 = io_x[26] ? _GEN711 : _GEN708;
wire  _GEN713 = io_x[22] ? _GEN712 : _GEN705;
wire  _GEN714 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN715 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN716 = io_x[30] ? _GEN715 : _GEN117;
wire  _GEN717 = io_x[26] ? _GEN716 : _GEN714;
wire  _GEN718 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN719 = io_x[30] ? _GEN718 : _GEN117;
wire  _GEN720 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN721 = io_x[26] ? _GEN720 : _GEN719;
wire  _GEN722 = io_x[22] ? _GEN721 : _GEN717;
wire  _GEN723 = io_x[13] ? _GEN722 : _GEN713;
wire  _GEN724 = io_x[33] ? _GEN723 : _GEN700;
wire  _GEN725 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN726 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN727 = io_x[30] ? _GEN726 : _GEN725;
wire  _GEN728 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN729 = io_x[30] ? _GEN117 : _GEN728;
wire  _GEN730 = io_x[26] ? _GEN729 : _GEN727;
wire  _GEN731 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN732 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN733 = io_x[26] ? _GEN732 : _GEN731;
wire  _GEN734 = io_x[22] ? _GEN733 : _GEN730;
wire  _GEN735 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN736 = io_x[30] ? _GEN735 : _GEN117;
wire  _GEN737 = io_x[26] ? _GEN119 : _GEN736;
wire  _GEN738 = io_x[22] ? _GEN204 : _GEN737;
wire  _GEN739 = io_x[13] ? _GEN738 : _GEN734;
wire  _GEN740 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN741 = io_x[30] ? _GEN106 : _GEN740;
wire  _GEN742 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN743 = io_x[30] ? _GEN117 : _GEN742;
wire  _GEN744 = io_x[26] ? _GEN743 : _GEN741;
wire  _GEN745 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN746 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN747 = io_x[30] ? _GEN746 : _GEN745;
wire  _GEN748 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN749 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN750 = io_x[30] ? _GEN749 : _GEN748;
wire  _GEN751 = io_x[26] ? _GEN750 : _GEN747;
wire  _GEN752 = io_x[22] ? _GEN751 : _GEN744;
wire  _GEN753 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN754 = io_x[30] ? _GEN753 : _GEN117;
wire  _GEN755 = io_x[26] ? _GEN754 : _GEN119;
wire  _GEN756 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN757 = io_x[30] ? _GEN756 : _GEN117;
wire  _GEN758 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN759 = io_x[30] ? _GEN758 : _GEN117;
wire  _GEN760 = io_x[26] ? _GEN759 : _GEN757;
wire  _GEN761 = io_x[22] ? _GEN760 : _GEN755;
wire  _GEN762 = io_x[13] ? _GEN761 : _GEN752;
wire  _GEN763 = io_x[33] ? _GEN762 : _GEN739;
wire  _GEN764 = io_x[69] ? _GEN763 : _GEN724;
wire  _GEN765 = io_x[71] ? _GEN764 : _GEN686;
wire  _GEN766 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN767 = io_x[30] ? _GEN106 : _GEN766;
wire  _GEN768 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN769 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN770 = io_x[30] ? _GEN769 : _GEN768;
wire  _GEN771 = io_x[26] ? _GEN770 : _GEN767;
wire  _GEN772 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN773 = io_x[30] ? _GEN117 : _GEN772;
wire  _GEN774 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN775 = io_x[30] ? _GEN117 : _GEN774;
wire  _GEN776 = io_x[26] ? _GEN775 : _GEN773;
wire  _GEN777 = io_x[22] ? _GEN776 : _GEN771;
wire  _GEN778 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN779 = io_x[30] ? _GEN778 : _GEN117;
wire  _GEN780 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN781 = io_x[30] ? _GEN117 : _GEN780;
wire  _GEN782 = io_x[26] ? _GEN781 : _GEN779;
wire  _GEN783 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN784 = io_x[30] ? _GEN783 : _GEN106;
wire  _GEN785 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN786 = io_x[30] ? _GEN785 : _GEN117;
wire  _GEN787 = io_x[26] ? _GEN786 : _GEN784;
wire  _GEN788 = io_x[22] ? _GEN787 : _GEN782;
wire  _GEN789 = io_x[13] ? _GEN788 : _GEN777;
wire  _GEN790 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN791 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN792 = io_x[30] ? _GEN791 : _GEN790;
wire  _GEN793 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN794 = io_x[30] ? _GEN117 : _GEN793;
wire  _GEN795 = io_x[26] ? _GEN794 : _GEN792;
wire  _GEN796 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN797 = io_x[30] ? _GEN117 : _GEN796;
wire  _GEN798 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN799 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN800 = io_x[30] ? _GEN799 : _GEN798;
wire  _GEN801 = io_x[26] ? _GEN800 : _GEN797;
wire  _GEN802 = io_x[22] ? _GEN801 : _GEN795;
wire  _GEN803 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN804 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN805 = io_x[30] ? _GEN804 : _GEN803;
wire  _GEN806 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN807 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN808 = io_x[30] ? _GEN807 : _GEN806;
wire  _GEN809 = io_x[26] ? _GEN808 : _GEN805;
wire  _GEN810 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN811 = io_x[30] ? _GEN106 : _GEN810;
wire  _GEN812 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN813 = io_x[30] ? _GEN812 : _GEN106;
wire  _GEN814 = io_x[26] ? _GEN813 : _GEN811;
wire  _GEN815 = io_x[22] ? _GEN814 : _GEN809;
wire  _GEN816 = io_x[13] ? _GEN815 : _GEN802;
wire  _GEN817 = io_x[33] ? _GEN816 : _GEN789;
wire  _GEN818 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN819 = io_x[30] ? _GEN117 : _GEN818;
wire  _GEN820 = io_x[26] ? _GEN119 : _GEN819;
wire  _GEN821 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN822 = io_x[30] ? _GEN821 : _GEN117;
wire  _GEN823 = io_x[26] ? _GEN822 : _GEN119;
wire  _GEN824 = io_x[22] ? _GEN823 : _GEN820;
wire  _GEN825 = io_x[26] ? _GEN108 : _GEN119;
wire  _GEN826 = io_x[22] ? _GEN314 : _GEN825;
wire  _GEN827 = io_x[13] ? _GEN826 : _GEN824;
wire  _GEN828 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN829 = io_x[30] ? _GEN106 : _GEN828;
wire  _GEN830 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN831 = io_x[30] ? _GEN830 : _GEN106;
wire  _GEN832 = io_x[26] ? _GEN831 : _GEN829;
wire  _GEN833 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN834 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN835 = io_x[30] ? _GEN106 : _GEN834;
wire  _GEN836 = io_x[26] ? _GEN835 : _GEN833;
wire  _GEN837 = io_x[22] ? _GEN836 : _GEN832;
wire  _GEN838 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN839 = io_x[30] ? _GEN838 : _GEN117;
wire  _GEN840 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN841 = io_x[26] ? _GEN840 : _GEN839;
wire  _GEN842 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN843 = io_x[30] ? _GEN842 : _GEN106;
wire  _GEN844 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN845 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN846 = io_x[30] ? _GEN845 : _GEN844;
wire  _GEN847 = io_x[26] ? _GEN846 : _GEN843;
wire  _GEN848 = io_x[22] ? _GEN847 : _GEN841;
wire  _GEN849 = io_x[13] ? _GEN848 : _GEN837;
wire  _GEN850 = io_x[33] ? _GEN849 : _GEN827;
wire  _GEN851 = io_x[69] ? _GEN850 : _GEN817;
wire  _GEN852 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN853 = io_x[30] ? _GEN106 : _GEN852;
wire  _GEN854 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN855 = io_x[30] ? _GEN854 : _GEN106;
wire  _GEN856 = io_x[26] ? _GEN855 : _GEN853;
wire  _GEN857 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN858 = io_x[30] ? _GEN117 : _GEN857;
wire  _GEN859 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN860 = io_x[30] ? _GEN859 : _GEN117;
wire  _GEN861 = io_x[26] ? _GEN860 : _GEN858;
wire  _GEN862 = io_x[22] ? _GEN861 : _GEN856;
wire  _GEN863 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN864 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN865 = io_x[30] ? _GEN864 : _GEN863;
wire  _GEN866 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN867 = io_x[30] ? _GEN866 : _GEN117;
wire  _GEN868 = io_x[26] ? _GEN867 : _GEN865;
wire  _GEN869 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN870 = io_x[30] ? _GEN869 : _GEN117;
wire  _GEN871 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN872 = io_x[30] ? _GEN871 : _GEN106;
wire  _GEN873 = io_x[26] ? _GEN872 : _GEN870;
wire  _GEN874 = io_x[22] ? _GEN873 : _GEN868;
wire  _GEN875 = io_x[13] ? _GEN874 : _GEN862;
wire  _GEN876 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN877 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN878 = io_x[30] ? _GEN877 : _GEN876;
wire  _GEN879 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN880 = io_x[30] ? _GEN117 : _GEN879;
wire  _GEN881 = io_x[26] ? _GEN880 : _GEN878;
wire  _GEN882 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN883 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN884 = io_x[30] ? _GEN883 : _GEN882;
wire  _GEN885 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN886 = io_x[30] ? _GEN885 : _GEN117;
wire  _GEN887 = io_x[26] ? _GEN886 : _GEN884;
wire  _GEN888 = io_x[22] ? _GEN887 : _GEN881;
wire  _GEN889 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN890 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN891 = io_x[30] ? _GEN890 : _GEN889;
wire  _GEN892 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN893 = io_x[30] ? _GEN892 : _GEN117;
wire  _GEN894 = io_x[26] ? _GEN893 : _GEN891;
wire  _GEN895 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN896 = io_x[30] ? _GEN895 : _GEN117;
wire  _GEN897 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN898 = io_x[30] ? _GEN897 : _GEN117;
wire  _GEN899 = io_x[26] ? _GEN898 : _GEN896;
wire  _GEN900 = io_x[22] ? _GEN899 : _GEN894;
wire  _GEN901 = io_x[13] ? _GEN900 : _GEN888;
wire  _GEN902 = io_x[33] ? _GEN901 : _GEN875;
wire  _GEN903 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN904 = io_x[30] ? _GEN106 : _GEN903;
wire  _GEN905 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN906 = io_x[30] ? _GEN905 : _GEN106;
wire  _GEN907 = io_x[26] ? _GEN906 : _GEN904;
wire  _GEN908 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN909 = io_x[30] ? _GEN117 : _GEN908;
wire  _GEN910 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN911 = io_x[30] ? _GEN106 : _GEN910;
wire  _GEN912 = io_x[26] ? _GEN911 : _GEN909;
wire  _GEN913 = io_x[22] ? _GEN912 : _GEN907;
wire  _GEN914 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN915 = io_x[30] ? _GEN106 : _GEN914;
wire  _GEN916 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN917 = io_x[30] ? _GEN117 : _GEN916;
wire  _GEN918 = io_x[26] ? _GEN917 : _GEN915;
wire  _GEN919 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN920 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN921 = io_x[30] ? _GEN920 : _GEN117;
wire  _GEN922 = io_x[26] ? _GEN921 : _GEN919;
wire  _GEN923 = io_x[22] ? _GEN922 : _GEN918;
wire  _GEN924 = io_x[13] ? _GEN923 : _GEN913;
wire  _GEN925 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN926 = io_x[30] ? _GEN106 : _GEN925;
wire  _GEN927 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN928 = io_x[30] ? _GEN106 : _GEN927;
wire  _GEN929 = io_x[26] ? _GEN928 : _GEN926;
wire  _GEN930 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN931 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN932 = io_x[30] ? _GEN931 : _GEN930;
wire  _GEN933 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN934 = io_x[30] ? _GEN117 : _GEN933;
wire  _GEN935 = io_x[26] ? _GEN934 : _GEN932;
wire  _GEN936 = io_x[22] ? _GEN935 : _GEN929;
wire  _GEN937 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN938 = io_x[30] ? _GEN937 : _GEN117;
wire  _GEN939 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN940 = io_x[30] ? _GEN939 : _GEN106;
wire  _GEN941 = io_x[26] ? _GEN940 : _GEN938;
wire  _GEN942 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN943 = io_x[30] ? _GEN942 : _GEN117;
wire  _GEN944 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN945 = io_x[30] ? _GEN944 : _GEN106;
wire  _GEN946 = io_x[26] ? _GEN945 : _GEN943;
wire  _GEN947 = io_x[22] ? _GEN946 : _GEN941;
wire  _GEN948 = io_x[13] ? _GEN947 : _GEN936;
wire  _GEN949 = io_x[33] ? _GEN948 : _GEN924;
wire  _GEN950 = io_x[69] ? _GEN949 : _GEN902;
wire  _GEN951 = io_x[71] ? _GEN950 : _GEN851;
wire  _GEN952 = io_x[72] ? _GEN951 : _GEN765;
wire  _GEN953 = io_x[13] ? _GEN563 : _GEN523;
wire  _GEN954 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN955 = io_x[30] ? _GEN117 : _GEN954;
wire  _GEN956 = io_x[26] ? _GEN108 : _GEN955;
wire  _GEN957 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN958 = io_x[30] ? _GEN117 : _GEN957;
wire  _GEN959 = io_x[26] ? _GEN958 : _GEN108;
wire  _GEN960 = io_x[22] ? _GEN959 : _GEN956;
wire  _GEN961 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN962 = io_x[30] ? _GEN961 : _GEN117;
wire  _GEN963 = io_x[26] ? _GEN962 : _GEN108;
wire  _GEN964 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN965 = io_x[26] ? _GEN964 : _GEN119;
wire  _GEN966 = io_x[22] ? _GEN965 : _GEN963;
wire  _GEN967 = io_x[13] ? _GEN966 : _GEN960;
wire  _GEN968 = io_x[33] ? _GEN967 : _GEN953;
wire  _GEN969 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN970 = io_x[30] ? _GEN106 : _GEN969;
wire  _GEN971 = io_x[26] ? _GEN108 : _GEN970;
wire  _GEN972 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN973 = io_x[22] ? _GEN972 : _GEN971;
wire  _GEN974 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN975 = io_x[26] ? _GEN974 : _GEN119;
wire  _GEN976 = io_x[22] ? _GEN975 : _GEN204;
wire  _GEN977 = io_x[13] ? _GEN976 : _GEN973;
wire  _GEN978 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN979 = io_x[30] ? _GEN117 : _GEN978;
wire  _GEN980 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN981 = io_x[30] ? _GEN980 : _GEN106;
wire  _GEN982 = io_x[26] ? _GEN981 : _GEN979;
wire  _GEN983 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN984 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN985 = io_x[30] ? _GEN117 : _GEN984;
wire  _GEN986 = io_x[26] ? _GEN985 : _GEN983;
wire  _GEN987 = io_x[22] ? _GEN986 : _GEN982;
wire  _GEN988 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN989 = io_x[30] ? _GEN117 : _GEN988;
wire  _GEN990 = io_x[26] ? _GEN119 : _GEN989;
wire  _GEN991 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN992 = io_x[30] ? _GEN991 : _GEN117;
wire  _GEN993 = io_x[26] ? _GEN992 : _GEN119;
wire  _GEN994 = io_x[22] ? _GEN993 : _GEN990;
wire  _GEN995 = io_x[13] ? _GEN994 : _GEN987;
wire  _GEN996 = io_x[33] ? _GEN995 : _GEN977;
wire  _GEN997 = io_x[69] ? _GEN996 : _GEN968;
wire  _GEN998 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN999 = io_x[30] ? _GEN117 : _GEN998;
wire  _GEN1000 = io_x[26] ? _GEN119 : _GEN999;
wire  _GEN1001 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN1002 = io_x[22] ? _GEN1001 : _GEN1000;
wire  _GEN1003 = io_x[22] ? _GEN314 : _GEN204;
wire  _GEN1004 = io_x[13] ? _GEN1003 : _GEN1002;
wire  _GEN1005 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1006 = io_x[26] ? _GEN1005 : _GEN108;
wire  _GEN1007 = io_x[22] ? _GEN1006 : _GEN314;
wire  _GEN1008 = io_x[13] ? _GEN523 : _GEN1007;
wire  _GEN1009 = io_x[33] ? _GEN1008 : _GEN1004;
wire  _GEN1010 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1011 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1012 = io_x[26] ? _GEN1011 : _GEN1010;
wire  _GEN1013 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1014 = io_x[30] ? _GEN117 : _GEN1013;
wire  _GEN1015 = io_x[26] ? _GEN1014 : _GEN108;
wire  _GEN1016 = io_x[22] ? _GEN1015 : _GEN1012;
wire  _GEN1017 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN1018 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1019 = io_x[30] ? _GEN1018 : _GEN117;
wire  _GEN1020 = io_x[26] ? _GEN1019 : _GEN119;
wire  _GEN1021 = io_x[22] ? _GEN1020 : _GEN1017;
wire  _GEN1022 = io_x[13] ? _GEN1021 : _GEN1016;
wire  _GEN1023 = io_x[26] ? _GEN108 : _GEN119;
wire  _GEN1024 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1025 = io_x[30] ? _GEN1024 : _GEN106;
wire  _GEN1026 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1027 = io_x[30] ? _GEN1026 : _GEN117;
wire  _GEN1028 = io_x[26] ? _GEN1027 : _GEN1025;
wire  _GEN1029 = io_x[22] ? _GEN1028 : _GEN1023;
wire  _GEN1030 = io_x[22] ? _GEN314 : _GEN204;
wire  _GEN1031 = io_x[13] ? _GEN1030 : _GEN1029;
wire  _GEN1032 = io_x[33] ? _GEN1031 : _GEN1022;
wire  _GEN1033 = io_x[69] ? _GEN1032 : _GEN1009;
wire  _GEN1034 = io_x[71] ? _GEN1033 : _GEN997;
wire  _GEN1035 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1036 = io_x[30] ? _GEN106 : _GEN1035;
wire  _GEN1037 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1038 = io_x[26] ? _GEN1037 : _GEN1036;
wire  _GEN1039 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1040 = io_x[26] ? _GEN119 : _GEN1039;
wire  _GEN1041 = io_x[22] ? _GEN1040 : _GEN1038;
wire  _GEN1042 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1043 = io_x[26] ? _GEN119 : _GEN1042;
wire  _GEN1044 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1045 = io_x[26] ? _GEN119 : _GEN1044;
wire  _GEN1046 = io_x[22] ? _GEN1045 : _GEN1043;
wire  _GEN1047 = io_x[13] ? _GEN1046 : _GEN1041;
wire  _GEN1048 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1049 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1050 = io_x[30] ? _GEN117 : _GEN1049;
wire  _GEN1051 = io_x[26] ? _GEN1050 : _GEN1048;
wire  _GEN1052 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1053 = io_x[30] ? _GEN1052 : _GEN117;
wire  _GEN1054 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1055 = io_x[26] ? _GEN1054 : _GEN1053;
wire  _GEN1056 = io_x[22] ? _GEN1055 : _GEN1051;
wire  _GEN1057 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1058 = io_x[30] ? _GEN1057 : _GEN106;
wire  _GEN1059 = io_x[26] ? _GEN108 : _GEN1058;
wire  _GEN1060 = io_x[22] ? _GEN1059 : _GEN204;
wire  _GEN1061 = io_x[13] ? _GEN1060 : _GEN1056;
wire  _GEN1062 = io_x[33] ? _GEN1061 : _GEN1047;
wire  _GEN1063 = io_x[13] ? _GEN563 : _GEN523;
wire  _GEN1064 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1065 = io_x[30] ? _GEN117 : _GEN1064;
wire  _GEN1066 = io_x[26] ? _GEN108 : _GEN1065;
wire  _GEN1067 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1068 = io_x[30] ? _GEN106 : _GEN1067;
wire  _GEN1069 = io_x[26] ? _GEN119 : _GEN1068;
wire  _GEN1070 = io_x[22] ? _GEN1069 : _GEN1066;
wire  _GEN1071 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1072 = io_x[30] ? _GEN1071 : _GEN117;
wire  _GEN1073 = io_x[26] ? _GEN1072 : _GEN108;
wire  _GEN1074 = io_x[22] ? _GEN1073 : _GEN204;
wire  _GEN1075 = io_x[13] ? _GEN1074 : _GEN1070;
wire  _GEN1076 = io_x[33] ? _GEN1075 : _GEN1063;
wire  _GEN1077 = io_x[69] ? _GEN1076 : _GEN1062;
wire  _GEN1078 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1079 = io_x[26] ? _GEN1078 : _GEN119;
wire  _GEN1080 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN1081 = io_x[22] ? _GEN1080 : _GEN1079;
wire  _GEN1082 = io_x[13] ? _GEN563 : _GEN1081;
wire  _GEN1083 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1084 = io_x[30] ? _GEN117 : _GEN1083;
wire  _GEN1085 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1086 = io_x[26] ? _GEN1085 : _GEN1084;
wire  _GEN1087 = io_x[22] ? _GEN1086 : _GEN204;
wire  _GEN1088 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN1089 = io_x[22] ? _GEN314 : _GEN1088;
wire  _GEN1090 = io_x[13] ? _GEN1089 : _GEN1087;
wire  _GEN1091 = io_x[33] ? _GEN1090 : _GEN1082;
wire  _GEN1092 = io_x[26] ? _GEN108 : _GEN119;
wire  _GEN1093 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1094 = io_x[30] ? _GEN1093 : _GEN117;
wire  _GEN1095 = io_x[26] ? _GEN1094 : _GEN119;
wire  _GEN1096 = io_x[22] ? _GEN1095 : _GEN1092;
wire  _GEN1097 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN1098 = io_x[22] ? _GEN1097 : _GEN314;
wire  _GEN1099 = io_x[13] ? _GEN1098 : _GEN1096;
wire  _GEN1100 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1101 = io_x[30] ? _GEN117 : _GEN1100;
wire  _GEN1102 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1103 = io_x[30] ? _GEN117 : _GEN1102;
wire  _GEN1104 = io_x[26] ? _GEN1103 : _GEN1101;
wire  _GEN1105 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1106 = io_x[30] ? _GEN117 : _GEN1105;
wire  _GEN1107 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1108 = io_x[26] ? _GEN1107 : _GEN1106;
wire  _GEN1109 = io_x[22] ? _GEN1108 : _GEN1104;
wire  _GEN1110 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1111 = io_x[30] ? _GEN1110 : _GEN117;
wire  _GEN1112 = io_x[26] ? _GEN119 : _GEN1111;
wire  _GEN1113 = io_x[22] ? _GEN1112 : _GEN314;
wire  _GEN1114 = io_x[13] ? _GEN1113 : _GEN1109;
wire  _GEN1115 = io_x[33] ? _GEN1114 : _GEN1099;
wire  _GEN1116 = io_x[69] ? _GEN1115 : _GEN1091;
wire  _GEN1117 = io_x[71] ? _GEN1116 : _GEN1077;
wire  _GEN1118 = io_x[72] ? _GEN1117 : _GEN1034;
wire  _GEN1119 = io_x[48] ? _GEN1118 : _GEN952;
wire  _GEN1120 = io_x[32] ? _GEN1119 : _GEN602;
wire  _GEN1121 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1122 = io_x[30] ? _GEN117 : _GEN1121;
wire  _GEN1123 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1124 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1125 = io_x[30] ? _GEN1124 : _GEN1123;
wire  _GEN1126 = io_x[26] ? _GEN1125 : _GEN1122;
wire  _GEN1127 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1128 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1129 = io_x[30] ? _GEN1128 : _GEN1127;
wire  _GEN1130 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1131 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1132 = io_x[30] ? _GEN1131 : _GEN1130;
wire  _GEN1133 = io_x[26] ? _GEN1132 : _GEN1129;
wire  _GEN1134 = io_x[22] ? _GEN1133 : _GEN1126;
wire  _GEN1135 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1136 = io_x[30] ? _GEN1135 : _GEN106;
wire  _GEN1137 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1138 = io_x[30] ? _GEN1137 : _GEN106;
wire  _GEN1139 = io_x[26] ? _GEN1138 : _GEN1136;
wire  _GEN1140 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1141 = io_x[30] ? _GEN1140 : _GEN106;
wire  _GEN1142 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1143 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1144 = io_x[30] ? _GEN1143 : _GEN1142;
wire  _GEN1145 = io_x[26] ? _GEN1144 : _GEN1141;
wire  _GEN1146 = io_x[22] ? _GEN1145 : _GEN1139;
wire  _GEN1147 = io_x[13] ? _GEN1146 : _GEN1134;
wire  _GEN1148 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1149 = io_x[30] ? _GEN117 : _GEN1148;
wire  _GEN1150 = io_x[26] ? _GEN1149 : _GEN108;
wire  _GEN1151 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1152 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1153 = io_x[30] ? _GEN1152 : _GEN1151;
wire  _GEN1154 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1155 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1156 = io_x[30] ? _GEN1155 : _GEN1154;
wire  _GEN1157 = io_x[26] ? _GEN1156 : _GEN1153;
wire  _GEN1158 = io_x[22] ? _GEN1157 : _GEN1150;
wire  _GEN1159 = io_x[26] ? _GEN108 : _GEN119;
wire  _GEN1160 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1161 = io_x[30] ? _GEN1160 : _GEN117;
wire  _GEN1162 = io_x[26] ? _GEN1161 : _GEN119;
wire  _GEN1163 = io_x[22] ? _GEN1162 : _GEN1159;
wire  _GEN1164 = io_x[13] ? _GEN1163 : _GEN1158;
wire  _GEN1165 = io_x[33] ? _GEN1164 : _GEN1147;
wire  _GEN1166 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1167 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1168 = io_x[30] ? _GEN1167 : _GEN1166;
wire  _GEN1169 = io_x[26] ? _GEN119 : _GEN1168;
wire  _GEN1170 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1171 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1172 = io_x[30] ? _GEN1171 : _GEN1170;
wire  _GEN1173 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1174 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1175 = io_x[30] ? _GEN1174 : _GEN1173;
wire  _GEN1176 = io_x[26] ? _GEN1175 : _GEN1172;
wire  _GEN1177 = io_x[22] ? _GEN1176 : _GEN1169;
wire  _GEN1178 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1179 = io_x[30] ? _GEN1178 : _GEN106;
wire  _GEN1180 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1181 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1182 = io_x[30] ? _GEN1181 : _GEN1180;
wire  _GEN1183 = io_x[26] ? _GEN1182 : _GEN1179;
wire  _GEN1184 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1185 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1186 = io_x[30] ? _GEN1185 : _GEN1184;
wire  _GEN1187 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1188 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1189 = io_x[30] ? _GEN1188 : _GEN1187;
wire  _GEN1190 = io_x[26] ? _GEN1189 : _GEN1186;
wire  _GEN1191 = io_x[22] ? _GEN1190 : _GEN1183;
wire  _GEN1192 = io_x[13] ? _GEN1191 : _GEN1177;
wire  _GEN1193 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1194 = io_x[30] ? _GEN117 : _GEN1193;
wire  _GEN1195 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1196 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1197 = io_x[30] ? _GEN1196 : _GEN1195;
wire  _GEN1198 = io_x[26] ? _GEN1197 : _GEN1194;
wire  _GEN1199 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1200 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1201 = io_x[30] ? _GEN1200 : _GEN1199;
wire  _GEN1202 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1203 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1204 = io_x[30] ? _GEN1203 : _GEN1202;
wire  _GEN1205 = io_x[26] ? _GEN1204 : _GEN1201;
wire  _GEN1206 = io_x[22] ? _GEN1205 : _GEN1198;
wire  _GEN1207 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1208 = io_x[30] ? _GEN1207 : _GEN117;
wire  _GEN1209 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1210 = io_x[30] ? _GEN1209 : _GEN117;
wire  _GEN1211 = io_x[26] ? _GEN1210 : _GEN1208;
wire  _GEN1212 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1213 = io_x[30] ? _GEN1212 : _GEN106;
wire  _GEN1214 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1215 = io_x[30] ? _GEN1214 : _GEN117;
wire  _GEN1216 = io_x[26] ? _GEN1215 : _GEN1213;
wire  _GEN1217 = io_x[22] ? _GEN1216 : _GEN1211;
wire  _GEN1218 = io_x[13] ? _GEN1217 : _GEN1206;
wire  _GEN1219 = io_x[33] ? _GEN1218 : _GEN1192;
wire  _GEN1220 = io_x[69] ? _GEN1219 : _GEN1165;
wire  _GEN1221 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1222 = io_x[30] ? _GEN117 : _GEN1221;
wire  _GEN1223 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1224 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1225 = io_x[30] ? _GEN1224 : _GEN1223;
wire  _GEN1226 = io_x[26] ? _GEN1225 : _GEN1222;
wire  _GEN1227 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1228 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1229 = io_x[30] ? _GEN1228 : _GEN1227;
wire  _GEN1230 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1231 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1232 = io_x[30] ? _GEN1231 : _GEN1230;
wire  _GEN1233 = io_x[26] ? _GEN1232 : _GEN1229;
wire  _GEN1234 = io_x[22] ? _GEN1233 : _GEN1226;
wire  _GEN1235 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1236 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1237 = io_x[30] ? _GEN1236 : _GEN106;
wire  _GEN1238 = io_x[26] ? _GEN1237 : _GEN1235;
wire  _GEN1239 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1240 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1241 = io_x[30] ? _GEN1240 : _GEN1239;
wire  _GEN1242 = io_x[26] ? _GEN1241 : _GEN108;
wire  _GEN1243 = io_x[22] ? _GEN1242 : _GEN1238;
wire  _GEN1244 = io_x[13] ? _GEN1243 : _GEN1234;
wire  _GEN1245 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1246 = io_x[30] ? _GEN117 : _GEN1245;
wire  _GEN1247 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1248 = io_x[30] ? _GEN106 : _GEN1247;
wire  _GEN1249 = io_x[26] ? _GEN1248 : _GEN1246;
wire  _GEN1250 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1251 = io_x[30] ? _GEN1250 : _GEN117;
wire  _GEN1252 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1253 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1254 = io_x[30] ? _GEN1253 : _GEN1252;
wire  _GEN1255 = io_x[26] ? _GEN1254 : _GEN1251;
wire  _GEN1256 = io_x[22] ? _GEN1255 : _GEN1249;
wire  _GEN1257 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1258 = io_x[30] ? _GEN1257 : _GEN117;
wire  _GEN1259 = io_x[26] ? _GEN1258 : _GEN108;
wire  _GEN1260 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1261 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1262 = io_x[30] ? _GEN1261 : _GEN117;
wire  _GEN1263 = io_x[26] ? _GEN1262 : _GEN1260;
wire  _GEN1264 = io_x[22] ? _GEN1263 : _GEN1259;
wire  _GEN1265 = io_x[13] ? _GEN1264 : _GEN1256;
wire  _GEN1266 = io_x[33] ? _GEN1265 : _GEN1244;
wire  _GEN1267 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1268 = io_x[30] ? _GEN117 : _GEN1267;
wire  _GEN1269 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1270 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1271 = io_x[30] ? _GEN1270 : _GEN1269;
wire  _GEN1272 = io_x[26] ? _GEN1271 : _GEN1268;
wire  _GEN1273 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1274 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1275 = io_x[30] ? _GEN1274 : _GEN1273;
wire  _GEN1276 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1277 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1278 = io_x[30] ? _GEN1277 : _GEN1276;
wire  _GEN1279 = io_x[26] ? _GEN1278 : _GEN1275;
wire  _GEN1280 = io_x[22] ? _GEN1279 : _GEN1272;
wire  _GEN1281 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1282 = io_x[30] ? _GEN1281 : _GEN117;
wire  _GEN1283 = io_x[26] ? _GEN1282 : _GEN119;
wire  _GEN1284 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1285 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1286 = io_x[30] ? _GEN1285 : _GEN1284;
wire  _GEN1287 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1288 = io_x[30] ? _GEN1287 : _GEN106;
wire  _GEN1289 = io_x[26] ? _GEN1288 : _GEN1286;
wire  _GEN1290 = io_x[22] ? _GEN1289 : _GEN1283;
wire  _GEN1291 = io_x[13] ? _GEN1290 : _GEN1280;
wire  _GEN1292 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1293 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1294 = io_x[30] ? _GEN1293 : _GEN117;
wire  _GEN1295 = io_x[26] ? _GEN1294 : _GEN1292;
wire  _GEN1296 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1297 = io_x[30] ? _GEN1296 : _GEN117;
wire  _GEN1298 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1299 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1300 = io_x[30] ? _GEN1299 : _GEN1298;
wire  _GEN1301 = io_x[26] ? _GEN1300 : _GEN1297;
wire  _GEN1302 = io_x[22] ? _GEN1301 : _GEN1295;
wire  _GEN1303 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1304 = io_x[30] ? _GEN1303 : _GEN117;
wire  _GEN1305 = io_x[26] ? _GEN1304 : _GEN108;
wire  _GEN1306 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1307 = io_x[30] ? _GEN1306 : _GEN117;
wire  _GEN1308 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1309 = io_x[30] ? _GEN1308 : _GEN106;
wire  _GEN1310 = io_x[26] ? _GEN1309 : _GEN1307;
wire  _GEN1311 = io_x[22] ? _GEN1310 : _GEN1305;
wire  _GEN1312 = io_x[13] ? _GEN1311 : _GEN1302;
wire  _GEN1313 = io_x[33] ? _GEN1312 : _GEN1291;
wire  _GEN1314 = io_x[69] ? _GEN1313 : _GEN1266;
wire  _GEN1315 = io_x[71] ? _GEN1314 : _GEN1220;
wire  _GEN1316 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1317 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1318 = io_x[30] ? _GEN1317 : _GEN1316;
wire  _GEN1319 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1320 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1321 = io_x[30] ? _GEN1320 : _GEN1319;
wire  _GEN1322 = io_x[26] ? _GEN1321 : _GEN1318;
wire  _GEN1323 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1324 = io_x[30] ? _GEN106 : _GEN1323;
wire  _GEN1325 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1326 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1327 = io_x[30] ? _GEN1326 : _GEN1325;
wire  _GEN1328 = io_x[26] ? _GEN1327 : _GEN1324;
wire  _GEN1329 = io_x[22] ? _GEN1328 : _GEN1322;
wire  _GEN1330 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1331 = io_x[30] ? _GEN117 : _GEN1330;
wire  _GEN1332 = io_x[26] ? _GEN119 : _GEN1331;
wire  _GEN1333 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1334 = io_x[30] ? _GEN1333 : _GEN117;
wire  _GEN1335 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1336 = io_x[30] ? _GEN1335 : _GEN106;
wire  _GEN1337 = io_x[26] ? _GEN1336 : _GEN1334;
wire  _GEN1338 = io_x[22] ? _GEN1337 : _GEN1332;
wire  _GEN1339 = io_x[13] ? _GEN1338 : _GEN1329;
wire  _GEN1340 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1341 = io_x[30] ? _GEN117 : _GEN1340;
wire  _GEN1342 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1343 = io_x[30] ? _GEN117 : _GEN1342;
wire  _GEN1344 = io_x[26] ? _GEN1343 : _GEN1341;
wire  _GEN1345 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1346 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1347 = io_x[30] ? _GEN1346 : _GEN1345;
wire  _GEN1348 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1349 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1350 = io_x[30] ? _GEN1349 : _GEN1348;
wire  _GEN1351 = io_x[26] ? _GEN1350 : _GEN1347;
wire  _GEN1352 = io_x[22] ? _GEN1351 : _GEN1344;
wire  _GEN1353 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1354 = io_x[30] ? _GEN1353 : _GEN106;
wire  _GEN1355 = io_x[26] ? _GEN1354 : _GEN108;
wire  _GEN1356 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1357 = io_x[30] ? _GEN1356 : _GEN117;
wire  _GEN1358 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1359 = io_x[30] ? _GEN1358 : _GEN117;
wire  _GEN1360 = io_x[26] ? _GEN1359 : _GEN1357;
wire  _GEN1361 = io_x[22] ? _GEN1360 : _GEN1355;
wire  _GEN1362 = io_x[13] ? _GEN1361 : _GEN1352;
wire  _GEN1363 = io_x[33] ? _GEN1362 : _GEN1339;
wire  _GEN1364 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1365 = io_x[30] ? _GEN106 : _GEN1364;
wire  _GEN1366 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1367 = io_x[30] ? _GEN117 : _GEN1366;
wire  _GEN1368 = io_x[26] ? _GEN1367 : _GEN1365;
wire  _GEN1369 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1370 = io_x[30] ? _GEN117 : _GEN1369;
wire  _GEN1371 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1372 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1373 = io_x[30] ? _GEN1372 : _GEN1371;
wire  _GEN1374 = io_x[26] ? _GEN1373 : _GEN1370;
wire  _GEN1375 = io_x[22] ? _GEN1374 : _GEN1368;
wire  _GEN1376 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1377 = io_x[30] ? _GEN1376 : _GEN106;
wire  _GEN1378 = io_x[26] ? _GEN1377 : _GEN108;
wire  _GEN1379 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1380 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1381 = io_x[30] ? _GEN1380 : _GEN1379;
wire  _GEN1382 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1383 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1384 = io_x[30] ? _GEN1383 : _GEN1382;
wire  _GEN1385 = io_x[26] ? _GEN1384 : _GEN1381;
wire  _GEN1386 = io_x[22] ? _GEN1385 : _GEN1378;
wire  _GEN1387 = io_x[13] ? _GEN1386 : _GEN1375;
wire  _GEN1388 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1389 = io_x[30] ? _GEN106 : _GEN1388;
wire  _GEN1390 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1391 = io_x[26] ? _GEN1390 : _GEN1389;
wire  _GEN1392 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1393 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1394 = io_x[30] ? _GEN1393 : _GEN1392;
wire  _GEN1395 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1396 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1397 = io_x[30] ? _GEN1396 : _GEN1395;
wire  _GEN1398 = io_x[26] ? _GEN1397 : _GEN1394;
wire  _GEN1399 = io_x[22] ? _GEN1398 : _GEN1391;
wire  _GEN1400 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1401 = io_x[30] ? _GEN1400 : _GEN117;
wire  _GEN1402 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1403 = io_x[30] ? _GEN1402 : _GEN106;
wire  _GEN1404 = io_x[26] ? _GEN1403 : _GEN1401;
wire  _GEN1405 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1406 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1407 = io_x[30] ? _GEN1406 : _GEN106;
wire  _GEN1408 = io_x[26] ? _GEN1407 : _GEN1405;
wire  _GEN1409 = io_x[22] ? _GEN1408 : _GEN1404;
wire  _GEN1410 = io_x[13] ? _GEN1409 : _GEN1399;
wire  _GEN1411 = io_x[33] ? _GEN1410 : _GEN1387;
wire  _GEN1412 = io_x[69] ? _GEN1411 : _GEN1363;
wire  _GEN1413 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1414 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1415 = io_x[30] ? _GEN1414 : _GEN1413;
wire  _GEN1416 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1417 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1418 = io_x[30] ? _GEN1417 : _GEN1416;
wire  _GEN1419 = io_x[26] ? _GEN1418 : _GEN1415;
wire  _GEN1420 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1421 = io_x[30] ? _GEN117 : _GEN1420;
wire  _GEN1422 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1423 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1424 = io_x[30] ? _GEN1423 : _GEN1422;
wire  _GEN1425 = io_x[26] ? _GEN1424 : _GEN1421;
wire  _GEN1426 = io_x[22] ? _GEN1425 : _GEN1419;
wire  _GEN1427 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1428 = io_x[26] ? _GEN108 : _GEN1427;
wire  _GEN1429 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1430 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1431 = io_x[30] ? _GEN1430 : _GEN1429;
wire  _GEN1432 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1433 = io_x[30] ? _GEN1432 : _GEN106;
wire  _GEN1434 = io_x[26] ? _GEN1433 : _GEN1431;
wire  _GEN1435 = io_x[22] ? _GEN1434 : _GEN1428;
wire  _GEN1436 = io_x[13] ? _GEN1435 : _GEN1426;
wire  _GEN1437 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1438 = io_x[30] ? _GEN106 : _GEN1437;
wire  _GEN1439 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1440 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1441 = io_x[30] ? _GEN1440 : _GEN1439;
wire  _GEN1442 = io_x[26] ? _GEN1441 : _GEN1438;
wire  _GEN1443 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1444 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1445 = io_x[30] ? _GEN1444 : _GEN1443;
wire  _GEN1446 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1447 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1448 = io_x[30] ? _GEN1447 : _GEN1446;
wire  _GEN1449 = io_x[26] ? _GEN1448 : _GEN1445;
wire  _GEN1450 = io_x[22] ? _GEN1449 : _GEN1442;
wire  _GEN1451 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1452 = io_x[30] ? _GEN1451 : _GEN117;
wire  _GEN1453 = io_x[26] ? _GEN108 : _GEN1452;
wire  _GEN1454 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1455 = io_x[30] ? _GEN1454 : _GEN117;
wire  _GEN1456 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1457 = io_x[30] ? _GEN1456 : _GEN117;
wire  _GEN1458 = io_x[26] ? _GEN1457 : _GEN1455;
wire  _GEN1459 = io_x[22] ? _GEN1458 : _GEN1453;
wire  _GEN1460 = io_x[13] ? _GEN1459 : _GEN1450;
wire  _GEN1461 = io_x[33] ? _GEN1460 : _GEN1436;
wire  _GEN1462 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1463 = io_x[30] ? _GEN117 : _GEN1462;
wire  _GEN1464 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1465 = io_x[30] ? _GEN117 : _GEN1464;
wire  _GEN1466 = io_x[26] ? _GEN1465 : _GEN1463;
wire  _GEN1467 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1468 = io_x[30] ? _GEN117 : _GEN1467;
wire  _GEN1469 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1470 = io_x[30] ? _GEN106 : _GEN1469;
wire  _GEN1471 = io_x[26] ? _GEN1470 : _GEN1468;
wire  _GEN1472 = io_x[22] ? _GEN1471 : _GEN1466;
wire  _GEN1473 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1474 = io_x[30] ? _GEN1473 : _GEN106;
wire  _GEN1475 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1476 = io_x[30] ? _GEN1475 : _GEN117;
wire  _GEN1477 = io_x[26] ? _GEN1476 : _GEN1474;
wire  _GEN1478 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1479 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1480 = io_x[30] ? _GEN1479 : _GEN1478;
wire  _GEN1481 = io_x[26] ? _GEN1480 : _GEN119;
wire  _GEN1482 = io_x[22] ? _GEN1481 : _GEN1477;
wire  _GEN1483 = io_x[13] ? _GEN1482 : _GEN1472;
wire  _GEN1484 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1485 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1486 = io_x[30] ? _GEN1485 : _GEN1484;
wire  _GEN1487 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1488 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1489 = io_x[30] ? _GEN1488 : _GEN1487;
wire  _GEN1490 = io_x[26] ? _GEN1489 : _GEN1486;
wire  _GEN1491 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1492 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1493 = io_x[30] ? _GEN1492 : _GEN1491;
wire  _GEN1494 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1495 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1496 = io_x[30] ? _GEN1495 : _GEN1494;
wire  _GEN1497 = io_x[26] ? _GEN1496 : _GEN1493;
wire  _GEN1498 = io_x[22] ? _GEN1497 : _GEN1490;
wire  _GEN1499 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1500 = io_x[30] ? _GEN1499 : _GEN117;
wire  _GEN1501 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1502 = io_x[30] ? _GEN1501 : _GEN106;
wire  _GEN1503 = io_x[26] ? _GEN1502 : _GEN1500;
wire  _GEN1504 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1505 = io_x[30] ? _GEN1504 : _GEN117;
wire  _GEN1506 = io_x[26] ? _GEN1505 : _GEN119;
wire  _GEN1507 = io_x[22] ? _GEN1506 : _GEN1503;
wire  _GEN1508 = io_x[13] ? _GEN1507 : _GEN1498;
wire  _GEN1509 = io_x[33] ? _GEN1508 : _GEN1483;
wire  _GEN1510 = io_x[69] ? _GEN1509 : _GEN1461;
wire  _GEN1511 = io_x[71] ? _GEN1510 : _GEN1412;
wire  _GEN1512 = io_x[72] ? _GEN1511 : _GEN1315;
wire  _GEN1513 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1514 = io_x[30] ? _GEN117 : _GEN1513;
wire  _GEN1515 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1516 = io_x[26] ? _GEN1515 : _GEN1514;
wire  _GEN1517 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1518 = io_x[30] ? _GEN117 : _GEN1517;
wire  _GEN1519 = io_x[26] ? _GEN1518 : _GEN108;
wire  _GEN1520 = io_x[22] ? _GEN1519 : _GEN1516;
wire  _GEN1521 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1522 = io_x[30] ? _GEN1521 : _GEN117;
wire  _GEN1523 = io_x[26] ? _GEN1522 : _GEN119;
wire  _GEN1524 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1525 = io_x[30] ? _GEN117 : _GEN1524;
wire  _GEN1526 = io_x[26] ? _GEN1525 : _GEN108;
wire  _GEN1527 = io_x[22] ? _GEN1526 : _GEN1523;
wire  _GEN1528 = io_x[13] ? _GEN1527 : _GEN1520;
wire  _GEN1529 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1530 = io_x[30] ? _GEN117 : _GEN1529;
wire  _GEN1531 = io_x[26] ? _GEN1530 : _GEN119;
wire  _GEN1532 = io_x[22] ? _GEN314 : _GEN1531;
wire  _GEN1533 = io_x[26] ? _GEN108 : _GEN119;
wire  _GEN1534 = io_x[22] ? _GEN204 : _GEN1533;
wire  _GEN1535 = io_x[13] ? _GEN1534 : _GEN1532;
wire  _GEN1536 = io_x[33] ? _GEN1535 : _GEN1528;
wire  _GEN1537 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1538 = io_x[26] ? _GEN108 : _GEN1537;
wire  _GEN1539 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1540 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1541 = io_x[26] ? _GEN1540 : _GEN1539;
wire  _GEN1542 = io_x[22] ? _GEN1541 : _GEN1538;
wire  _GEN1543 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN1544 = io_x[22] ? _GEN1543 : _GEN314;
wire  _GEN1545 = io_x[13] ? _GEN1544 : _GEN1542;
wire  _GEN1546 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1547 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1548 = io_x[30] ? _GEN1547 : _GEN1546;
wire  _GEN1549 = io_x[26] ? _GEN1548 : _GEN119;
wire  _GEN1550 = io_x[22] ? _GEN314 : _GEN1549;
wire  _GEN1551 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1552 = io_x[30] ? _GEN1551 : _GEN117;
wire  _GEN1553 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1554 = io_x[30] ? _GEN1553 : _GEN117;
wire  _GEN1555 = io_x[26] ? _GEN1554 : _GEN1552;
wire  _GEN1556 = io_x[22] ? _GEN1555 : _GEN314;
wire  _GEN1557 = io_x[13] ? _GEN1556 : _GEN1550;
wire  _GEN1558 = io_x[33] ? _GEN1557 : _GEN1545;
wire  _GEN1559 = io_x[69] ? _GEN1558 : _GEN1536;
wire  _GEN1560 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1561 = io_x[30] ? _GEN117 : _GEN1560;
wire  _GEN1562 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1563 = io_x[30] ? _GEN117 : _GEN1562;
wire  _GEN1564 = io_x[26] ? _GEN1563 : _GEN1561;
wire  _GEN1565 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1566 = io_x[30] ? _GEN106 : _GEN1565;
wire  _GEN1567 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1568 = io_x[30] ? _GEN117 : _GEN1567;
wire  _GEN1569 = io_x[26] ? _GEN1568 : _GEN1566;
wire  _GEN1570 = io_x[22] ? _GEN1569 : _GEN1564;
wire  _GEN1571 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1572 = io_x[30] ? _GEN1571 : _GEN117;
wire  _GEN1573 = io_x[26] ? _GEN1572 : _GEN119;
wire  _GEN1574 = io_x[22] ? _GEN1573 : _GEN314;
wire  _GEN1575 = io_x[13] ? _GEN1574 : _GEN1570;
wire  _GEN1576 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1577 = io_x[26] ? _GEN119 : _GEN1576;
wire  _GEN1578 = io_x[22] ? _GEN1577 : _GEN204;
wire  _GEN1579 = io_x[13] ? _GEN1578 : _GEN563;
wire  _GEN1580 = io_x[33] ? _GEN1579 : _GEN1575;
wire  _GEN1581 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1582 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1583 = io_x[26] ? _GEN1582 : _GEN1581;
wire  _GEN1584 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1585 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1586 = io_x[30] ? _GEN1585 : _GEN1584;
wire  _GEN1587 = io_x[26] ? _GEN1586 : _GEN108;
wire  _GEN1588 = io_x[22] ? _GEN1587 : _GEN1583;
wire  _GEN1589 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1590 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1591 = io_x[26] ? _GEN1590 : _GEN1589;
wire  _GEN1592 = io_x[22] ? _GEN1591 : _GEN314;
wire  _GEN1593 = io_x[13] ? _GEN1592 : _GEN1588;
wire  _GEN1594 = io_x[22] ? _GEN314 : _GEN204;
wire  _GEN1595 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1596 = io_x[30] ? _GEN1595 : _GEN117;
wire  _GEN1597 = io_x[26] ? _GEN1596 : _GEN119;
wire  _GEN1598 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1599 = io_x[30] ? _GEN117 : _GEN1598;
wire  _GEN1600 = io_x[26] ? _GEN1599 : _GEN108;
wire  _GEN1601 = io_x[22] ? _GEN1600 : _GEN1597;
wire  _GEN1602 = io_x[13] ? _GEN1601 : _GEN1594;
wire  _GEN1603 = io_x[33] ? _GEN1602 : _GEN1593;
wire  _GEN1604 = io_x[69] ? _GEN1603 : _GEN1580;
wire  _GEN1605 = io_x[71] ? _GEN1604 : _GEN1559;
wire  _GEN1606 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1607 = io_x[30] ? _GEN117 : _GEN1606;
wire  _GEN1608 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1609 = io_x[30] ? _GEN1608 : _GEN117;
wire  _GEN1610 = io_x[26] ? _GEN1609 : _GEN1607;
wire  _GEN1611 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1612 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1613 = io_x[30] ? _GEN1612 : _GEN106;
wire  _GEN1614 = io_x[26] ? _GEN1613 : _GEN1611;
wire  _GEN1615 = io_x[22] ? _GEN1614 : _GEN1610;
wire  _GEN1616 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1617 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1618 = io_x[30] ? _GEN1617 : _GEN106;
wire  _GEN1619 = io_x[26] ? _GEN1618 : _GEN1616;
wire  _GEN1620 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1621 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1622 = io_x[30] ? _GEN1621 : _GEN117;
wire  _GEN1623 = io_x[26] ? _GEN1622 : _GEN1620;
wire  _GEN1624 = io_x[22] ? _GEN1623 : _GEN1619;
wire  _GEN1625 = io_x[13] ? _GEN1624 : _GEN1615;
wire  _GEN1626 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1627 = io_x[26] ? _GEN1626 : _GEN119;
wire  _GEN1628 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1629 = io_x[30] ? _GEN117 : _GEN1628;
wire  _GEN1630 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1631 = io_x[26] ? _GEN1630 : _GEN1629;
wire  _GEN1632 = io_x[22] ? _GEN1631 : _GEN1627;
wire  _GEN1633 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1634 = io_x[26] ? _GEN108 : _GEN1633;
wire  _GEN1635 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1636 = io_x[30] ? _GEN1635 : _GEN117;
wire  _GEN1637 = io_x[26] ? _GEN1636 : _GEN119;
wire  _GEN1638 = io_x[22] ? _GEN1637 : _GEN1634;
wire  _GEN1639 = io_x[13] ? _GEN1638 : _GEN1632;
wire  _GEN1640 = io_x[33] ? _GEN1639 : _GEN1625;
wire  _GEN1641 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1642 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1643 = io_x[30] ? _GEN1642 : _GEN1641;
wire  _GEN1644 = io_x[26] ? _GEN1643 : _GEN108;
wire  _GEN1645 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1646 = io_x[26] ? _GEN1645 : _GEN119;
wire  _GEN1647 = io_x[22] ? _GEN1646 : _GEN1644;
wire  _GEN1648 = io_x[13] ? _GEN523 : _GEN1647;
wire  _GEN1649 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1650 = io_x[26] ? _GEN1649 : _GEN119;
wire  _GEN1651 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1652 = io_x[30] ? _GEN1651 : _GEN117;
wire  _GEN1653 = io_x[26] ? _GEN108 : _GEN1652;
wire  _GEN1654 = io_x[22] ? _GEN1653 : _GEN1650;
wire  _GEN1655 = io_x[13] ? _GEN1654 : _GEN523;
wire  _GEN1656 = io_x[33] ? _GEN1655 : _GEN1648;
wire  _GEN1657 = io_x[69] ? _GEN1656 : _GEN1640;
wire  _GEN1658 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1659 = io_x[30] ? _GEN117 : _GEN1658;
wire  _GEN1660 = io_x[26] ? _GEN108 : _GEN1659;
wire  _GEN1661 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1662 = io_x[30] ? _GEN1661 : _GEN106;
wire  _GEN1663 = io_x[26] ? _GEN1662 : _GEN119;
wire  _GEN1664 = io_x[22] ? _GEN1663 : _GEN1660;
wire  _GEN1665 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN1666 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1667 = io_x[30] ? _GEN1666 : _GEN117;
wire  _GEN1668 = io_x[26] ? _GEN1667 : _GEN119;
wire  _GEN1669 = io_x[22] ? _GEN1668 : _GEN1665;
wire  _GEN1670 = io_x[13] ? _GEN1669 : _GEN1664;
wire  _GEN1671 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1672 = io_x[30] ? _GEN117 : _GEN1671;
wire  _GEN1673 = io_x[26] ? _GEN108 : _GEN1672;
wire  _GEN1674 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1675 = io_x[30] ? _GEN1674 : _GEN106;
wire  _GEN1676 = io_x[26] ? _GEN1675 : _GEN108;
wire  _GEN1677 = io_x[22] ? _GEN1676 : _GEN1673;
wire  _GEN1678 = io_x[22] ? _GEN204 : _GEN314;
wire  _GEN1679 = io_x[13] ? _GEN1678 : _GEN1677;
wire  _GEN1680 = io_x[33] ? _GEN1679 : _GEN1670;
wire  _GEN1681 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1682 = io_x[30] ? _GEN117 : _GEN1681;
wire  _GEN1683 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1684 = io_x[26] ? _GEN1683 : _GEN1682;
wire  _GEN1685 = io_x[22] ? _GEN314 : _GEN1684;
wire  _GEN1686 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1687 = io_x[26] ? _GEN1686 : _GEN119;
wire  _GEN1688 = io_x[22] ? _GEN1687 : _GEN314;
wire  _GEN1689 = io_x[13] ? _GEN1688 : _GEN1685;
wire  _GEN1690 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1691 = io_x[30] ? _GEN117 : _GEN1690;
wire  _GEN1692 = io_x[26] ? _GEN1691 : _GEN119;
wire  _GEN1693 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1694 = io_x[30] ? _GEN1693 : _GEN117;
wire  _GEN1695 = io_x[26] ? _GEN1694 : _GEN108;
wire  _GEN1696 = io_x[22] ? _GEN1695 : _GEN1692;
wire  _GEN1697 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1698 = io_x[30] ? _GEN1697 : _GEN117;
wire  _GEN1699 = io_x[26] ? _GEN1698 : _GEN119;
wire  _GEN1700 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1701 = io_x[30] ? _GEN1700 : _GEN106;
wire  _GEN1702 = io_x[26] ? _GEN1701 : _GEN108;
wire  _GEN1703 = io_x[22] ? _GEN1702 : _GEN1699;
wire  _GEN1704 = io_x[13] ? _GEN1703 : _GEN1696;
wire  _GEN1705 = io_x[33] ? _GEN1704 : _GEN1689;
wire  _GEN1706 = io_x[69] ? _GEN1705 : _GEN1680;
wire  _GEN1707 = io_x[71] ? _GEN1706 : _GEN1657;
wire  _GEN1708 = io_x[72] ? _GEN1707 : _GEN1605;
wire  _GEN1709 = io_x[48] ? _GEN1708 : _GEN1512;
wire  _GEN1710 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1711 = io_x[30] ? _GEN117 : _GEN1710;
wire  _GEN1712 = io_x[26] ? _GEN119 : _GEN1711;
wire  _GEN1713 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1714 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1715 = io_x[30] ? _GEN1714 : _GEN1713;
wire  _GEN1716 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1717 = io_x[30] ? _GEN1716 : _GEN106;
wire  _GEN1718 = io_x[26] ? _GEN1717 : _GEN1715;
wire  _GEN1719 = io_x[22] ? _GEN1718 : _GEN1712;
wire  _GEN1720 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1721 = io_x[30] ? _GEN1720 : _GEN117;
wire  _GEN1722 = io_x[26] ? _GEN1721 : _GEN119;
wire  _GEN1723 = io_x[22] ? _GEN1722 : _GEN314;
wire  _GEN1724 = io_x[13] ? _GEN1723 : _GEN1719;
wire  _GEN1725 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1726 = io_x[30] ? _GEN117 : _GEN1725;
wire  _GEN1727 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1728 = io_x[30] ? _GEN106 : _GEN1727;
wire  _GEN1729 = io_x[26] ? _GEN1728 : _GEN1726;
wire  _GEN1730 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1731 = io_x[30] ? _GEN106 : _GEN1730;
wire  _GEN1732 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1733 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1734 = io_x[30] ? _GEN1733 : _GEN1732;
wire  _GEN1735 = io_x[26] ? _GEN1734 : _GEN1731;
wire  _GEN1736 = io_x[22] ? _GEN1735 : _GEN1729;
wire  _GEN1737 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1738 = io_x[30] ? _GEN1737 : _GEN106;
wire  _GEN1739 = io_x[26] ? _GEN1738 : _GEN119;
wire  _GEN1740 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1741 = io_x[30] ? _GEN1740 : _GEN117;
wire  _GEN1742 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1743 = io_x[30] ? _GEN1742 : _GEN117;
wire  _GEN1744 = io_x[26] ? _GEN1743 : _GEN1741;
wire  _GEN1745 = io_x[22] ? _GEN1744 : _GEN1739;
wire  _GEN1746 = io_x[13] ? _GEN1745 : _GEN1736;
wire  _GEN1747 = io_x[33] ? _GEN1746 : _GEN1724;
wire  _GEN1748 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1749 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1750 = io_x[30] ? _GEN1749 : _GEN1748;
wire  _GEN1751 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1752 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1753 = io_x[30] ? _GEN1752 : _GEN1751;
wire  _GEN1754 = io_x[26] ? _GEN1753 : _GEN1750;
wire  _GEN1755 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1756 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1757 = io_x[30] ? _GEN1756 : _GEN1755;
wire  _GEN1758 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1759 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1760 = io_x[30] ? _GEN1759 : _GEN1758;
wire  _GEN1761 = io_x[26] ? _GEN1760 : _GEN1757;
wire  _GEN1762 = io_x[22] ? _GEN1761 : _GEN1754;
wire  _GEN1763 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1764 = io_x[30] ? _GEN1763 : _GEN117;
wire  _GEN1765 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1766 = io_x[30] ? _GEN1765 : _GEN117;
wire  _GEN1767 = io_x[26] ? _GEN1766 : _GEN1764;
wire  _GEN1768 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1769 = io_x[30] ? _GEN1768 : _GEN106;
wire  _GEN1770 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1771 = io_x[30] ? _GEN1770 : _GEN106;
wire  _GEN1772 = io_x[26] ? _GEN1771 : _GEN1769;
wire  _GEN1773 = io_x[22] ? _GEN1772 : _GEN1767;
wire  _GEN1774 = io_x[13] ? _GEN1773 : _GEN1762;
wire  _GEN1775 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1776 = io_x[30] ? _GEN117 : _GEN1775;
wire  _GEN1777 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1778 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1779 = io_x[30] ? _GEN1778 : _GEN1777;
wire  _GEN1780 = io_x[26] ? _GEN1779 : _GEN1776;
wire  _GEN1781 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1782 = io_x[30] ? _GEN1781 : _GEN106;
wire  _GEN1783 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1784 = io_x[30] ? _GEN106 : _GEN1783;
wire  _GEN1785 = io_x[26] ? _GEN1784 : _GEN1782;
wire  _GEN1786 = io_x[22] ? _GEN1785 : _GEN1780;
wire  _GEN1787 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1788 = io_x[30] ? _GEN1787 : _GEN106;
wire  _GEN1789 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1790 = io_x[30] ? _GEN1789 : _GEN106;
wire  _GEN1791 = io_x[26] ? _GEN1790 : _GEN1788;
wire  _GEN1792 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1793 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1794 = io_x[30] ? _GEN1793 : _GEN1792;
wire  _GEN1795 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1796 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1797 = io_x[30] ? _GEN1796 : _GEN1795;
wire  _GEN1798 = io_x[26] ? _GEN1797 : _GEN1794;
wire  _GEN1799 = io_x[22] ? _GEN1798 : _GEN1791;
wire  _GEN1800 = io_x[13] ? _GEN1799 : _GEN1786;
wire  _GEN1801 = io_x[33] ? _GEN1800 : _GEN1774;
wire  _GEN1802 = io_x[69] ? _GEN1801 : _GEN1747;
wire  _GEN1803 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1804 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1805 = io_x[30] ? _GEN1804 : _GEN1803;
wire  _GEN1806 = io_x[26] ? _GEN119 : _GEN1805;
wire  _GEN1807 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1808 = io_x[30] ? _GEN1807 : _GEN117;
wire  _GEN1809 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1810 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1811 = io_x[30] ? _GEN1810 : _GEN1809;
wire  _GEN1812 = io_x[26] ? _GEN1811 : _GEN1808;
wire  _GEN1813 = io_x[22] ? _GEN1812 : _GEN1806;
wire  _GEN1814 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1815 = io_x[30] ? _GEN1814 : _GEN117;
wire  _GEN1816 = io_x[26] ? _GEN119 : _GEN1815;
wire  _GEN1817 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1818 = io_x[30] ? _GEN1817 : _GEN117;
wire  _GEN1819 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1820 = io_x[30] ? _GEN1819 : _GEN117;
wire  _GEN1821 = io_x[26] ? _GEN1820 : _GEN1818;
wire  _GEN1822 = io_x[22] ? _GEN1821 : _GEN1816;
wire  _GEN1823 = io_x[13] ? _GEN1822 : _GEN1813;
wire  _GEN1824 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1825 = io_x[30] ? _GEN117 : _GEN1824;
wire  _GEN1826 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1827 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1828 = io_x[30] ? _GEN1827 : _GEN1826;
wire  _GEN1829 = io_x[26] ? _GEN1828 : _GEN1825;
wire  _GEN1830 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1831 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1832 = io_x[30] ? _GEN1831 : _GEN1830;
wire  _GEN1833 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1834 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1835 = io_x[30] ? _GEN1834 : _GEN1833;
wire  _GEN1836 = io_x[26] ? _GEN1835 : _GEN1832;
wire  _GEN1837 = io_x[22] ? _GEN1836 : _GEN1829;
wire  _GEN1838 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1839 = io_x[30] ? _GEN1838 : _GEN117;
wire  _GEN1840 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1841 = io_x[26] ? _GEN1840 : _GEN1839;
wire  _GEN1842 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1843 = io_x[30] ? _GEN1842 : _GEN117;
wire  _GEN1844 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1845 = io_x[30] ? _GEN1844 : _GEN117;
wire  _GEN1846 = io_x[26] ? _GEN1845 : _GEN1843;
wire  _GEN1847 = io_x[22] ? _GEN1846 : _GEN1841;
wire  _GEN1848 = io_x[13] ? _GEN1847 : _GEN1837;
wire  _GEN1849 = io_x[33] ? _GEN1848 : _GEN1823;
wire  _GEN1850 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1851 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1852 = io_x[30] ? _GEN1851 : _GEN117;
wire  _GEN1853 = io_x[26] ? _GEN1852 : _GEN1850;
wire  _GEN1854 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN1855 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1856 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1857 = io_x[30] ? _GEN1856 : _GEN1855;
wire  _GEN1858 = io_x[26] ? _GEN1857 : _GEN1854;
wire  _GEN1859 = io_x[22] ? _GEN1858 : _GEN1853;
wire  _GEN1860 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1861 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1862 = io_x[30] ? _GEN1861 : _GEN1860;
wire  _GEN1863 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1864 = io_x[30] ? _GEN1863 : _GEN106;
wire  _GEN1865 = io_x[26] ? _GEN1864 : _GEN1862;
wire  _GEN1866 = io_x[22] ? _GEN1865 : _GEN204;
wire  _GEN1867 = io_x[13] ? _GEN1866 : _GEN1859;
wire  _GEN1868 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1869 = io_x[30] ? _GEN117 : _GEN1868;
wire  _GEN1870 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1871 = io_x[30] ? _GEN1870 : _GEN117;
wire  _GEN1872 = io_x[26] ? _GEN1871 : _GEN1869;
wire  _GEN1873 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1874 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1875 = io_x[30] ? _GEN1874 : _GEN1873;
wire  _GEN1876 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1877 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1878 = io_x[30] ? _GEN1877 : _GEN1876;
wire  _GEN1879 = io_x[26] ? _GEN1878 : _GEN1875;
wire  _GEN1880 = io_x[22] ? _GEN1879 : _GEN1872;
wire  _GEN1881 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1882 = io_x[30] ? _GEN1881 : _GEN106;
wire  _GEN1883 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1884 = io_x[30] ? _GEN1883 : _GEN117;
wire  _GEN1885 = io_x[26] ? _GEN1884 : _GEN1882;
wire  _GEN1886 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1887 = io_x[30] ? _GEN106 : _GEN1886;
wire  _GEN1888 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1889 = io_x[30] ? _GEN1888 : _GEN117;
wire  _GEN1890 = io_x[26] ? _GEN1889 : _GEN1887;
wire  _GEN1891 = io_x[22] ? _GEN1890 : _GEN1885;
wire  _GEN1892 = io_x[13] ? _GEN1891 : _GEN1880;
wire  _GEN1893 = io_x[33] ? _GEN1892 : _GEN1867;
wire  _GEN1894 = io_x[69] ? _GEN1893 : _GEN1849;
wire  _GEN1895 = io_x[71] ? _GEN1894 : _GEN1802;
wire  _GEN1896 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1897 = io_x[30] ? _GEN117 : _GEN1896;
wire  _GEN1898 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1899 = io_x[30] ? _GEN117 : _GEN1898;
wire  _GEN1900 = io_x[26] ? _GEN1899 : _GEN1897;
wire  _GEN1901 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1902 = io_x[30] ? _GEN1901 : _GEN117;
wire  _GEN1903 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1904 = io_x[30] ? _GEN117 : _GEN1903;
wire  _GEN1905 = io_x[26] ? _GEN1904 : _GEN1902;
wire  _GEN1906 = io_x[22] ? _GEN1905 : _GEN1900;
wire  _GEN1907 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1908 = io_x[30] ? _GEN1907 : _GEN106;
wire  _GEN1909 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1910 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1911 = io_x[30] ? _GEN1910 : _GEN1909;
wire  _GEN1912 = io_x[26] ? _GEN1911 : _GEN1908;
wire  _GEN1913 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1914 = io_x[30] ? _GEN1913 : _GEN117;
wire  _GEN1915 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1916 = io_x[30] ? _GEN1915 : _GEN106;
wire  _GEN1917 = io_x[26] ? _GEN1916 : _GEN1914;
wire  _GEN1918 = io_x[22] ? _GEN1917 : _GEN1912;
wire  _GEN1919 = io_x[13] ? _GEN1918 : _GEN1906;
wire  _GEN1920 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1921 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1922 = io_x[30] ? _GEN1921 : _GEN1920;
wire  _GEN1923 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1924 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1925 = io_x[30] ? _GEN1924 : _GEN1923;
wire  _GEN1926 = io_x[26] ? _GEN1925 : _GEN1922;
wire  _GEN1927 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1928 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1929 = io_x[30] ? _GEN1928 : _GEN1927;
wire  _GEN1930 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1931 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1932 = io_x[30] ? _GEN1931 : _GEN1930;
wire  _GEN1933 = io_x[26] ? _GEN1932 : _GEN1929;
wire  _GEN1934 = io_x[22] ? _GEN1933 : _GEN1926;
wire  _GEN1935 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1936 = io_x[30] ? _GEN1935 : _GEN117;
wire  _GEN1937 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1938 = io_x[30] ? _GEN1937 : _GEN106;
wire  _GEN1939 = io_x[26] ? _GEN1938 : _GEN1936;
wire  _GEN1940 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1941 = io_x[30] ? _GEN1940 : _GEN106;
wire  _GEN1942 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1943 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1944 = io_x[30] ? _GEN1943 : _GEN1942;
wire  _GEN1945 = io_x[26] ? _GEN1944 : _GEN1941;
wire  _GEN1946 = io_x[22] ? _GEN1945 : _GEN1939;
wire  _GEN1947 = io_x[13] ? _GEN1946 : _GEN1934;
wire  _GEN1948 = io_x[33] ? _GEN1947 : _GEN1919;
wire  _GEN1949 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1950 = io_x[30] ? _GEN117 : _GEN1949;
wire  _GEN1951 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1952 = io_x[30] ? _GEN1951 : _GEN106;
wire  _GEN1953 = io_x[26] ? _GEN1952 : _GEN1950;
wire  _GEN1954 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1955 = io_x[30] ? _GEN1954 : _GEN117;
wire  _GEN1956 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1957 = io_x[30] ? _GEN1956 : _GEN117;
wire  _GEN1958 = io_x[26] ? _GEN1957 : _GEN1955;
wire  _GEN1959 = io_x[22] ? _GEN1958 : _GEN1953;
wire  _GEN1960 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1961 = io_x[30] ? _GEN1960 : _GEN117;
wire  _GEN1962 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1963 = io_x[30] ? _GEN1962 : _GEN117;
wire  _GEN1964 = io_x[26] ? _GEN1963 : _GEN1961;
wire  _GEN1965 = io_x[22] ? _GEN1964 : _GEN204;
wire  _GEN1966 = io_x[13] ? _GEN1965 : _GEN1959;
wire  _GEN1967 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1968 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1969 = io_x[30] ? _GEN1968 : _GEN1967;
wire  _GEN1970 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1971 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1972 = io_x[30] ? _GEN1971 : _GEN1970;
wire  _GEN1973 = io_x[26] ? _GEN1972 : _GEN1969;
wire  _GEN1974 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1975 = io_x[30] ? _GEN106 : _GEN1974;
wire  _GEN1976 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1977 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1978 = io_x[30] ? _GEN1977 : _GEN1976;
wire  _GEN1979 = io_x[26] ? _GEN1978 : _GEN1975;
wire  _GEN1980 = io_x[22] ? _GEN1979 : _GEN1973;
wire  _GEN1981 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1982 = io_x[30] ? _GEN1981 : _GEN117;
wire  _GEN1983 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1984 = io_x[30] ? _GEN1983 : _GEN117;
wire  _GEN1985 = io_x[26] ? _GEN1984 : _GEN1982;
wire  _GEN1986 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1987 = io_x[30] ? _GEN1986 : _GEN117;
wire  _GEN1988 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN1989 = io_x[30] ? _GEN1988 : _GEN117;
wire  _GEN1990 = io_x[26] ? _GEN1989 : _GEN1987;
wire  _GEN1991 = io_x[22] ? _GEN1990 : _GEN1985;
wire  _GEN1992 = io_x[13] ? _GEN1991 : _GEN1980;
wire  _GEN1993 = io_x[33] ? _GEN1992 : _GEN1966;
wire  _GEN1994 = io_x[69] ? _GEN1993 : _GEN1948;
wire  _GEN1995 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN1996 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN1997 = io_x[30] ? _GEN1996 : _GEN117;
wire  _GEN1998 = io_x[26] ? _GEN1997 : _GEN1995;
wire  _GEN1999 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2000 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2001 = io_x[30] ? _GEN2000 : _GEN1999;
wire  _GEN2002 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2003 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2004 = io_x[30] ? _GEN2003 : _GEN2002;
wire  _GEN2005 = io_x[26] ? _GEN2004 : _GEN2001;
wire  _GEN2006 = io_x[22] ? _GEN2005 : _GEN1998;
wire  _GEN2007 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2008 = io_x[30] ? _GEN117 : _GEN2007;
wire  _GEN2009 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2010 = io_x[30] ? _GEN2009 : _GEN117;
wire  _GEN2011 = io_x[26] ? _GEN2010 : _GEN2008;
wire  _GEN2012 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2013 = io_x[30] ? _GEN2012 : _GEN106;
wire  _GEN2014 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2015 = io_x[30] ? _GEN2014 : _GEN117;
wire  _GEN2016 = io_x[26] ? _GEN2015 : _GEN2013;
wire  _GEN2017 = io_x[22] ? _GEN2016 : _GEN2011;
wire  _GEN2018 = io_x[13] ? _GEN2017 : _GEN2006;
wire  _GEN2019 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2020 = io_x[30] ? _GEN117 : _GEN2019;
wire  _GEN2021 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2022 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2023 = io_x[30] ? _GEN2022 : _GEN2021;
wire  _GEN2024 = io_x[26] ? _GEN2023 : _GEN2020;
wire  _GEN2025 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2026 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2027 = io_x[30] ? _GEN2026 : _GEN2025;
wire  _GEN2028 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2029 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2030 = io_x[30] ? _GEN2029 : _GEN2028;
wire  _GEN2031 = io_x[26] ? _GEN2030 : _GEN2027;
wire  _GEN2032 = io_x[22] ? _GEN2031 : _GEN2024;
wire  _GEN2033 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2034 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2035 = io_x[30] ? _GEN2034 : _GEN2033;
wire  _GEN2036 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2037 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2038 = io_x[30] ? _GEN2037 : _GEN2036;
wire  _GEN2039 = io_x[26] ? _GEN2038 : _GEN2035;
wire  _GEN2040 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2041 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2042 = io_x[30] ? _GEN2041 : _GEN2040;
wire  _GEN2043 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2044 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2045 = io_x[30] ? _GEN2044 : _GEN2043;
wire  _GEN2046 = io_x[26] ? _GEN2045 : _GEN2042;
wire  _GEN2047 = io_x[22] ? _GEN2046 : _GEN2039;
wire  _GEN2048 = io_x[13] ? _GEN2047 : _GEN2032;
wire  _GEN2049 = io_x[33] ? _GEN2048 : _GEN2018;
wire  _GEN2050 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2051 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2052 = io_x[30] ? _GEN2051 : _GEN2050;
wire  _GEN2053 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2054 = io_x[30] ? _GEN117 : _GEN2053;
wire  _GEN2055 = io_x[26] ? _GEN2054 : _GEN2052;
wire  _GEN2056 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2057 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2058 = io_x[30] ? _GEN2057 : _GEN2056;
wire  _GEN2059 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2060 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2061 = io_x[30] ? _GEN2060 : _GEN2059;
wire  _GEN2062 = io_x[26] ? _GEN2061 : _GEN2058;
wire  _GEN2063 = io_x[22] ? _GEN2062 : _GEN2055;
wire  _GEN2064 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN2065 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2066 = io_x[30] ? _GEN2065 : _GEN117;
wire  _GEN2067 = io_x[26] ? _GEN2066 : _GEN2064;
wire  _GEN2068 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2069 = io_x[30] ? _GEN2068 : _GEN106;
wire  _GEN2070 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2071 = io_x[30] ? _GEN2070 : _GEN117;
wire  _GEN2072 = io_x[26] ? _GEN2071 : _GEN2069;
wire  _GEN2073 = io_x[22] ? _GEN2072 : _GEN2067;
wire  _GEN2074 = io_x[13] ? _GEN2073 : _GEN2063;
wire  _GEN2075 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2076 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2077 = io_x[30] ? _GEN2076 : _GEN2075;
wire  _GEN2078 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2079 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2080 = io_x[30] ? _GEN2079 : _GEN2078;
wire  _GEN2081 = io_x[26] ? _GEN2080 : _GEN2077;
wire  _GEN2082 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2083 = io_x[30] ? _GEN117 : _GEN2082;
wire  _GEN2084 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2085 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2086 = io_x[30] ? _GEN2085 : _GEN2084;
wire  _GEN2087 = io_x[26] ? _GEN2086 : _GEN2083;
wire  _GEN2088 = io_x[22] ? _GEN2087 : _GEN2081;
wire  _GEN2089 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2090 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2091 = io_x[30] ? _GEN2090 : _GEN2089;
wire  _GEN2092 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2093 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2094 = io_x[30] ? _GEN2093 : _GEN2092;
wire  _GEN2095 = io_x[26] ? _GEN2094 : _GEN2091;
wire  _GEN2096 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2097 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2098 = io_x[30] ? _GEN2097 : _GEN2096;
wire  _GEN2099 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2100 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2101 = io_x[30] ? _GEN2100 : _GEN2099;
wire  _GEN2102 = io_x[26] ? _GEN2101 : _GEN2098;
wire  _GEN2103 = io_x[22] ? _GEN2102 : _GEN2095;
wire  _GEN2104 = io_x[13] ? _GEN2103 : _GEN2088;
wire  _GEN2105 = io_x[33] ? _GEN2104 : _GEN2074;
wire  _GEN2106 = io_x[69] ? _GEN2105 : _GEN2049;
wire  _GEN2107 = io_x[71] ? _GEN2106 : _GEN1994;
wire  _GEN2108 = io_x[72] ? _GEN2107 : _GEN1895;
wire  _GEN2109 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN2110 = io_x[26] ? _GEN2109 : _GEN108;
wire  _GEN2111 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN2112 = io_x[26] ? _GEN2111 : _GEN119;
wire  _GEN2113 = io_x[22] ? _GEN2112 : _GEN2110;
wire  _GEN2114 = io_x[13] ? _GEN523 : _GEN2113;
wire  _GEN2115 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2116 = io_x[30] ? _GEN117 : _GEN2115;
wire  _GEN2117 = io_x[26] ? _GEN2116 : _GEN108;
wire  _GEN2118 = io_x[26] ? _GEN108 : _GEN119;
wire  _GEN2119 = io_x[22] ? _GEN2118 : _GEN2117;
wire  _GEN2120 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN2121 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2122 = io_x[30] ? _GEN2121 : _GEN117;
wire  _GEN2123 = io_x[26] ? _GEN2122 : _GEN2120;
wire  _GEN2124 = io_x[22] ? _GEN2123 : _GEN314;
wire  _GEN2125 = io_x[13] ? _GEN2124 : _GEN2119;
wire  _GEN2126 = io_x[33] ? _GEN2125 : _GEN2114;
wire  _GEN2127 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2128 = io_x[30] ? _GEN117 : _GEN2127;
wire  _GEN2129 = io_x[26] ? _GEN108 : _GEN2128;
wire  _GEN2130 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2131 = io_x[30] ? _GEN2130 : _GEN117;
wire  _GEN2132 = io_x[26] ? _GEN2131 : _GEN119;
wire  _GEN2133 = io_x[22] ? _GEN2132 : _GEN2129;
wire  _GEN2134 = io_x[22] ? _GEN204 : _GEN314;
wire  _GEN2135 = io_x[13] ? _GEN2134 : _GEN2133;
wire  _GEN2136 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2137 = io_x[30] ? _GEN106 : _GEN2136;
wire  _GEN2138 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2139 = io_x[30] ? _GEN106 : _GEN2138;
wire  _GEN2140 = io_x[26] ? _GEN2139 : _GEN2137;
wire  _GEN2141 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2142 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2143 = io_x[30] ? _GEN2142 : _GEN2141;
wire  _GEN2144 = io_x[26] ? _GEN2143 : _GEN119;
wire  _GEN2145 = io_x[22] ? _GEN2144 : _GEN2140;
wire  _GEN2146 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN2147 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN2148 = io_x[26] ? _GEN2147 : _GEN2146;
wire  _GEN2149 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2150 = io_x[30] ? _GEN2149 : _GEN106;
wire  _GEN2151 = io_x[26] ? _GEN2150 : _GEN108;
wire  _GEN2152 = io_x[22] ? _GEN2151 : _GEN2148;
wire  _GEN2153 = io_x[13] ? _GEN2152 : _GEN2145;
wire  _GEN2154 = io_x[33] ? _GEN2153 : _GEN2135;
wire  _GEN2155 = io_x[69] ? _GEN2154 : _GEN2126;
wire  _GEN2156 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2157 = io_x[30] ? _GEN117 : _GEN2156;
wire  _GEN2158 = io_x[26] ? _GEN2157 : _GEN119;
wire  _GEN2159 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2160 = io_x[30] ? _GEN117 : _GEN2159;
wire  _GEN2161 = io_x[26] ? _GEN119 : _GEN2160;
wire  _GEN2162 = io_x[22] ? _GEN2161 : _GEN2158;
wire  _GEN2163 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2164 = io_x[30] ? _GEN2163 : _GEN117;
wire  _GEN2165 = io_x[26] ? _GEN2164 : _GEN119;
wire  _GEN2166 = io_x[22] ? _GEN2165 : _GEN314;
wire  _GEN2167 = io_x[13] ? _GEN2166 : _GEN2162;
wire  _GEN2168 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2169 = io_x[30] ? _GEN117 : _GEN2168;
wire  _GEN2170 = io_x[26] ? _GEN119 : _GEN2169;
wire  _GEN2171 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2172 = io_x[30] ? _GEN117 : _GEN2171;
wire  _GEN2173 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN2174 = io_x[26] ? _GEN2173 : _GEN2172;
wire  _GEN2175 = io_x[22] ? _GEN2174 : _GEN2170;
wire  _GEN2176 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2177 = io_x[30] ? _GEN2176 : _GEN117;
wire  _GEN2178 = io_x[26] ? _GEN2177 : _GEN119;
wire  _GEN2179 = io_x[22] ? _GEN2178 : _GEN314;
wire  _GEN2180 = io_x[13] ? _GEN2179 : _GEN2175;
wire  _GEN2181 = io_x[33] ? _GEN2180 : _GEN2167;
wire  _GEN2182 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN2183 = io_x[26] ? _GEN108 : _GEN2182;
wire  _GEN2184 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2185 = io_x[30] ? _GEN2184 : _GEN117;
wire  _GEN2186 = io_x[26] ? _GEN2185 : _GEN119;
wire  _GEN2187 = io_x[22] ? _GEN2186 : _GEN2183;
wire  _GEN2188 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2189 = io_x[30] ? _GEN2188 : _GEN117;
wire  _GEN2190 = io_x[26] ? _GEN2189 : _GEN108;
wire  _GEN2191 = io_x[22] ? _GEN2190 : _GEN314;
wire  _GEN2192 = io_x[13] ? _GEN2191 : _GEN2187;
wire  _GEN2193 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN2194 = io_x[26] ? _GEN119 : _GEN2193;
wire  _GEN2195 = io_x[22] ? _GEN2194 : _GEN204;
wire  _GEN2196 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2197 = io_x[30] ? _GEN2196 : _GEN117;
wire  _GEN2198 = io_x[26] ? _GEN2197 : _GEN119;
wire  _GEN2199 = io_x[22] ? _GEN2198 : _GEN204;
wire  _GEN2200 = io_x[13] ? _GEN2199 : _GEN2195;
wire  _GEN2201 = io_x[33] ? _GEN2200 : _GEN2192;
wire  _GEN2202 = io_x[69] ? _GEN2201 : _GEN2181;
wire  _GEN2203 = io_x[71] ? _GEN2202 : _GEN2155;
wire  _GEN2204 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2205 = io_x[30] ? _GEN117 : _GEN2204;
wire  _GEN2206 = io_x[26] ? _GEN119 : _GEN2205;
wire  _GEN2207 = io_x[22] ? _GEN314 : _GEN2206;
wire  _GEN2208 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN2209 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2210 = io_x[30] ? _GEN117 : _GEN2209;
wire  _GEN2211 = io_x[26] ? _GEN2210 : _GEN2208;
wire  _GEN2212 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2213 = io_x[30] ? _GEN2212 : _GEN117;
wire  _GEN2214 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2215 = io_x[30] ? _GEN2214 : _GEN117;
wire  _GEN2216 = io_x[26] ? _GEN2215 : _GEN2213;
wire  _GEN2217 = io_x[22] ? _GEN2216 : _GEN2211;
wire  _GEN2218 = io_x[13] ? _GEN2217 : _GEN2207;
wire  _GEN2219 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2220 = io_x[30] ? _GEN2219 : _GEN117;
wire  _GEN2221 = io_x[26] ? _GEN2220 : _GEN119;
wire  _GEN2222 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2223 = io_x[30] ? _GEN117 : _GEN2222;
wire  _GEN2224 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2225 = io_x[30] ? _GEN117 : _GEN2224;
wire  _GEN2226 = io_x[26] ? _GEN2225 : _GEN2223;
wire  _GEN2227 = io_x[22] ? _GEN2226 : _GEN2221;
wire  _GEN2228 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2229 = io_x[30] ? _GEN2228 : _GEN117;
wire  _GEN2230 = io_x[26] ? _GEN2229 : _GEN108;
wire  _GEN2231 = io_x[22] ? _GEN2230 : _GEN314;
wire  _GEN2232 = io_x[13] ? _GEN2231 : _GEN2227;
wire  _GEN2233 = io_x[33] ? _GEN2232 : _GEN2218;
wire  _GEN2234 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2235 = io_x[30] ? _GEN117 : _GEN2234;
wire  _GEN2236 = io_x[26] ? _GEN119 : _GEN2235;
wire  _GEN2237 = io_x[26] ? _GEN119 : _GEN108;
wire  _GEN2238 = io_x[22] ? _GEN2237 : _GEN2236;
wire  _GEN2239 = io_x[26] ? _GEN108 : _GEN119;
wire  _GEN2240 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN2241 = io_x[26] ? _GEN2240 : _GEN119;
wire  _GEN2242 = io_x[22] ? _GEN2241 : _GEN2239;
wire  _GEN2243 = io_x[13] ? _GEN2242 : _GEN2238;
wire  _GEN2244 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2245 = io_x[30] ? _GEN117 : _GEN2244;
wire  _GEN2246 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN2247 = io_x[26] ? _GEN2246 : _GEN2245;
wire  _GEN2248 = io_x[30] ? _GEN117 : _GEN106;
wire  _GEN2249 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN2250 = io_x[26] ? _GEN2249 : _GEN2248;
wire  _GEN2251 = io_x[22] ? _GEN2250 : _GEN2247;
wire  _GEN2252 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN2253 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2254 = io_x[30] ? _GEN117 : _GEN2253;
wire  _GEN2255 = io_x[26] ? _GEN2254 : _GEN2252;
wire  _GEN2256 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN2257 = io_x[26] ? _GEN2256 : _GEN119;
wire  _GEN2258 = io_x[22] ? _GEN2257 : _GEN2255;
wire  _GEN2259 = io_x[13] ? _GEN2258 : _GEN2251;
wire  _GEN2260 = io_x[33] ? _GEN2259 : _GEN2243;
wire  _GEN2261 = io_x[69] ? _GEN2260 : _GEN2233;
wire  _GEN2262 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2263 = io_x[30] ? _GEN117 : _GEN2262;
wire  _GEN2264 = io_x[26] ? _GEN119 : _GEN2263;
wire  _GEN2265 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2266 = io_x[30] ? _GEN2265 : _GEN117;
wire  _GEN2267 = io_x[26] ? _GEN2266 : _GEN119;
wire  _GEN2268 = io_x[22] ? _GEN2267 : _GEN2264;
wire  _GEN2269 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2270 = io_x[30] ? _GEN2269 : _GEN117;
wire  _GEN2271 = io_x[26] ? _GEN2270 : _GEN108;
wire  _GEN2272 = io_x[22] ? _GEN2271 : _GEN314;
wire  _GEN2273 = io_x[13] ? _GEN2272 : _GEN2268;
wire  _GEN2274 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2275 = io_x[30] ? _GEN2274 : _GEN106;
wire  _GEN2276 = io_x[26] ? _GEN2275 : _GEN108;
wire  _GEN2277 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2278 = io_x[30] ? _GEN106 : _GEN2277;
wire  _GEN2279 = io_x[26] ? _GEN108 : _GEN2278;
wire  _GEN2280 = io_x[22] ? _GEN2279 : _GEN2276;
wire  _GEN2281 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2282 = io_x[30] ? _GEN2281 : _GEN117;
wire  _GEN2283 = io_x[26] ? _GEN2282 : _GEN108;
wire  _GEN2284 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2285 = io_x[30] ? _GEN2284 : _GEN117;
wire  _GEN2286 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2287 = io_x[30] ? _GEN2286 : _GEN117;
wire  _GEN2288 = io_x[26] ? _GEN2287 : _GEN2285;
wire  _GEN2289 = io_x[22] ? _GEN2288 : _GEN2283;
wire  _GEN2290 = io_x[13] ? _GEN2289 : _GEN2280;
wire  _GEN2291 = io_x[33] ? _GEN2290 : _GEN2273;
wire  _GEN2292 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2293 = io_x[30] ? _GEN117 : _GEN2292;
wire  _GEN2294 = io_x[26] ? _GEN119 : _GEN2293;
wire  _GEN2295 = io_x[22] ? _GEN2294 : _GEN314;
wire  _GEN2296 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2297 = io_x[30] ? _GEN117 : _GEN2296;
wire  _GEN2298 = io_x[26] ? _GEN119 : _GEN2297;
wire  _GEN2299 = io_x[22] ? _GEN314 : _GEN2298;
wire  _GEN2300 = io_x[13] ? _GEN2299 : _GEN2295;
wire  _GEN2301 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2302 = io_x[30] ? _GEN117 : _GEN2301;
wire  _GEN2303 = io_x[30] ? _GEN106 : _GEN117;
wire  _GEN2304 = io_x[26] ? _GEN2303 : _GEN2302;
wire  _GEN2305 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2306 = io_x[30] ? _GEN106 : _GEN2305;
wire  _GEN2307 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2308 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2309 = io_x[30] ? _GEN2308 : _GEN2307;
wire  _GEN2310 = io_x[26] ? _GEN2309 : _GEN2306;
wire  _GEN2311 = io_x[22] ? _GEN2310 : _GEN2304;
wire  _GEN2312 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2313 = io_x[30] ? _GEN2312 : _GEN117;
wire  _GEN2314 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2315 = io_x[30] ? _GEN2314 : _GEN117;
wire  _GEN2316 = io_x[26] ? _GEN2315 : _GEN2313;
wire  _GEN2317 = io_x[76] ? _GEN103 : _GEN104;
wire  _GEN2318 = io_x[76] ? _GEN104 : _GEN103;
wire  _GEN2319 = io_x[30] ? _GEN2318 : _GEN2317;
wire  _GEN2320 = io_x[26] ? _GEN2319 : _GEN119;
wire  _GEN2321 = io_x[22] ? _GEN2320 : _GEN2316;
wire  _GEN2322 = io_x[13] ? _GEN2321 : _GEN2311;
wire  _GEN2323 = io_x[33] ? _GEN2322 : _GEN2300;
wire  _GEN2324 = io_x[69] ? _GEN2323 : _GEN2291;
wire  _GEN2325 = io_x[71] ? _GEN2324 : _GEN2261;
wire  _GEN2326 = io_x[72] ? _GEN2325 : _GEN2203;
wire  _GEN2327 = io_x[48] ? _GEN2326 : _GEN2108;
wire  _GEN2328 = io_x[32] ? _GEN2327 : _GEN1709;
wire  _GEN2329 = io_x[18] ? _GEN2328 : _GEN1120;
assign io_y[17] = _GEN2329;
wire  _GEN2330 = 1'b0;
wire  _GEN2331 = 1'b1;
wire  _GEN2332 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2333 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2334 = io_x[29] ? _GEN2333 : _GEN2332;
wire  _GEN2335 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2336 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2337 = io_x[29] ? _GEN2336 : _GEN2335;
wire  _GEN2338 = io_x[17] ? _GEN2337 : _GEN2334;
wire  _GEN2339 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2340 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2341 = io_x[29] ? _GEN2340 : _GEN2339;
wire  _GEN2342 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2343 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2344 = io_x[29] ? _GEN2343 : _GEN2342;
wire  _GEN2345 = io_x[17] ? _GEN2344 : _GEN2341;
wire  _GEN2346 = io_x[21] ? _GEN2345 : _GEN2338;
wire  _GEN2347 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2348 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2349 = io_x[29] ? _GEN2348 : _GEN2347;
wire  _GEN2350 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2351 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2352 = io_x[29] ? _GEN2351 : _GEN2350;
wire  _GEN2353 = io_x[17] ? _GEN2352 : _GEN2349;
wire  _GEN2354 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2355 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2356 = io_x[29] ? _GEN2355 : _GEN2354;
wire  _GEN2357 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2358 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2359 = io_x[29] ? _GEN2358 : _GEN2357;
wire  _GEN2360 = io_x[17] ? _GEN2359 : _GEN2356;
wire  _GEN2361 = io_x[21] ? _GEN2360 : _GEN2353;
wire  _GEN2362 = io_x[9] ? _GEN2361 : _GEN2346;
wire  _GEN2363 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2364 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2365 = io_x[29] ? _GEN2364 : _GEN2363;
wire  _GEN2366 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2367 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2368 = io_x[29] ? _GEN2367 : _GEN2366;
wire  _GEN2369 = io_x[17] ? _GEN2368 : _GEN2365;
wire  _GEN2370 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2371 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2372 = io_x[29] ? _GEN2371 : _GEN2370;
wire  _GEN2373 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2374 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2375 = io_x[29] ? _GEN2374 : _GEN2373;
wire  _GEN2376 = io_x[17] ? _GEN2375 : _GEN2372;
wire  _GEN2377 = io_x[21] ? _GEN2376 : _GEN2369;
wire  _GEN2378 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2379 = 1'b0;
wire  _GEN2380 = io_x[29] ? _GEN2379 : _GEN2378;
wire  _GEN2381 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2382 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2383 = io_x[29] ? _GEN2382 : _GEN2381;
wire  _GEN2384 = io_x[17] ? _GEN2383 : _GEN2380;
wire  _GEN2385 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2386 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2387 = io_x[29] ? _GEN2386 : _GEN2385;
wire  _GEN2388 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2389 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2390 = io_x[29] ? _GEN2389 : _GEN2388;
wire  _GEN2391 = io_x[17] ? _GEN2390 : _GEN2387;
wire  _GEN2392 = io_x[21] ? _GEN2391 : _GEN2384;
wire  _GEN2393 = io_x[9] ? _GEN2392 : _GEN2377;
wire  _GEN2394 = io_x[1] ? _GEN2393 : _GEN2362;
wire  _GEN2395 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2396 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2397 = io_x[29] ? _GEN2396 : _GEN2395;
wire  _GEN2398 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2399 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2400 = io_x[29] ? _GEN2399 : _GEN2398;
wire  _GEN2401 = io_x[17] ? _GEN2400 : _GEN2397;
wire  _GEN2402 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2403 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2404 = io_x[29] ? _GEN2403 : _GEN2402;
wire  _GEN2405 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2406 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2407 = io_x[29] ? _GEN2406 : _GEN2405;
wire  _GEN2408 = io_x[17] ? _GEN2407 : _GEN2404;
wire  _GEN2409 = io_x[21] ? _GEN2408 : _GEN2401;
wire  _GEN2410 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2411 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2412 = io_x[29] ? _GEN2411 : _GEN2410;
wire  _GEN2413 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2414 = io_x[29] ? _GEN2413 : _GEN2379;
wire  _GEN2415 = io_x[17] ? _GEN2414 : _GEN2412;
wire  _GEN2416 = 1'b1;
wire  _GEN2417 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2418 = io_x[29] ? _GEN2417 : _GEN2416;
wire  _GEN2419 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2420 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2421 = io_x[29] ? _GEN2420 : _GEN2419;
wire  _GEN2422 = io_x[17] ? _GEN2421 : _GEN2418;
wire  _GEN2423 = io_x[21] ? _GEN2422 : _GEN2415;
wire  _GEN2424 = io_x[9] ? _GEN2423 : _GEN2409;
wire  _GEN2425 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2426 = io_x[29] ? _GEN2379 : _GEN2425;
wire  _GEN2427 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2428 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2429 = io_x[29] ? _GEN2428 : _GEN2427;
wire  _GEN2430 = io_x[17] ? _GEN2429 : _GEN2426;
wire  _GEN2431 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2432 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2433 = io_x[29] ? _GEN2432 : _GEN2431;
wire  _GEN2434 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2435 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2436 = io_x[29] ? _GEN2435 : _GEN2434;
wire  _GEN2437 = io_x[17] ? _GEN2436 : _GEN2433;
wire  _GEN2438 = io_x[21] ? _GEN2437 : _GEN2430;
wire  _GEN2439 = 1'b1;
wire  _GEN2440 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2441 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2442 = io_x[29] ? _GEN2441 : _GEN2440;
wire  _GEN2443 = io_x[17] ? _GEN2442 : _GEN2439;
wire  _GEN2444 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2445 = io_x[29] ? _GEN2444 : _GEN2416;
wire  _GEN2446 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2447 = io_x[29] ? _GEN2446 : _GEN2379;
wire  _GEN2448 = io_x[17] ? _GEN2447 : _GEN2445;
wire  _GEN2449 = io_x[21] ? _GEN2448 : _GEN2443;
wire  _GEN2450 = io_x[9] ? _GEN2449 : _GEN2438;
wire  _GEN2451 = io_x[1] ? _GEN2450 : _GEN2424;
wire  _GEN2452 = io_x[75] ? _GEN2451 : _GEN2394;
wire  _GEN2453 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2454 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2455 = io_x[29] ? _GEN2454 : _GEN2453;
wire  _GEN2456 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2457 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2458 = io_x[29] ? _GEN2457 : _GEN2456;
wire  _GEN2459 = io_x[17] ? _GEN2458 : _GEN2455;
wire  _GEN2460 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2461 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2462 = io_x[29] ? _GEN2461 : _GEN2460;
wire  _GEN2463 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2464 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2465 = io_x[29] ? _GEN2464 : _GEN2463;
wire  _GEN2466 = io_x[17] ? _GEN2465 : _GEN2462;
wire  _GEN2467 = io_x[21] ? _GEN2466 : _GEN2459;
wire  _GEN2468 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2469 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2470 = io_x[29] ? _GEN2469 : _GEN2468;
wire  _GEN2471 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2472 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2473 = io_x[29] ? _GEN2472 : _GEN2471;
wire  _GEN2474 = io_x[17] ? _GEN2473 : _GEN2470;
wire  _GEN2475 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2476 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2477 = io_x[29] ? _GEN2476 : _GEN2475;
wire  _GEN2478 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2479 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2480 = io_x[29] ? _GEN2479 : _GEN2478;
wire  _GEN2481 = io_x[17] ? _GEN2480 : _GEN2477;
wire  _GEN2482 = io_x[21] ? _GEN2481 : _GEN2474;
wire  _GEN2483 = io_x[9] ? _GEN2482 : _GEN2467;
wire  _GEN2484 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2485 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2486 = io_x[29] ? _GEN2485 : _GEN2484;
wire  _GEN2487 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2488 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2489 = io_x[29] ? _GEN2488 : _GEN2487;
wire  _GEN2490 = io_x[17] ? _GEN2489 : _GEN2486;
wire  _GEN2491 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2492 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2493 = io_x[29] ? _GEN2492 : _GEN2491;
wire  _GEN2494 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2495 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2496 = io_x[29] ? _GEN2495 : _GEN2494;
wire  _GEN2497 = io_x[17] ? _GEN2496 : _GEN2493;
wire  _GEN2498 = io_x[21] ? _GEN2497 : _GEN2490;
wire  _GEN2499 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2500 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2501 = io_x[29] ? _GEN2500 : _GEN2499;
wire  _GEN2502 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2503 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2504 = io_x[29] ? _GEN2503 : _GEN2502;
wire  _GEN2505 = io_x[17] ? _GEN2504 : _GEN2501;
wire  _GEN2506 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2507 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2508 = io_x[29] ? _GEN2507 : _GEN2506;
wire  _GEN2509 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2510 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2511 = io_x[29] ? _GEN2510 : _GEN2509;
wire  _GEN2512 = io_x[17] ? _GEN2511 : _GEN2508;
wire  _GEN2513 = io_x[21] ? _GEN2512 : _GEN2505;
wire  _GEN2514 = io_x[9] ? _GEN2513 : _GEN2498;
wire  _GEN2515 = io_x[1] ? _GEN2514 : _GEN2483;
wire  _GEN2516 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2517 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2518 = io_x[29] ? _GEN2517 : _GEN2516;
wire  _GEN2519 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2520 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2521 = io_x[29] ? _GEN2520 : _GEN2519;
wire  _GEN2522 = io_x[17] ? _GEN2521 : _GEN2518;
wire  _GEN2523 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2524 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2525 = io_x[29] ? _GEN2524 : _GEN2523;
wire  _GEN2526 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2527 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2528 = io_x[29] ? _GEN2527 : _GEN2526;
wire  _GEN2529 = io_x[17] ? _GEN2528 : _GEN2525;
wire  _GEN2530 = io_x[21] ? _GEN2529 : _GEN2522;
wire  _GEN2531 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2532 = io_x[29] ? _GEN2531 : _GEN2379;
wire  _GEN2533 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2534 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2535 = io_x[29] ? _GEN2534 : _GEN2533;
wire  _GEN2536 = io_x[17] ? _GEN2535 : _GEN2532;
wire  _GEN2537 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2538 = io_x[29] ? _GEN2537 : _GEN2416;
wire  _GEN2539 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2540 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2541 = io_x[29] ? _GEN2540 : _GEN2539;
wire  _GEN2542 = io_x[17] ? _GEN2541 : _GEN2538;
wire  _GEN2543 = io_x[21] ? _GEN2542 : _GEN2536;
wire  _GEN2544 = io_x[9] ? _GEN2543 : _GEN2530;
wire  _GEN2545 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2546 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2547 = io_x[29] ? _GEN2546 : _GEN2545;
wire  _GEN2548 = io_x[17] ? _GEN2547 : _GEN2439;
wire  _GEN2549 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2550 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2551 = io_x[29] ? _GEN2550 : _GEN2549;
wire  _GEN2552 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2553 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2554 = io_x[29] ? _GEN2553 : _GEN2552;
wire  _GEN2555 = io_x[17] ? _GEN2554 : _GEN2551;
wire  _GEN2556 = io_x[21] ? _GEN2555 : _GEN2548;
wire  _GEN2557 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2558 = io_x[29] ? _GEN2557 : _GEN2379;
wire  _GEN2559 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2560 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2561 = io_x[29] ? _GEN2560 : _GEN2559;
wire  _GEN2562 = io_x[17] ? _GEN2561 : _GEN2558;
wire  _GEN2563 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2564 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2565 = io_x[29] ? _GEN2564 : _GEN2563;
wire  _GEN2566 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2567 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2568 = io_x[29] ? _GEN2567 : _GEN2566;
wire  _GEN2569 = io_x[17] ? _GEN2568 : _GEN2565;
wire  _GEN2570 = io_x[21] ? _GEN2569 : _GEN2562;
wire  _GEN2571 = io_x[9] ? _GEN2570 : _GEN2556;
wire  _GEN2572 = io_x[1] ? _GEN2571 : _GEN2544;
wire  _GEN2573 = io_x[75] ? _GEN2572 : _GEN2515;
wire  _GEN2574 = io_x[32] ? _GEN2573 : _GEN2452;
wire  _GEN2575 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2576 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2577 = io_x[29] ? _GEN2576 : _GEN2575;
wire  _GEN2578 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2579 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2580 = io_x[29] ? _GEN2579 : _GEN2578;
wire  _GEN2581 = io_x[17] ? _GEN2580 : _GEN2577;
wire  _GEN2582 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2583 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2584 = io_x[29] ? _GEN2583 : _GEN2582;
wire  _GEN2585 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2586 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2587 = io_x[29] ? _GEN2586 : _GEN2585;
wire  _GEN2588 = io_x[17] ? _GEN2587 : _GEN2584;
wire  _GEN2589 = io_x[21] ? _GEN2588 : _GEN2581;
wire  _GEN2590 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2591 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2592 = io_x[29] ? _GEN2591 : _GEN2590;
wire  _GEN2593 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2594 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2595 = io_x[29] ? _GEN2594 : _GEN2593;
wire  _GEN2596 = io_x[17] ? _GEN2595 : _GEN2592;
wire  _GEN2597 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2598 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2599 = io_x[29] ? _GEN2598 : _GEN2597;
wire  _GEN2600 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2601 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2602 = io_x[29] ? _GEN2601 : _GEN2600;
wire  _GEN2603 = io_x[17] ? _GEN2602 : _GEN2599;
wire  _GEN2604 = io_x[21] ? _GEN2603 : _GEN2596;
wire  _GEN2605 = io_x[9] ? _GEN2604 : _GEN2589;
wire  _GEN2606 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2607 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2608 = io_x[29] ? _GEN2607 : _GEN2606;
wire  _GEN2609 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2610 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2611 = io_x[29] ? _GEN2610 : _GEN2609;
wire  _GEN2612 = io_x[17] ? _GEN2611 : _GEN2608;
wire  _GEN2613 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2614 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2615 = io_x[29] ? _GEN2614 : _GEN2613;
wire  _GEN2616 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2617 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2618 = io_x[29] ? _GEN2617 : _GEN2616;
wire  _GEN2619 = io_x[17] ? _GEN2618 : _GEN2615;
wire  _GEN2620 = io_x[21] ? _GEN2619 : _GEN2612;
wire  _GEN2621 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2622 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2623 = io_x[29] ? _GEN2622 : _GEN2621;
wire  _GEN2624 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2625 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2626 = io_x[29] ? _GEN2625 : _GEN2624;
wire  _GEN2627 = io_x[17] ? _GEN2626 : _GEN2623;
wire  _GEN2628 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2629 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2630 = io_x[29] ? _GEN2629 : _GEN2628;
wire  _GEN2631 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2632 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2633 = io_x[29] ? _GEN2632 : _GEN2631;
wire  _GEN2634 = io_x[17] ? _GEN2633 : _GEN2630;
wire  _GEN2635 = io_x[21] ? _GEN2634 : _GEN2627;
wire  _GEN2636 = io_x[9] ? _GEN2635 : _GEN2620;
wire  _GEN2637 = io_x[1] ? _GEN2636 : _GEN2605;
wire  _GEN2638 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2639 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2640 = io_x[29] ? _GEN2639 : _GEN2638;
wire  _GEN2641 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2642 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2643 = io_x[29] ? _GEN2642 : _GEN2641;
wire  _GEN2644 = io_x[17] ? _GEN2643 : _GEN2640;
wire  _GEN2645 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2646 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2647 = io_x[29] ? _GEN2646 : _GEN2645;
wire  _GEN2648 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2649 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2650 = io_x[29] ? _GEN2649 : _GEN2648;
wire  _GEN2651 = io_x[17] ? _GEN2650 : _GEN2647;
wire  _GEN2652 = io_x[21] ? _GEN2651 : _GEN2644;
wire  _GEN2653 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2654 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2655 = io_x[29] ? _GEN2654 : _GEN2653;
wire  _GEN2656 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2657 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2658 = io_x[29] ? _GEN2657 : _GEN2656;
wire  _GEN2659 = io_x[17] ? _GEN2658 : _GEN2655;
wire  _GEN2660 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2661 = io_x[29] ? _GEN2660 : _GEN2416;
wire  _GEN2662 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2663 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2664 = io_x[29] ? _GEN2663 : _GEN2662;
wire  _GEN2665 = io_x[17] ? _GEN2664 : _GEN2661;
wire  _GEN2666 = io_x[21] ? _GEN2665 : _GEN2659;
wire  _GEN2667 = io_x[9] ? _GEN2666 : _GEN2652;
wire  _GEN2668 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2669 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2670 = io_x[29] ? _GEN2669 : _GEN2668;
wire  _GEN2671 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2672 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2673 = io_x[29] ? _GEN2672 : _GEN2671;
wire  _GEN2674 = io_x[17] ? _GEN2673 : _GEN2670;
wire  _GEN2675 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2676 = io_x[29] ? _GEN2379 : _GEN2675;
wire  _GEN2677 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2678 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2679 = io_x[29] ? _GEN2678 : _GEN2677;
wire  _GEN2680 = io_x[17] ? _GEN2679 : _GEN2676;
wire  _GEN2681 = io_x[21] ? _GEN2680 : _GEN2674;
wire  _GEN2682 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2683 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2684 = io_x[29] ? _GEN2683 : _GEN2682;
wire  _GEN2685 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2686 = io_x[29] ? _GEN2379 : _GEN2685;
wire  _GEN2687 = io_x[17] ? _GEN2686 : _GEN2684;
wire  _GEN2688 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2689 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2690 = io_x[29] ? _GEN2689 : _GEN2688;
wire  _GEN2691 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2692 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2693 = io_x[29] ? _GEN2692 : _GEN2691;
wire  _GEN2694 = io_x[17] ? _GEN2693 : _GEN2690;
wire  _GEN2695 = io_x[21] ? _GEN2694 : _GEN2687;
wire  _GEN2696 = io_x[9] ? _GEN2695 : _GEN2681;
wire  _GEN2697 = io_x[1] ? _GEN2696 : _GEN2667;
wire  _GEN2698 = io_x[75] ? _GEN2697 : _GEN2637;
wire  _GEN2699 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2700 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2701 = io_x[29] ? _GEN2700 : _GEN2699;
wire  _GEN2702 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2703 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2704 = io_x[29] ? _GEN2703 : _GEN2702;
wire  _GEN2705 = io_x[17] ? _GEN2704 : _GEN2701;
wire  _GEN2706 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2707 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2708 = io_x[29] ? _GEN2707 : _GEN2706;
wire  _GEN2709 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2710 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2711 = io_x[29] ? _GEN2710 : _GEN2709;
wire  _GEN2712 = io_x[17] ? _GEN2711 : _GEN2708;
wire  _GEN2713 = io_x[21] ? _GEN2712 : _GEN2705;
wire  _GEN2714 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2715 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2716 = io_x[29] ? _GEN2715 : _GEN2714;
wire  _GEN2717 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2718 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2719 = io_x[29] ? _GEN2718 : _GEN2717;
wire  _GEN2720 = io_x[17] ? _GEN2719 : _GEN2716;
wire  _GEN2721 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2722 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2723 = io_x[29] ? _GEN2722 : _GEN2721;
wire  _GEN2724 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2725 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2726 = io_x[29] ? _GEN2725 : _GEN2724;
wire  _GEN2727 = io_x[17] ? _GEN2726 : _GEN2723;
wire  _GEN2728 = io_x[21] ? _GEN2727 : _GEN2720;
wire  _GEN2729 = io_x[9] ? _GEN2728 : _GEN2713;
wire  _GEN2730 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2731 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2732 = io_x[29] ? _GEN2731 : _GEN2730;
wire  _GEN2733 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2734 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2735 = io_x[29] ? _GEN2734 : _GEN2733;
wire  _GEN2736 = io_x[17] ? _GEN2735 : _GEN2732;
wire  _GEN2737 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2738 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2739 = io_x[29] ? _GEN2738 : _GEN2737;
wire  _GEN2740 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2741 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2742 = io_x[29] ? _GEN2741 : _GEN2740;
wire  _GEN2743 = io_x[17] ? _GEN2742 : _GEN2739;
wire  _GEN2744 = io_x[21] ? _GEN2743 : _GEN2736;
wire  _GEN2745 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2746 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2747 = io_x[29] ? _GEN2746 : _GEN2745;
wire  _GEN2748 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2749 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2750 = io_x[29] ? _GEN2749 : _GEN2748;
wire  _GEN2751 = io_x[17] ? _GEN2750 : _GEN2747;
wire  _GEN2752 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2753 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2754 = io_x[29] ? _GEN2753 : _GEN2752;
wire  _GEN2755 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2756 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2757 = io_x[29] ? _GEN2756 : _GEN2755;
wire  _GEN2758 = io_x[17] ? _GEN2757 : _GEN2754;
wire  _GEN2759 = io_x[21] ? _GEN2758 : _GEN2751;
wire  _GEN2760 = io_x[9] ? _GEN2759 : _GEN2744;
wire  _GEN2761 = io_x[1] ? _GEN2760 : _GEN2729;
wire  _GEN2762 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2763 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2764 = io_x[29] ? _GEN2763 : _GEN2762;
wire  _GEN2765 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2766 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2767 = io_x[29] ? _GEN2766 : _GEN2765;
wire  _GEN2768 = io_x[17] ? _GEN2767 : _GEN2764;
wire  _GEN2769 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2770 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2771 = io_x[29] ? _GEN2770 : _GEN2769;
wire  _GEN2772 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2773 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2774 = io_x[29] ? _GEN2773 : _GEN2772;
wire  _GEN2775 = io_x[17] ? _GEN2774 : _GEN2771;
wire  _GEN2776 = io_x[21] ? _GEN2775 : _GEN2768;
wire  _GEN2777 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2778 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2779 = io_x[29] ? _GEN2778 : _GEN2777;
wire  _GEN2780 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2781 = io_x[29] ? _GEN2780 : _GEN2416;
wire  _GEN2782 = io_x[17] ? _GEN2781 : _GEN2779;
wire  _GEN2783 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2784 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2785 = io_x[29] ? _GEN2784 : _GEN2783;
wire  _GEN2786 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2787 = io_x[29] ? _GEN2416 : _GEN2786;
wire  _GEN2788 = io_x[17] ? _GEN2787 : _GEN2785;
wire  _GEN2789 = io_x[21] ? _GEN2788 : _GEN2782;
wire  _GEN2790 = io_x[9] ? _GEN2789 : _GEN2776;
wire  _GEN2791 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2792 = io_x[29] ? _GEN2416 : _GEN2791;
wire  _GEN2793 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2794 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2795 = io_x[29] ? _GEN2794 : _GEN2793;
wire  _GEN2796 = io_x[17] ? _GEN2795 : _GEN2792;
wire  _GEN2797 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2798 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2799 = io_x[29] ? _GEN2798 : _GEN2797;
wire  _GEN2800 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2801 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2802 = io_x[29] ? _GEN2801 : _GEN2800;
wire  _GEN2803 = io_x[17] ? _GEN2802 : _GEN2799;
wire  _GEN2804 = io_x[21] ? _GEN2803 : _GEN2796;
wire  _GEN2805 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2806 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2807 = io_x[29] ? _GEN2806 : _GEN2805;
wire  _GEN2808 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2809 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2810 = io_x[29] ? _GEN2809 : _GEN2808;
wire  _GEN2811 = io_x[17] ? _GEN2810 : _GEN2807;
wire  _GEN2812 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2813 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2814 = io_x[29] ? _GEN2813 : _GEN2812;
wire  _GEN2815 = io_x[25] ? _GEN2330 : _GEN2331;
wire  _GEN2816 = io_x[25] ? _GEN2331 : _GEN2330;
wire  _GEN2817 = io_x[29] ? _GEN2816 : _GEN2815;
wire  _GEN2818 = io_x[17] ? _GEN2817 : _GEN2814;
wire  _GEN2819 = io_x[21] ? _GEN2818 : _GEN2811;
wire  _GEN2820 = io_x[9] ? _GEN2819 : _GEN2804;
wire  _GEN2821 = io_x[1] ? _GEN2820 : _GEN2790;
wire  _GEN2822 = io_x[75] ? _GEN2821 : _GEN2761;
wire  _GEN2823 = io_x[32] ? _GEN2822 : _GEN2698;
wire  _GEN2824 = io_x[37] ? _GEN2823 : _GEN2574;
assign io_y[16] = _GEN2824;
wire  _GEN2825 = 1'b0;
wire  _GEN2826 = 1'b1;
wire  _GEN2827 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2828 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2829 = io_x[28] ? _GEN2828 : _GEN2827;
wire  _GEN2830 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2831 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2832 = io_x[28] ? _GEN2831 : _GEN2830;
wire  _GEN2833 = io_x[74] ? _GEN2832 : _GEN2829;
wire  _GEN2834 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2835 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2836 = io_x[28] ? _GEN2835 : _GEN2834;
wire  _GEN2837 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2838 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2839 = io_x[28] ? _GEN2838 : _GEN2837;
wire  _GEN2840 = io_x[74] ? _GEN2839 : _GEN2836;
wire  _GEN2841 = io_x[24] ? _GEN2840 : _GEN2833;
wire  _GEN2842 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2843 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2844 = io_x[28] ? _GEN2843 : _GEN2842;
wire  _GEN2845 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2846 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2847 = io_x[28] ? _GEN2846 : _GEN2845;
wire  _GEN2848 = io_x[74] ? _GEN2847 : _GEN2844;
wire  _GEN2849 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2850 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2851 = io_x[28] ? _GEN2850 : _GEN2849;
wire  _GEN2852 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2853 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2854 = io_x[28] ? _GEN2853 : _GEN2852;
wire  _GEN2855 = io_x[74] ? _GEN2854 : _GEN2851;
wire  _GEN2856 = io_x[24] ? _GEN2855 : _GEN2848;
wire  _GEN2857 = io_x[80] ? _GEN2856 : _GEN2841;
wire  _GEN2858 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2859 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2860 = io_x[28] ? _GEN2859 : _GEN2858;
wire  _GEN2861 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2862 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2863 = io_x[28] ? _GEN2862 : _GEN2861;
wire  _GEN2864 = io_x[74] ? _GEN2863 : _GEN2860;
wire  _GEN2865 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2866 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2867 = io_x[28] ? _GEN2866 : _GEN2865;
wire  _GEN2868 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2869 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2870 = io_x[28] ? _GEN2869 : _GEN2868;
wire  _GEN2871 = io_x[74] ? _GEN2870 : _GEN2867;
wire  _GEN2872 = io_x[24] ? _GEN2871 : _GEN2864;
wire  _GEN2873 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2874 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2875 = io_x[28] ? _GEN2874 : _GEN2873;
wire  _GEN2876 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2877 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2878 = io_x[28] ? _GEN2877 : _GEN2876;
wire  _GEN2879 = io_x[74] ? _GEN2878 : _GEN2875;
wire  _GEN2880 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2881 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2882 = io_x[28] ? _GEN2881 : _GEN2880;
wire  _GEN2883 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2884 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2885 = io_x[28] ? _GEN2884 : _GEN2883;
wire  _GEN2886 = io_x[74] ? _GEN2885 : _GEN2882;
wire  _GEN2887 = io_x[24] ? _GEN2886 : _GEN2879;
wire  _GEN2888 = io_x[80] ? _GEN2887 : _GEN2872;
wire  _GEN2889 = io_x[20] ? _GEN2888 : _GEN2857;
wire  _GEN2890 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2891 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2892 = io_x[28] ? _GEN2891 : _GEN2890;
wire  _GEN2893 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2894 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2895 = io_x[28] ? _GEN2894 : _GEN2893;
wire  _GEN2896 = io_x[74] ? _GEN2895 : _GEN2892;
wire  _GEN2897 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2898 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2899 = io_x[28] ? _GEN2898 : _GEN2897;
wire  _GEN2900 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2901 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2902 = io_x[28] ? _GEN2901 : _GEN2900;
wire  _GEN2903 = io_x[74] ? _GEN2902 : _GEN2899;
wire  _GEN2904 = io_x[24] ? _GEN2903 : _GEN2896;
wire  _GEN2905 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2906 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2907 = io_x[28] ? _GEN2906 : _GEN2905;
wire  _GEN2908 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2909 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2910 = io_x[28] ? _GEN2909 : _GEN2908;
wire  _GEN2911 = io_x[74] ? _GEN2910 : _GEN2907;
wire  _GEN2912 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2913 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2914 = io_x[28] ? _GEN2913 : _GEN2912;
wire  _GEN2915 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2916 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2917 = io_x[28] ? _GEN2916 : _GEN2915;
wire  _GEN2918 = io_x[74] ? _GEN2917 : _GEN2914;
wire  _GEN2919 = io_x[24] ? _GEN2918 : _GEN2911;
wire  _GEN2920 = io_x[80] ? _GEN2919 : _GEN2904;
wire  _GEN2921 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2922 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2923 = io_x[28] ? _GEN2922 : _GEN2921;
wire  _GEN2924 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2925 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2926 = io_x[28] ? _GEN2925 : _GEN2924;
wire  _GEN2927 = io_x[74] ? _GEN2926 : _GEN2923;
wire  _GEN2928 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2929 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2930 = io_x[28] ? _GEN2929 : _GEN2928;
wire  _GEN2931 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2932 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2933 = io_x[28] ? _GEN2932 : _GEN2931;
wire  _GEN2934 = io_x[74] ? _GEN2933 : _GEN2930;
wire  _GEN2935 = io_x[24] ? _GEN2934 : _GEN2927;
wire  _GEN2936 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2937 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2938 = io_x[28] ? _GEN2937 : _GEN2936;
wire  _GEN2939 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2940 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2941 = io_x[28] ? _GEN2940 : _GEN2939;
wire  _GEN2942 = io_x[74] ? _GEN2941 : _GEN2938;
wire  _GEN2943 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2944 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2945 = io_x[28] ? _GEN2944 : _GEN2943;
wire  _GEN2946 = io_x[16] ? _GEN2825 : _GEN2826;
wire  _GEN2947 = io_x[16] ? _GEN2826 : _GEN2825;
wire  _GEN2948 = io_x[28] ? _GEN2947 : _GEN2946;
wire  _GEN2949 = io_x[74] ? _GEN2948 : _GEN2945;
wire  _GEN2950 = io_x[24] ? _GEN2949 : _GEN2942;
wire  _GEN2951 = io_x[80] ? _GEN2950 : _GEN2935;
wire  _GEN2952 = io_x[20] ? _GEN2951 : _GEN2920;
wire  _GEN2953 = io_x[18] ? _GEN2952 : _GEN2889;
assign io_y[15] = _GEN2953;
wire  _GEN2954 = 1'b0;
wire  _GEN2955 = 1'b1;
wire  _GEN2956 = io_x[73] ? _GEN2955 : _GEN2954;
wire  _GEN2957 = io_x[73] ? _GEN2955 : _GEN2954;
wire  _GEN2958 = io_x[45] ? _GEN2957 : _GEN2956;
wire  _GEN2959 = io_x[73] ? _GEN2955 : _GEN2954;
wire  _GEN2960 = io_x[73] ? _GEN2955 : _GEN2954;
wire  _GEN2961 = io_x[45] ? _GEN2960 : _GEN2959;
wire  _GEN2962 = io_x[15] ? _GEN2961 : _GEN2958;
assign io_y[14] = _GEN2962;
wire  _GEN2963 = 1'b0;
wire  _GEN2964 = 1'b1;
wire  _GEN2965 = io_x[72] ? _GEN2964 : _GEN2963;
wire  _GEN2966 = io_x[72] ? _GEN2964 : _GEN2963;
wire  _GEN2967 = io_x[40] ? _GEN2966 : _GEN2965;
wire  _GEN2968 = io_x[72] ? _GEN2964 : _GEN2963;
wire  _GEN2969 = io_x[72] ? _GEN2964 : _GEN2963;
wire  _GEN2970 = io_x[40] ? _GEN2969 : _GEN2968;
wire  _GEN2971 = io_x[81] ? _GEN2970 : _GEN2967;
wire  _GEN2972 = io_x[72] ? _GEN2964 : _GEN2963;
wire  _GEN2973 = io_x[72] ? _GEN2964 : _GEN2963;
wire  _GEN2974 = io_x[40] ? _GEN2973 : _GEN2972;
wire  _GEN2975 = io_x[72] ? _GEN2964 : _GEN2963;
wire  _GEN2976 = io_x[72] ? _GEN2964 : _GEN2963;
wire  _GEN2977 = io_x[40] ? _GEN2976 : _GEN2975;
wire  _GEN2978 = io_x[81] ? _GEN2977 : _GEN2974;
wire  _GEN2979 = io_x[19] ? _GEN2978 : _GEN2971;
assign io_y[13] = _GEN2979;
wire  _GEN2980 = 1'b0;
wire  _GEN2981 = 1'b1;
wire  _GEN2982 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN2983 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN2984 = io_x[38] ? _GEN2983 : _GEN2982;
wire  _GEN2985 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN2986 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN2987 = io_x[38] ? _GEN2986 : _GEN2985;
wire  _GEN2988 = io_x[41] ? _GEN2987 : _GEN2984;
wire  _GEN2989 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN2990 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN2991 = io_x[38] ? _GEN2990 : _GEN2989;
wire  _GEN2992 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN2993 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN2994 = io_x[38] ? _GEN2993 : _GEN2992;
wire  _GEN2995 = io_x[41] ? _GEN2994 : _GEN2991;
wire  _GEN2996 = io_x[43] ? _GEN2995 : _GEN2988;
wire  _GEN2997 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN2998 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN2999 = io_x[38] ? _GEN2998 : _GEN2997;
wire  _GEN3000 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN3001 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN3002 = io_x[38] ? _GEN3001 : _GEN3000;
wire  _GEN3003 = io_x[41] ? _GEN3002 : _GEN2999;
wire  _GEN3004 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN3005 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN3006 = io_x[38] ? _GEN3005 : _GEN3004;
wire  _GEN3007 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN3008 = io_x[71] ? _GEN2981 : _GEN2980;
wire  _GEN3009 = io_x[38] ? _GEN3008 : _GEN3007;
wire  _GEN3010 = io_x[41] ? _GEN3009 : _GEN3006;
wire  _GEN3011 = io_x[43] ? _GEN3010 : _GEN3003;
wire  _GEN3012 = io_x[75] ? _GEN3011 : _GEN2996;
assign io_y[12] = _GEN3012;
wire  _GEN3013 = 1'b0;
wire  _GEN3014 = 1'b1;
wire  _GEN3015 = io_x[70] ? _GEN3014 : _GEN3013;
wire  _GEN3016 = io_x[70] ? _GEN3014 : _GEN3013;
wire  _GEN3017 = io_x[37] ? _GEN3016 : _GEN3015;
assign io_y[11] = _GEN3017;
wire  _GEN3018 = 1'b0;
wire  _GEN3019 = 1'b1;
wire  _GEN3020 = io_x[69] ? _GEN3019 : _GEN3018;
wire  _GEN3021 = io_x[69] ? _GEN3019 : _GEN3018;
wire  _GEN3022 = io_x[43] ? _GEN3021 : _GEN3020;
assign io_y[10] = _GEN3022;
wire  _GEN3023 = 1'b0;
wire  _GEN3024 = 1'b1;
wire  _GEN3025 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3026 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3027 = io_x[11] ? _GEN3026 : _GEN3025;
wire  _GEN3028 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3029 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3030 = io_x[11] ? _GEN3029 : _GEN3028;
wire  _GEN3031 = io_x[15] ? _GEN3030 : _GEN3027;
wire  _GEN3032 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3033 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3034 = io_x[11] ? _GEN3033 : _GEN3032;
wire  _GEN3035 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3036 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3037 = io_x[11] ? _GEN3036 : _GEN3035;
wire  _GEN3038 = io_x[15] ? _GEN3037 : _GEN3034;
wire  _GEN3039 = io_x[3] ? _GEN3038 : _GEN3031;
wire  _GEN3040 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3041 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3042 = io_x[11] ? _GEN3041 : _GEN3040;
wire  _GEN3043 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3044 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3045 = io_x[11] ? _GEN3044 : _GEN3043;
wire  _GEN3046 = io_x[15] ? _GEN3045 : _GEN3042;
wire  _GEN3047 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3048 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3049 = io_x[11] ? _GEN3048 : _GEN3047;
wire  _GEN3050 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3051 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3052 = io_x[11] ? _GEN3051 : _GEN3050;
wire  _GEN3053 = io_x[15] ? _GEN3052 : _GEN3049;
wire  _GEN3054 = io_x[3] ? _GEN3053 : _GEN3046;
wire  _GEN3055 = io_x[9] ? _GEN3054 : _GEN3039;
wire  _GEN3056 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3057 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3058 = io_x[11] ? _GEN3057 : _GEN3056;
wire  _GEN3059 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3060 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3061 = io_x[11] ? _GEN3060 : _GEN3059;
wire  _GEN3062 = io_x[15] ? _GEN3061 : _GEN3058;
wire  _GEN3063 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3064 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3065 = io_x[11] ? _GEN3064 : _GEN3063;
wire  _GEN3066 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3067 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3068 = io_x[11] ? _GEN3067 : _GEN3066;
wire  _GEN3069 = io_x[15] ? _GEN3068 : _GEN3065;
wire  _GEN3070 = io_x[3] ? _GEN3069 : _GEN3062;
wire  _GEN3071 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3072 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3073 = io_x[11] ? _GEN3072 : _GEN3071;
wire  _GEN3074 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3075 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3076 = io_x[11] ? _GEN3075 : _GEN3074;
wire  _GEN3077 = io_x[15] ? _GEN3076 : _GEN3073;
wire  _GEN3078 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3079 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3080 = io_x[11] ? _GEN3079 : _GEN3078;
wire  _GEN3081 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3082 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3083 = io_x[11] ? _GEN3082 : _GEN3081;
wire  _GEN3084 = io_x[15] ? _GEN3083 : _GEN3080;
wire  _GEN3085 = io_x[3] ? _GEN3084 : _GEN3077;
wire  _GEN3086 = io_x[9] ? _GEN3085 : _GEN3070;
wire  _GEN3087 = io_x[48] ? _GEN3086 : _GEN3055;
wire  _GEN3088 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3089 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3090 = io_x[11] ? _GEN3089 : _GEN3088;
wire  _GEN3091 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3092 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3093 = io_x[11] ? _GEN3092 : _GEN3091;
wire  _GEN3094 = io_x[15] ? _GEN3093 : _GEN3090;
wire  _GEN3095 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3096 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3097 = io_x[11] ? _GEN3096 : _GEN3095;
wire  _GEN3098 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3099 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3100 = io_x[11] ? _GEN3099 : _GEN3098;
wire  _GEN3101 = io_x[15] ? _GEN3100 : _GEN3097;
wire  _GEN3102 = io_x[3] ? _GEN3101 : _GEN3094;
wire  _GEN3103 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3104 = 1'b1;
wire  _GEN3105 = io_x[11] ? _GEN3104 : _GEN3103;
wire  _GEN3106 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3107 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3108 = io_x[11] ? _GEN3107 : _GEN3106;
wire  _GEN3109 = io_x[15] ? _GEN3108 : _GEN3105;
wire  _GEN3110 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3111 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3112 = io_x[11] ? _GEN3111 : _GEN3110;
wire  _GEN3113 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3114 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3115 = io_x[11] ? _GEN3114 : _GEN3113;
wire  _GEN3116 = io_x[15] ? _GEN3115 : _GEN3112;
wire  _GEN3117 = io_x[3] ? _GEN3116 : _GEN3109;
wire  _GEN3118 = io_x[9] ? _GEN3117 : _GEN3102;
wire  _GEN3119 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3120 = io_x[11] ? _GEN3104 : _GEN3119;
wire  _GEN3121 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3122 = io_x[11] ? _GEN3121 : _GEN3104;
wire  _GEN3123 = io_x[15] ? _GEN3122 : _GEN3120;
wire  _GEN3124 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3125 = 1'b0;
wire  _GEN3126 = io_x[11] ? _GEN3125 : _GEN3124;
wire  _GEN3127 = io_x[11] ? _GEN3104 : _GEN3125;
wire  _GEN3128 = io_x[15] ? _GEN3127 : _GEN3126;
wire  _GEN3129 = io_x[3] ? _GEN3128 : _GEN3123;
wire  _GEN3130 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3131 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3132 = io_x[11] ? _GEN3131 : _GEN3130;
wire  _GEN3133 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3134 = io_x[11] ? _GEN3133 : _GEN3104;
wire  _GEN3135 = io_x[15] ? _GEN3134 : _GEN3132;
wire  _GEN3136 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3137 = io_x[11] ? _GEN3125 : _GEN3136;
wire  _GEN3138 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3139 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3140 = io_x[11] ? _GEN3139 : _GEN3138;
wire  _GEN3141 = io_x[15] ? _GEN3140 : _GEN3137;
wire  _GEN3142 = io_x[3] ? _GEN3141 : _GEN3135;
wire  _GEN3143 = io_x[9] ? _GEN3142 : _GEN3129;
wire  _GEN3144 = io_x[48] ? _GEN3143 : _GEN3118;
wire  _GEN3145 = io_x[45] ? _GEN3144 : _GEN3087;
wire  _GEN3146 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3147 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3148 = io_x[11] ? _GEN3147 : _GEN3146;
wire  _GEN3149 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3150 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3151 = io_x[11] ? _GEN3150 : _GEN3149;
wire  _GEN3152 = io_x[15] ? _GEN3151 : _GEN3148;
wire  _GEN3153 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3154 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3155 = io_x[11] ? _GEN3154 : _GEN3153;
wire  _GEN3156 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3157 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3158 = io_x[11] ? _GEN3157 : _GEN3156;
wire  _GEN3159 = io_x[15] ? _GEN3158 : _GEN3155;
wire  _GEN3160 = io_x[3] ? _GEN3159 : _GEN3152;
wire  _GEN3161 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3162 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3163 = io_x[11] ? _GEN3162 : _GEN3161;
wire  _GEN3164 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3165 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3166 = io_x[11] ? _GEN3165 : _GEN3164;
wire  _GEN3167 = io_x[15] ? _GEN3166 : _GEN3163;
wire  _GEN3168 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3169 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3170 = io_x[11] ? _GEN3169 : _GEN3168;
wire  _GEN3171 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3172 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3173 = io_x[11] ? _GEN3172 : _GEN3171;
wire  _GEN3174 = io_x[15] ? _GEN3173 : _GEN3170;
wire  _GEN3175 = io_x[3] ? _GEN3174 : _GEN3167;
wire  _GEN3176 = io_x[9] ? _GEN3175 : _GEN3160;
wire  _GEN3177 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3178 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3179 = io_x[11] ? _GEN3178 : _GEN3177;
wire  _GEN3180 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3181 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3182 = io_x[11] ? _GEN3181 : _GEN3180;
wire  _GEN3183 = io_x[15] ? _GEN3182 : _GEN3179;
wire  _GEN3184 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3185 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3186 = io_x[11] ? _GEN3185 : _GEN3184;
wire  _GEN3187 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3188 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3189 = io_x[11] ? _GEN3188 : _GEN3187;
wire  _GEN3190 = io_x[15] ? _GEN3189 : _GEN3186;
wire  _GEN3191 = io_x[3] ? _GEN3190 : _GEN3183;
wire  _GEN3192 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3193 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3194 = io_x[11] ? _GEN3193 : _GEN3192;
wire  _GEN3195 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3196 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3197 = io_x[11] ? _GEN3196 : _GEN3195;
wire  _GEN3198 = io_x[15] ? _GEN3197 : _GEN3194;
wire  _GEN3199 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3200 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3201 = io_x[11] ? _GEN3200 : _GEN3199;
wire  _GEN3202 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3203 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3204 = io_x[11] ? _GEN3203 : _GEN3202;
wire  _GEN3205 = io_x[15] ? _GEN3204 : _GEN3201;
wire  _GEN3206 = io_x[3] ? _GEN3205 : _GEN3198;
wire  _GEN3207 = io_x[9] ? _GEN3206 : _GEN3191;
wire  _GEN3208 = io_x[48] ? _GEN3207 : _GEN3176;
wire  _GEN3209 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3210 = io_x[11] ? _GEN3104 : _GEN3209;
wire  _GEN3211 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3212 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3213 = io_x[11] ? _GEN3212 : _GEN3211;
wire  _GEN3214 = io_x[15] ? _GEN3213 : _GEN3210;
wire  _GEN3215 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3216 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3217 = io_x[11] ? _GEN3216 : _GEN3215;
wire  _GEN3218 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3219 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3220 = io_x[11] ? _GEN3219 : _GEN3218;
wire  _GEN3221 = io_x[15] ? _GEN3220 : _GEN3217;
wire  _GEN3222 = io_x[3] ? _GEN3221 : _GEN3214;
wire  _GEN3223 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3224 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3225 = io_x[11] ? _GEN3224 : _GEN3223;
wire  _GEN3226 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3227 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3228 = io_x[11] ? _GEN3227 : _GEN3226;
wire  _GEN3229 = io_x[15] ? _GEN3228 : _GEN3225;
wire  _GEN3230 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3231 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3232 = io_x[11] ? _GEN3231 : _GEN3230;
wire  _GEN3233 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3234 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3235 = io_x[11] ? _GEN3234 : _GEN3233;
wire  _GEN3236 = io_x[15] ? _GEN3235 : _GEN3232;
wire  _GEN3237 = io_x[3] ? _GEN3236 : _GEN3229;
wire  _GEN3238 = io_x[9] ? _GEN3237 : _GEN3222;
wire  _GEN3239 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3240 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3241 = io_x[11] ? _GEN3240 : _GEN3239;
wire  _GEN3242 = 1'b0;
wire  _GEN3243 = io_x[15] ? _GEN3242 : _GEN3241;
wire  _GEN3244 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3245 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3246 = io_x[11] ? _GEN3245 : _GEN3244;
wire  _GEN3247 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3248 = io_x[11] ? _GEN3104 : _GEN3247;
wire  _GEN3249 = io_x[15] ? _GEN3248 : _GEN3246;
wire  _GEN3250 = io_x[3] ? _GEN3249 : _GEN3243;
wire  _GEN3251 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3252 = io_x[11] ? _GEN3251 : _GEN3104;
wire  _GEN3253 = io_x[11] ? _GEN3125 : _GEN3104;
wire  _GEN3254 = io_x[15] ? _GEN3253 : _GEN3252;
wire  _GEN3255 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3256 = io_x[11] ? _GEN3255 : _GEN3104;
wire  _GEN3257 = io_x[7] ? _GEN3023 : _GEN3024;
wire  _GEN3258 = io_x[7] ? _GEN3024 : _GEN3023;
wire  _GEN3259 = io_x[11] ? _GEN3258 : _GEN3257;
wire  _GEN3260 = io_x[15] ? _GEN3259 : _GEN3256;
wire  _GEN3261 = io_x[3] ? _GEN3260 : _GEN3254;
wire  _GEN3262 = io_x[9] ? _GEN3261 : _GEN3250;
wire  _GEN3263 = io_x[48] ? _GEN3262 : _GEN3238;
wire  _GEN3264 = io_x[45] ? _GEN3263 : _GEN3208;
wire  _GEN3265 = io_x[34] ? _GEN3264 : _GEN3145;
assign io_y[9] = _GEN3265;
wire  _GEN3266 = 1'b0;
wire  _GEN3267 = 1'b1;
wire  _GEN3268 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3269 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3270 = io_x[14] ? _GEN3269 : _GEN3268;
wire  _GEN3271 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3272 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3273 = io_x[14] ? _GEN3272 : _GEN3271;
wire  _GEN3274 = io_x[2] ? _GEN3273 : _GEN3270;
wire  _GEN3275 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3276 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3277 = io_x[14] ? _GEN3276 : _GEN3275;
wire  _GEN3278 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3279 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3280 = io_x[14] ? _GEN3279 : _GEN3278;
wire  _GEN3281 = io_x[2] ? _GEN3280 : _GEN3277;
wire  _GEN3282 = io_x[6] ? _GEN3281 : _GEN3274;
wire  _GEN3283 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3284 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3285 = io_x[14] ? _GEN3284 : _GEN3283;
wire  _GEN3286 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3287 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3288 = io_x[14] ? _GEN3287 : _GEN3286;
wire  _GEN3289 = io_x[2] ? _GEN3288 : _GEN3285;
wire  _GEN3290 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3291 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3292 = io_x[14] ? _GEN3291 : _GEN3290;
wire  _GEN3293 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3294 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3295 = io_x[14] ? _GEN3294 : _GEN3293;
wire  _GEN3296 = io_x[2] ? _GEN3295 : _GEN3292;
wire  _GEN3297 = io_x[6] ? _GEN3296 : _GEN3289;
wire  _GEN3298 = io_x[44] ? _GEN3297 : _GEN3282;
wire  _GEN3299 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3300 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3301 = io_x[14] ? _GEN3300 : _GEN3299;
wire  _GEN3302 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3303 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3304 = io_x[14] ? _GEN3303 : _GEN3302;
wire  _GEN3305 = io_x[2] ? _GEN3304 : _GEN3301;
wire  _GEN3306 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3307 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3308 = io_x[14] ? _GEN3307 : _GEN3306;
wire  _GEN3309 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3310 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3311 = io_x[14] ? _GEN3310 : _GEN3309;
wire  _GEN3312 = io_x[2] ? _GEN3311 : _GEN3308;
wire  _GEN3313 = io_x[6] ? _GEN3312 : _GEN3305;
wire  _GEN3314 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3315 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3316 = io_x[14] ? _GEN3315 : _GEN3314;
wire  _GEN3317 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3318 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3319 = io_x[14] ? _GEN3318 : _GEN3317;
wire  _GEN3320 = io_x[2] ? _GEN3319 : _GEN3316;
wire  _GEN3321 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3322 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3323 = io_x[14] ? _GEN3322 : _GEN3321;
wire  _GEN3324 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3325 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3326 = io_x[14] ? _GEN3325 : _GEN3324;
wire  _GEN3327 = io_x[2] ? _GEN3326 : _GEN3323;
wire  _GEN3328 = io_x[6] ? _GEN3327 : _GEN3320;
wire  _GEN3329 = io_x[44] ? _GEN3328 : _GEN3313;
wire  _GEN3330 = io_x[75] ? _GEN3329 : _GEN3298;
wire  _GEN3331 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3332 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3333 = io_x[14] ? _GEN3332 : _GEN3331;
wire  _GEN3334 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3335 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3336 = io_x[14] ? _GEN3335 : _GEN3334;
wire  _GEN3337 = io_x[2] ? _GEN3336 : _GEN3333;
wire  _GEN3338 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3339 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3340 = io_x[14] ? _GEN3339 : _GEN3338;
wire  _GEN3341 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3342 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3343 = io_x[14] ? _GEN3342 : _GEN3341;
wire  _GEN3344 = io_x[2] ? _GEN3343 : _GEN3340;
wire  _GEN3345 = io_x[6] ? _GEN3344 : _GEN3337;
wire  _GEN3346 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3347 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3348 = io_x[14] ? _GEN3347 : _GEN3346;
wire  _GEN3349 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3350 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3351 = io_x[14] ? _GEN3350 : _GEN3349;
wire  _GEN3352 = io_x[2] ? _GEN3351 : _GEN3348;
wire  _GEN3353 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3354 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3355 = io_x[14] ? _GEN3354 : _GEN3353;
wire  _GEN3356 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3357 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3358 = io_x[14] ? _GEN3357 : _GEN3356;
wire  _GEN3359 = io_x[2] ? _GEN3358 : _GEN3355;
wire  _GEN3360 = io_x[6] ? _GEN3359 : _GEN3352;
wire  _GEN3361 = io_x[44] ? _GEN3360 : _GEN3345;
wire  _GEN3362 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3363 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3364 = io_x[14] ? _GEN3363 : _GEN3362;
wire  _GEN3365 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3366 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3367 = io_x[14] ? _GEN3366 : _GEN3365;
wire  _GEN3368 = io_x[2] ? _GEN3367 : _GEN3364;
wire  _GEN3369 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3370 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3371 = io_x[14] ? _GEN3370 : _GEN3369;
wire  _GEN3372 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3373 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3374 = io_x[14] ? _GEN3373 : _GEN3372;
wire  _GEN3375 = io_x[2] ? _GEN3374 : _GEN3371;
wire  _GEN3376 = io_x[6] ? _GEN3375 : _GEN3368;
wire  _GEN3377 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3378 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3379 = io_x[14] ? _GEN3378 : _GEN3377;
wire  _GEN3380 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3381 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3382 = io_x[14] ? _GEN3381 : _GEN3380;
wire  _GEN3383 = io_x[2] ? _GEN3382 : _GEN3379;
wire  _GEN3384 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3385 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3386 = io_x[14] ? _GEN3385 : _GEN3384;
wire  _GEN3387 = io_x[10] ? _GEN3266 : _GEN3267;
wire  _GEN3388 = io_x[10] ? _GEN3267 : _GEN3266;
wire  _GEN3389 = io_x[14] ? _GEN3388 : _GEN3387;
wire  _GEN3390 = io_x[2] ? _GEN3389 : _GEN3386;
wire  _GEN3391 = io_x[6] ? _GEN3390 : _GEN3383;
wire  _GEN3392 = io_x[44] ? _GEN3391 : _GEN3376;
wire  _GEN3393 = io_x[75] ? _GEN3392 : _GEN3361;
wire  _GEN3394 = io_x[19] ? _GEN3393 : _GEN3330;
assign io_y[8] = _GEN3394;
wire  _GEN3395 = 1'b0;
wire  _GEN3396 = 1'b1;
wire  _GEN3397 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3398 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3399 = io_x[13] ? _GEN3398 : _GEN3397;
wire  _GEN3400 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3401 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3402 = io_x[13] ? _GEN3401 : _GEN3400;
wire  _GEN3403 = io_x[1] ? _GEN3402 : _GEN3399;
wire  _GEN3404 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3405 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3406 = io_x[13] ? _GEN3405 : _GEN3404;
wire  _GEN3407 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3408 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3409 = io_x[13] ? _GEN3408 : _GEN3407;
wire  _GEN3410 = io_x[1] ? _GEN3409 : _GEN3406;
wire  _GEN3411 = io_x[5] ? _GEN3410 : _GEN3403;
wire  _GEN3412 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3413 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3414 = io_x[13] ? _GEN3413 : _GEN3412;
wire  _GEN3415 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3416 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3417 = io_x[13] ? _GEN3416 : _GEN3415;
wire  _GEN3418 = io_x[1] ? _GEN3417 : _GEN3414;
wire  _GEN3419 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3420 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3421 = io_x[13] ? _GEN3420 : _GEN3419;
wire  _GEN3422 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3423 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3424 = io_x[13] ? _GEN3423 : _GEN3422;
wire  _GEN3425 = io_x[1] ? _GEN3424 : _GEN3421;
wire  _GEN3426 = io_x[5] ? _GEN3425 : _GEN3418;
wire  _GEN3427 = io_x[2] ? _GEN3426 : _GEN3411;
wire  _GEN3428 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3429 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3430 = io_x[13] ? _GEN3429 : _GEN3428;
wire  _GEN3431 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3432 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3433 = io_x[13] ? _GEN3432 : _GEN3431;
wire  _GEN3434 = io_x[1] ? _GEN3433 : _GEN3430;
wire  _GEN3435 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3436 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3437 = io_x[13] ? _GEN3436 : _GEN3435;
wire  _GEN3438 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3439 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3440 = io_x[13] ? _GEN3439 : _GEN3438;
wire  _GEN3441 = io_x[1] ? _GEN3440 : _GEN3437;
wire  _GEN3442 = io_x[5] ? _GEN3441 : _GEN3434;
wire  _GEN3443 = 1'b1;
wire  _GEN3444 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3445 = io_x[13] ? _GEN3444 : _GEN3443;
wire  _GEN3446 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3447 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3448 = io_x[13] ? _GEN3447 : _GEN3446;
wire  _GEN3449 = io_x[1] ? _GEN3448 : _GEN3445;
wire  _GEN3450 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3451 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3452 = io_x[13] ? _GEN3451 : _GEN3450;
wire  _GEN3453 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3454 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3455 = io_x[13] ? _GEN3454 : _GEN3453;
wire  _GEN3456 = io_x[1] ? _GEN3455 : _GEN3452;
wire  _GEN3457 = io_x[5] ? _GEN3456 : _GEN3449;
wire  _GEN3458 = io_x[2] ? _GEN3457 : _GEN3442;
wire  _GEN3459 = io_x[43] ? _GEN3458 : _GEN3427;
wire  _GEN3460 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3461 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3462 = io_x[13] ? _GEN3461 : _GEN3460;
wire  _GEN3463 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3464 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3465 = io_x[13] ? _GEN3464 : _GEN3463;
wire  _GEN3466 = io_x[1] ? _GEN3465 : _GEN3462;
wire  _GEN3467 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3468 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3469 = io_x[13] ? _GEN3468 : _GEN3467;
wire  _GEN3470 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3471 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3472 = io_x[13] ? _GEN3471 : _GEN3470;
wire  _GEN3473 = io_x[1] ? _GEN3472 : _GEN3469;
wire  _GEN3474 = io_x[5] ? _GEN3473 : _GEN3466;
wire  _GEN3475 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3476 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3477 = io_x[13] ? _GEN3476 : _GEN3475;
wire  _GEN3478 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3479 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3480 = io_x[13] ? _GEN3479 : _GEN3478;
wire  _GEN3481 = io_x[1] ? _GEN3480 : _GEN3477;
wire  _GEN3482 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3483 = io_x[13] ? _GEN3443 : _GEN3482;
wire  _GEN3484 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3485 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3486 = io_x[13] ? _GEN3485 : _GEN3484;
wire  _GEN3487 = io_x[1] ? _GEN3486 : _GEN3483;
wire  _GEN3488 = io_x[5] ? _GEN3487 : _GEN3481;
wire  _GEN3489 = io_x[2] ? _GEN3488 : _GEN3474;
wire  _GEN3490 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3491 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3492 = io_x[13] ? _GEN3491 : _GEN3490;
wire  _GEN3493 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3494 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3495 = io_x[13] ? _GEN3494 : _GEN3493;
wire  _GEN3496 = io_x[1] ? _GEN3495 : _GEN3492;
wire  _GEN3497 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3498 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3499 = io_x[13] ? _GEN3498 : _GEN3497;
wire  _GEN3500 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3501 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3502 = io_x[13] ? _GEN3501 : _GEN3500;
wire  _GEN3503 = io_x[1] ? _GEN3502 : _GEN3499;
wire  _GEN3504 = io_x[5] ? _GEN3503 : _GEN3496;
wire  _GEN3505 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3506 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3507 = io_x[13] ? _GEN3506 : _GEN3505;
wire  _GEN3508 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3509 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3510 = io_x[13] ? _GEN3509 : _GEN3508;
wire  _GEN3511 = io_x[1] ? _GEN3510 : _GEN3507;
wire  _GEN3512 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3513 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3514 = io_x[13] ? _GEN3513 : _GEN3512;
wire  _GEN3515 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3516 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3517 = io_x[13] ? _GEN3516 : _GEN3515;
wire  _GEN3518 = io_x[1] ? _GEN3517 : _GEN3514;
wire  _GEN3519 = io_x[5] ? _GEN3518 : _GEN3511;
wire  _GEN3520 = io_x[2] ? _GEN3519 : _GEN3504;
wire  _GEN3521 = io_x[43] ? _GEN3520 : _GEN3489;
wire  _GEN3522 = io_x[48] ? _GEN3521 : _GEN3459;
wire  _GEN3523 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3524 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3525 = io_x[13] ? _GEN3524 : _GEN3523;
wire  _GEN3526 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3527 = 1'b0;
wire  _GEN3528 = io_x[13] ? _GEN3527 : _GEN3526;
wire  _GEN3529 = io_x[1] ? _GEN3528 : _GEN3525;
wire  _GEN3530 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3531 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3532 = io_x[13] ? _GEN3531 : _GEN3530;
wire  _GEN3533 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3534 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3535 = io_x[13] ? _GEN3534 : _GEN3533;
wire  _GEN3536 = io_x[1] ? _GEN3535 : _GEN3532;
wire  _GEN3537 = io_x[5] ? _GEN3536 : _GEN3529;
wire  _GEN3538 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3539 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3540 = io_x[13] ? _GEN3539 : _GEN3538;
wire  _GEN3541 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3542 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3543 = io_x[13] ? _GEN3542 : _GEN3541;
wire  _GEN3544 = io_x[1] ? _GEN3543 : _GEN3540;
wire  _GEN3545 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3546 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3547 = io_x[13] ? _GEN3546 : _GEN3545;
wire  _GEN3548 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3549 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3550 = io_x[13] ? _GEN3549 : _GEN3548;
wire  _GEN3551 = io_x[1] ? _GEN3550 : _GEN3547;
wire  _GEN3552 = io_x[5] ? _GEN3551 : _GEN3544;
wire  _GEN3553 = io_x[2] ? _GEN3552 : _GEN3537;
wire  _GEN3554 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3555 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3556 = io_x[13] ? _GEN3555 : _GEN3554;
wire  _GEN3557 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3558 = io_x[13] ? _GEN3557 : _GEN3527;
wire  _GEN3559 = io_x[1] ? _GEN3558 : _GEN3556;
wire  _GEN3560 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3561 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3562 = io_x[13] ? _GEN3561 : _GEN3560;
wire  _GEN3563 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3564 = io_x[13] ? _GEN3443 : _GEN3563;
wire  _GEN3565 = io_x[1] ? _GEN3564 : _GEN3562;
wire  _GEN3566 = io_x[5] ? _GEN3565 : _GEN3559;
wire  _GEN3567 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3568 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3569 = io_x[13] ? _GEN3568 : _GEN3567;
wire  _GEN3570 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3571 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3572 = io_x[13] ? _GEN3571 : _GEN3570;
wire  _GEN3573 = io_x[1] ? _GEN3572 : _GEN3569;
wire  _GEN3574 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3575 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3576 = io_x[13] ? _GEN3575 : _GEN3574;
wire  _GEN3577 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3578 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3579 = io_x[13] ? _GEN3578 : _GEN3577;
wire  _GEN3580 = io_x[1] ? _GEN3579 : _GEN3576;
wire  _GEN3581 = io_x[5] ? _GEN3580 : _GEN3573;
wire  _GEN3582 = io_x[2] ? _GEN3581 : _GEN3566;
wire  _GEN3583 = io_x[43] ? _GEN3582 : _GEN3553;
wire  _GEN3584 = 1'b1;
wire  _GEN3585 = 1'b1;
wire  _GEN3586 = 1'b0;
wire  _GEN3587 = 1'b1;
wire  _GEN3588 = io_x[1] ? _GEN3587 : _GEN3586;
wire  _GEN3589 = io_x[5] ? _GEN3588 : _GEN3585;
wire  _GEN3590 = io_x[2] ? _GEN3589 : _GEN3584;
wire  _GEN3591 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3592 = io_x[13] ? _GEN3443 : _GEN3591;
wire  _GEN3593 = io_x[1] ? _GEN3592 : _GEN3587;
wire  _GEN3594 = io_x[1] ? _GEN3586 : _GEN3587;
wire  _GEN3595 = io_x[5] ? _GEN3594 : _GEN3593;
wire  _GEN3596 = io_x[2] ? _GEN3595 : _GEN3584;
wire  _GEN3597 = io_x[43] ? _GEN3596 : _GEN3590;
wire  _GEN3598 = io_x[48] ? _GEN3597 : _GEN3583;
wire  _GEN3599 = io_x[81] ? _GEN3598 : _GEN3522;
wire  _GEN3600 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3601 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3602 = io_x[13] ? _GEN3601 : _GEN3600;
wire  _GEN3603 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3604 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3605 = io_x[13] ? _GEN3604 : _GEN3603;
wire  _GEN3606 = io_x[1] ? _GEN3605 : _GEN3602;
wire  _GEN3607 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3608 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3609 = io_x[13] ? _GEN3608 : _GEN3607;
wire  _GEN3610 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3611 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3612 = io_x[13] ? _GEN3611 : _GEN3610;
wire  _GEN3613 = io_x[1] ? _GEN3612 : _GEN3609;
wire  _GEN3614 = io_x[5] ? _GEN3613 : _GEN3606;
wire  _GEN3615 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3616 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3617 = io_x[13] ? _GEN3616 : _GEN3615;
wire  _GEN3618 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3619 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3620 = io_x[13] ? _GEN3619 : _GEN3618;
wire  _GEN3621 = io_x[1] ? _GEN3620 : _GEN3617;
wire  _GEN3622 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3623 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3624 = io_x[13] ? _GEN3623 : _GEN3622;
wire  _GEN3625 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3626 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3627 = io_x[13] ? _GEN3626 : _GEN3625;
wire  _GEN3628 = io_x[1] ? _GEN3627 : _GEN3624;
wire  _GEN3629 = io_x[5] ? _GEN3628 : _GEN3621;
wire  _GEN3630 = io_x[2] ? _GEN3629 : _GEN3614;
wire  _GEN3631 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3632 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3633 = io_x[13] ? _GEN3632 : _GEN3631;
wire  _GEN3634 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3635 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3636 = io_x[13] ? _GEN3635 : _GEN3634;
wire  _GEN3637 = io_x[1] ? _GEN3636 : _GEN3633;
wire  _GEN3638 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3639 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3640 = io_x[13] ? _GEN3639 : _GEN3638;
wire  _GEN3641 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3642 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3643 = io_x[13] ? _GEN3642 : _GEN3641;
wire  _GEN3644 = io_x[1] ? _GEN3643 : _GEN3640;
wire  _GEN3645 = io_x[5] ? _GEN3644 : _GEN3637;
wire  _GEN3646 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3647 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3648 = io_x[13] ? _GEN3647 : _GEN3646;
wire  _GEN3649 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3650 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3651 = io_x[13] ? _GEN3650 : _GEN3649;
wire  _GEN3652 = io_x[1] ? _GEN3651 : _GEN3648;
wire  _GEN3653 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3654 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3655 = io_x[13] ? _GEN3654 : _GEN3653;
wire  _GEN3656 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3657 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3658 = io_x[13] ? _GEN3657 : _GEN3656;
wire  _GEN3659 = io_x[1] ? _GEN3658 : _GEN3655;
wire  _GEN3660 = io_x[5] ? _GEN3659 : _GEN3652;
wire  _GEN3661 = io_x[2] ? _GEN3660 : _GEN3645;
wire  _GEN3662 = io_x[43] ? _GEN3661 : _GEN3630;
wire  _GEN3663 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3664 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3665 = io_x[13] ? _GEN3664 : _GEN3663;
wire  _GEN3666 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3667 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3668 = io_x[13] ? _GEN3667 : _GEN3666;
wire  _GEN3669 = io_x[1] ? _GEN3668 : _GEN3665;
wire  _GEN3670 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3671 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3672 = io_x[13] ? _GEN3671 : _GEN3670;
wire  _GEN3673 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3674 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3675 = io_x[13] ? _GEN3674 : _GEN3673;
wire  _GEN3676 = io_x[1] ? _GEN3675 : _GEN3672;
wire  _GEN3677 = io_x[5] ? _GEN3676 : _GEN3669;
wire  _GEN3678 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3679 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3680 = io_x[13] ? _GEN3679 : _GEN3678;
wire  _GEN3681 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3682 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3683 = io_x[13] ? _GEN3682 : _GEN3681;
wire  _GEN3684 = io_x[1] ? _GEN3683 : _GEN3680;
wire  _GEN3685 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3686 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3687 = io_x[13] ? _GEN3686 : _GEN3685;
wire  _GEN3688 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3689 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3690 = io_x[13] ? _GEN3689 : _GEN3688;
wire  _GEN3691 = io_x[1] ? _GEN3690 : _GEN3687;
wire  _GEN3692 = io_x[5] ? _GEN3691 : _GEN3684;
wire  _GEN3693 = io_x[2] ? _GEN3692 : _GEN3677;
wire  _GEN3694 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3695 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3696 = io_x[13] ? _GEN3695 : _GEN3694;
wire  _GEN3697 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3698 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3699 = io_x[13] ? _GEN3698 : _GEN3697;
wire  _GEN3700 = io_x[1] ? _GEN3699 : _GEN3696;
wire  _GEN3701 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3702 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3703 = io_x[13] ? _GEN3702 : _GEN3701;
wire  _GEN3704 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3705 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3706 = io_x[13] ? _GEN3705 : _GEN3704;
wire  _GEN3707 = io_x[1] ? _GEN3706 : _GEN3703;
wire  _GEN3708 = io_x[5] ? _GEN3707 : _GEN3700;
wire  _GEN3709 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3710 = io_x[13] ? _GEN3443 : _GEN3709;
wire  _GEN3711 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3712 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3713 = io_x[13] ? _GEN3712 : _GEN3711;
wire  _GEN3714 = io_x[1] ? _GEN3713 : _GEN3710;
wire  _GEN3715 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3716 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3717 = io_x[13] ? _GEN3716 : _GEN3715;
wire  _GEN3718 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3719 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3720 = io_x[13] ? _GEN3719 : _GEN3718;
wire  _GEN3721 = io_x[1] ? _GEN3720 : _GEN3717;
wire  _GEN3722 = io_x[5] ? _GEN3721 : _GEN3714;
wire  _GEN3723 = io_x[2] ? _GEN3722 : _GEN3708;
wire  _GEN3724 = io_x[43] ? _GEN3723 : _GEN3693;
wire  _GEN3725 = io_x[48] ? _GEN3724 : _GEN3662;
wire  _GEN3726 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3727 = io_x[13] ? _GEN3443 : _GEN3726;
wire  _GEN3728 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3729 = io_x[13] ? _GEN3443 : _GEN3728;
wire  _GEN3730 = io_x[1] ? _GEN3729 : _GEN3727;
wire  _GEN3731 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3732 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3733 = io_x[13] ? _GEN3732 : _GEN3731;
wire  _GEN3734 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3735 = io_x[13] ? _GEN3527 : _GEN3734;
wire  _GEN3736 = io_x[1] ? _GEN3735 : _GEN3733;
wire  _GEN3737 = io_x[5] ? _GEN3736 : _GEN3730;
wire  _GEN3738 = io_x[13] ? _GEN3443 : _GEN3527;
wire  _GEN3739 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3740 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3741 = io_x[13] ? _GEN3740 : _GEN3739;
wire  _GEN3742 = io_x[1] ? _GEN3741 : _GEN3738;
wire  _GEN3743 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3744 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3745 = io_x[13] ? _GEN3744 : _GEN3743;
wire  _GEN3746 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3747 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3748 = io_x[13] ? _GEN3747 : _GEN3746;
wire  _GEN3749 = io_x[1] ? _GEN3748 : _GEN3745;
wire  _GEN3750 = io_x[5] ? _GEN3749 : _GEN3742;
wire  _GEN3751 = io_x[2] ? _GEN3750 : _GEN3737;
wire  _GEN3752 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3753 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3754 = io_x[13] ? _GEN3753 : _GEN3752;
wire  _GEN3755 = io_x[1] ? _GEN3586 : _GEN3754;
wire  _GEN3756 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3757 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3758 = io_x[13] ? _GEN3757 : _GEN3756;
wire  _GEN3759 = io_x[1] ? _GEN3758 : _GEN3586;
wire  _GEN3760 = io_x[5] ? _GEN3759 : _GEN3755;
wire  _GEN3761 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3762 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3763 = io_x[13] ? _GEN3762 : _GEN3761;
wire  _GEN3764 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3765 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3766 = io_x[13] ? _GEN3765 : _GEN3764;
wire  _GEN3767 = io_x[1] ? _GEN3766 : _GEN3763;
wire  _GEN3768 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3769 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3770 = io_x[13] ? _GEN3769 : _GEN3768;
wire  _GEN3771 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3772 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3773 = io_x[13] ? _GEN3772 : _GEN3771;
wire  _GEN3774 = io_x[1] ? _GEN3773 : _GEN3770;
wire  _GEN3775 = io_x[5] ? _GEN3774 : _GEN3767;
wire  _GEN3776 = io_x[2] ? _GEN3775 : _GEN3760;
wire  _GEN3777 = io_x[43] ? _GEN3776 : _GEN3751;
wire  _GEN3778 = 1'b0;
wire  _GEN3779 = io_x[2] ? _GEN3584 : _GEN3778;
wire  _GEN3780 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3781 = io_x[13] ? _GEN3780 : _GEN3443;
wire  _GEN3782 = io_x[1] ? _GEN3587 : _GEN3781;
wire  _GEN3783 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3784 = io_x[13] ? _GEN3783 : _GEN3443;
wire  _GEN3785 = io_x[13] ? _GEN3443 : _GEN3527;
wire  _GEN3786 = io_x[1] ? _GEN3785 : _GEN3784;
wire  _GEN3787 = io_x[5] ? _GEN3786 : _GEN3782;
wire  _GEN3788 = io_x[13] ? _GEN3527 : _GEN3443;
wire  _GEN3789 = io_x[1] ? _GEN3788 : _GEN3587;
wire  _GEN3790 = io_x[13] ? _GEN3527 : _GEN3443;
wire  _GEN3791 = io_x[9] ? _GEN3395 : _GEN3396;
wire  _GEN3792 = io_x[9] ? _GEN3396 : _GEN3395;
wire  _GEN3793 = io_x[13] ? _GEN3792 : _GEN3791;
wire  _GEN3794 = io_x[1] ? _GEN3793 : _GEN3790;
wire  _GEN3795 = io_x[5] ? _GEN3794 : _GEN3789;
wire  _GEN3796 = io_x[2] ? _GEN3795 : _GEN3787;
wire  _GEN3797 = io_x[43] ? _GEN3796 : _GEN3779;
wire  _GEN3798 = io_x[48] ? _GEN3797 : _GEN3777;
wire  _GEN3799 = io_x[81] ? _GEN3798 : _GEN3725;
wire  _GEN3800 = io_x[40] ? _GEN3799 : _GEN3599;
assign io_y[7] = _GEN3800;
wire  _GEN3801 = 1'b0;
wire  _GEN3802 = 1'b1;
wire  _GEN3803 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3804 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3805 = io_x[4] ? _GEN3804 : _GEN3803;
wire  _GEN3806 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3807 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3808 = io_x[4] ? _GEN3807 : _GEN3806;
wire  _GEN3809 = io_x[12] ? _GEN3808 : _GEN3805;
wire  _GEN3810 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3811 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3812 = io_x[4] ? _GEN3811 : _GEN3810;
wire  _GEN3813 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3814 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3815 = io_x[4] ? _GEN3814 : _GEN3813;
wire  _GEN3816 = io_x[12] ? _GEN3815 : _GEN3812;
wire  _GEN3817 = io_x[0] ? _GEN3816 : _GEN3809;
wire  _GEN3818 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3819 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3820 = io_x[4] ? _GEN3819 : _GEN3818;
wire  _GEN3821 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3822 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3823 = io_x[4] ? _GEN3822 : _GEN3821;
wire  _GEN3824 = io_x[12] ? _GEN3823 : _GEN3820;
wire  _GEN3825 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3826 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3827 = io_x[4] ? _GEN3826 : _GEN3825;
wire  _GEN3828 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3829 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3830 = io_x[4] ? _GEN3829 : _GEN3828;
wire  _GEN3831 = io_x[12] ? _GEN3830 : _GEN3827;
wire  _GEN3832 = io_x[0] ? _GEN3831 : _GEN3824;
wire  _GEN3833 = io_x[42] ? _GEN3832 : _GEN3817;
wire  _GEN3834 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3835 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3836 = io_x[4] ? _GEN3835 : _GEN3834;
wire  _GEN3837 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3838 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3839 = io_x[4] ? _GEN3838 : _GEN3837;
wire  _GEN3840 = io_x[12] ? _GEN3839 : _GEN3836;
wire  _GEN3841 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3842 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3843 = io_x[4] ? _GEN3842 : _GEN3841;
wire  _GEN3844 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3845 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3846 = io_x[4] ? _GEN3845 : _GEN3844;
wire  _GEN3847 = io_x[12] ? _GEN3846 : _GEN3843;
wire  _GEN3848 = io_x[0] ? _GEN3847 : _GEN3840;
wire  _GEN3849 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3850 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3851 = io_x[4] ? _GEN3850 : _GEN3849;
wire  _GEN3852 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3853 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3854 = io_x[4] ? _GEN3853 : _GEN3852;
wire  _GEN3855 = io_x[12] ? _GEN3854 : _GEN3851;
wire  _GEN3856 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3857 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3858 = io_x[4] ? _GEN3857 : _GEN3856;
wire  _GEN3859 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3860 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3861 = io_x[4] ? _GEN3860 : _GEN3859;
wire  _GEN3862 = io_x[12] ? _GEN3861 : _GEN3858;
wire  _GEN3863 = io_x[0] ? _GEN3862 : _GEN3855;
wire  _GEN3864 = io_x[42] ? _GEN3863 : _GEN3848;
wire  _GEN3865 = io_x[48] ? _GEN3864 : _GEN3833;
wire  _GEN3866 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3867 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3868 = io_x[4] ? _GEN3867 : _GEN3866;
wire  _GEN3869 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3870 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3871 = io_x[4] ? _GEN3870 : _GEN3869;
wire  _GEN3872 = io_x[12] ? _GEN3871 : _GEN3868;
wire  _GEN3873 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3874 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3875 = io_x[4] ? _GEN3874 : _GEN3873;
wire  _GEN3876 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3877 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3878 = io_x[4] ? _GEN3877 : _GEN3876;
wire  _GEN3879 = io_x[12] ? _GEN3878 : _GEN3875;
wire  _GEN3880 = io_x[0] ? _GEN3879 : _GEN3872;
wire  _GEN3881 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3882 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3883 = io_x[4] ? _GEN3882 : _GEN3881;
wire  _GEN3884 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3885 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3886 = io_x[4] ? _GEN3885 : _GEN3884;
wire  _GEN3887 = io_x[12] ? _GEN3886 : _GEN3883;
wire  _GEN3888 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3889 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3890 = io_x[4] ? _GEN3889 : _GEN3888;
wire  _GEN3891 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3892 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3893 = io_x[4] ? _GEN3892 : _GEN3891;
wire  _GEN3894 = io_x[12] ? _GEN3893 : _GEN3890;
wire  _GEN3895 = io_x[0] ? _GEN3894 : _GEN3887;
wire  _GEN3896 = io_x[42] ? _GEN3895 : _GEN3880;
wire  _GEN3897 = 1'b0;
wire  _GEN3898 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3899 = io_x[4] ? _GEN3898 : _GEN3897;
wire  _GEN3900 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3901 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3902 = io_x[4] ? _GEN3901 : _GEN3900;
wire  _GEN3903 = io_x[12] ? _GEN3902 : _GEN3899;
wire  _GEN3904 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3905 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3906 = io_x[4] ? _GEN3905 : _GEN3904;
wire  _GEN3907 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3908 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3909 = io_x[4] ? _GEN3908 : _GEN3907;
wire  _GEN3910 = io_x[12] ? _GEN3909 : _GEN3906;
wire  _GEN3911 = io_x[0] ? _GEN3910 : _GEN3903;
wire  _GEN3912 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3913 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3914 = io_x[4] ? _GEN3913 : _GEN3912;
wire  _GEN3915 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3916 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3917 = io_x[4] ? _GEN3916 : _GEN3915;
wire  _GEN3918 = io_x[12] ? _GEN3917 : _GEN3914;
wire  _GEN3919 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3920 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3921 = io_x[4] ? _GEN3920 : _GEN3919;
wire  _GEN3922 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3923 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3924 = io_x[4] ? _GEN3923 : _GEN3922;
wire  _GEN3925 = io_x[12] ? _GEN3924 : _GEN3921;
wire  _GEN3926 = io_x[0] ? _GEN3925 : _GEN3918;
wire  _GEN3927 = io_x[42] ? _GEN3926 : _GEN3911;
wire  _GEN3928 = io_x[48] ? _GEN3927 : _GEN3896;
wire  _GEN3929 = io_x[2] ? _GEN3928 : _GEN3865;
wire  _GEN3930 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3931 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3932 = io_x[4] ? _GEN3931 : _GEN3930;
wire  _GEN3933 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3934 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3935 = io_x[4] ? _GEN3934 : _GEN3933;
wire  _GEN3936 = io_x[12] ? _GEN3935 : _GEN3932;
wire  _GEN3937 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3938 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3939 = io_x[4] ? _GEN3938 : _GEN3937;
wire  _GEN3940 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3941 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3942 = io_x[4] ? _GEN3941 : _GEN3940;
wire  _GEN3943 = io_x[12] ? _GEN3942 : _GEN3939;
wire  _GEN3944 = io_x[0] ? _GEN3943 : _GEN3936;
wire  _GEN3945 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3946 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3947 = io_x[4] ? _GEN3946 : _GEN3945;
wire  _GEN3948 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3949 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3950 = io_x[4] ? _GEN3949 : _GEN3948;
wire  _GEN3951 = io_x[12] ? _GEN3950 : _GEN3947;
wire  _GEN3952 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3953 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3954 = io_x[4] ? _GEN3953 : _GEN3952;
wire  _GEN3955 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3956 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3957 = io_x[4] ? _GEN3956 : _GEN3955;
wire  _GEN3958 = io_x[12] ? _GEN3957 : _GEN3954;
wire  _GEN3959 = io_x[0] ? _GEN3958 : _GEN3951;
wire  _GEN3960 = io_x[42] ? _GEN3959 : _GEN3944;
wire  _GEN3961 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3962 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3963 = io_x[4] ? _GEN3962 : _GEN3961;
wire  _GEN3964 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3965 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3966 = io_x[4] ? _GEN3965 : _GEN3964;
wire  _GEN3967 = io_x[12] ? _GEN3966 : _GEN3963;
wire  _GEN3968 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3969 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3970 = io_x[4] ? _GEN3969 : _GEN3968;
wire  _GEN3971 = 1'b1;
wire  _GEN3972 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3973 = io_x[4] ? _GEN3972 : _GEN3971;
wire  _GEN3974 = io_x[12] ? _GEN3973 : _GEN3970;
wire  _GEN3975 = io_x[0] ? _GEN3974 : _GEN3967;
wire  _GEN3976 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3977 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3978 = io_x[4] ? _GEN3977 : _GEN3976;
wire  _GEN3979 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3980 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3981 = io_x[4] ? _GEN3980 : _GEN3979;
wire  _GEN3982 = io_x[12] ? _GEN3981 : _GEN3978;
wire  _GEN3983 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3984 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3985 = io_x[4] ? _GEN3984 : _GEN3983;
wire  _GEN3986 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3987 = io_x[4] ? _GEN3897 : _GEN3986;
wire  _GEN3988 = io_x[12] ? _GEN3987 : _GEN3985;
wire  _GEN3989 = io_x[0] ? _GEN3988 : _GEN3982;
wire  _GEN3990 = io_x[42] ? _GEN3989 : _GEN3975;
wire  _GEN3991 = io_x[48] ? _GEN3990 : _GEN3960;
wire  _GEN3992 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3993 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3994 = io_x[4] ? _GEN3993 : _GEN3992;
wire  _GEN3995 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN3996 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN3997 = io_x[4] ? _GEN3996 : _GEN3995;
wire  _GEN3998 = io_x[12] ? _GEN3997 : _GEN3994;
wire  _GEN3999 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4000 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4001 = io_x[4] ? _GEN4000 : _GEN3999;
wire  _GEN4002 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4003 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4004 = io_x[4] ? _GEN4003 : _GEN4002;
wire  _GEN4005 = io_x[12] ? _GEN4004 : _GEN4001;
wire  _GEN4006 = io_x[0] ? _GEN4005 : _GEN3998;
wire  _GEN4007 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4008 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4009 = io_x[4] ? _GEN4008 : _GEN4007;
wire  _GEN4010 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4011 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4012 = io_x[4] ? _GEN4011 : _GEN4010;
wire  _GEN4013 = io_x[12] ? _GEN4012 : _GEN4009;
wire  _GEN4014 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4015 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4016 = io_x[4] ? _GEN4015 : _GEN4014;
wire  _GEN4017 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4018 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4019 = io_x[4] ? _GEN4018 : _GEN4017;
wire  _GEN4020 = io_x[12] ? _GEN4019 : _GEN4016;
wire  _GEN4021 = io_x[0] ? _GEN4020 : _GEN4013;
wire  _GEN4022 = io_x[42] ? _GEN4021 : _GEN4006;
wire  _GEN4023 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4024 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4025 = io_x[4] ? _GEN4024 : _GEN4023;
wire  _GEN4026 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4027 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4028 = io_x[4] ? _GEN4027 : _GEN4026;
wire  _GEN4029 = io_x[12] ? _GEN4028 : _GEN4025;
wire  _GEN4030 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4031 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4032 = io_x[4] ? _GEN4031 : _GEN4030;
wire  _GEN4033 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4034 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4035 = io_x[4] ? _GEN4034 : _GEN4033;
wire  _GEN4036 = io_x[12] ? _GEN4035 : _GEN4032;
wire  _GEN4037 = io_x[0] ? _GEN4036 : _GEN4029;
wire  _GEN4038 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4039 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4040 = io_x[4] ? _GEN4039 : _GEN4038;
wire  _GEN4041 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4042 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4043 = io_x[4] ? _GEN4042 : _GEN4041;
wire  _GEN4044 = io_x[12] ? _GEN4043 : _GEN4040;
wire  _GEN4045 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4046 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4047 = io_x[4] ? _GEN4046 : _GEN4045;
wire  _GEN4048 = io_x[8] ? _GEN3801 : _GEN3802;
wire  _GEN4049 = io_x[8] ? _GEN3802 : _GEN3801;
wire  _GEN4050 = io_x[4] ? _GEN4049 : _GEN4048;
wire  _GEN4051 = io_x[12] ? _GEN4050 : _GEN4047;
wire  _GEN4052 = io_x[0] ? _GEN4051 : _GEN4044;
wire  _GEN4053 = io_x[42] ? _GEN4052 : _GEN4037;
wire  _GEN4054 = io_x[48] ? _GEN4053 : _GEN4022;
wire  _GEN4055 = io_x[2] ? _GEN4054 : _GEN3991;
wire  _GEN4056 = io_x[34] ? _GEN4055 : _GEN3929;
assign io_y[6] = _GEN4056;
wire  _GEN4057 = 1'b0;
wire  _GEN4058 = 1'b1;
wire  _GEN4059 = io_x[41] ? _GEN4058 : _GEN4057;
wire  _GEN4060 = io_x[41] ? _GEN4058 : _GEN4057;
wire  _GEN4061 = io_x[42] ? _GEN4060 : _GEN4059;
wire  _GEN4062 = io_x[41] ? _GEN4058 : _GEN4057;
wire  _GEN4063 = io_x[41] ? _GEN4058 : _GEN4057;
wire  _GEN4064 = io_x[42] ? _GEN4063 : _GEN4062;
wire  _GEN4065 = io_x[15] ? _GEN4064 : _GEN4061;
assign io_y[5] = _GEN4065;
wire  _GEN4066 = 1'b0;
wire  _GEN4067 = 1'b1;
wire  _GEN4068 = io_x[40] ? _GEN4067 : _GEN4066;
wire  _GEN4069 = io_x[40] ? _GEN4067 : _GEN4066;
wire  _GEN4070 = io_x[78] ? _GEN4069 : _GEN4068;
wire  _GEN4071 = io_x[40] ? _GEN4067 : _GEN4066;
wire  _GEN4072 = io_x[40] ? _GEN4067 : _GEN4066;
wire  _GEN4073 = io_x[78] ? _GEN4072 : _GEN4071;
wire  _GEN4074 = io_x[39] ? _GEN4073 : _GEN4070;
assign io_y[4] = _GEN4074;
wire  _GEN4075 = 1'b0;
wire  _GEN4076 = 1'b1;
wire  _GEN4077 = io_x[39] ? _GEN4076 : _GEN4075;
wire  _GEN4078 = io_x[39] ? _GEN4076 : _GEN4075;
wire  _GEN4079 = io_x[72] ? _GEN4078 : _GEN4077;
wire  _GEN4080 = io_x[39] ? _GEN4076 : _GEN4075;
wire  _GEN4081 = io_x[39] ? _GEN4076 : _GEN4075;
wire  _GEN4082 = io_x[72] ? _GEN4081 : _GEN4080;
wire  _GEN4083 = io_x[40] ? _GEN4082 : _GEN4079;
assign io_y[3] = _GEN4083;
wire  _GEN4084 = 1'b0;
wire  _GEN4085 = 1'b1;
wire  _GEN4086 = io_x[38] ? _GEN4085 : _GEN4084;
wire  _GEN4087 = io_x[38] ? _GEN4085 : _GEN4084;
wire  _GEN4088 = io_x[77] ? _GEN4087 : _GEN4086;
wire  _GEN4089 = io_x[38] ? _GEN4085 : _GEN4084;
wire  _GEN4090 = io_x[38] ? _GEN4085 : _GEN4084;
wire  _GEN4091 = io_x[77] ? _GEN4090 : _GEN4089;
wire  _GEN4092 = io_x[43] ? _GEN4091 : _GEN4088;
wire  _GEN4093 = io_x[38] ? _GEN4085 : _GEN4084;
wire  _GEN4094 = io_x[38] ? _GEN4085 : _GEN4084;
wire  _GEN4095 = io_x[77] ? _GEN4094 : _GEN4093;
wire  _GEN4096 = io_x[38] ? _GEN4085 : _GEN4084;
wire  _GEN4097 = io_x[38] ? _GEN4085 : _GEN4084;
wire  _GEN4098 = io_x[77] ? _GEN4097 : _GEN4096;
wire  _GEN4099 = io_x[43] ? _GEN4098 : _GEN4095;
wire  _GEN4100 = io_x[81] ? _GEN4099 : _GEN4092;
assign io_y[2] = _GEN4100;
wire  _GEN4101 = 1'b0;
wire  _GEN4102 = 1'b1;
wire  _GEN4103 = io_x[37] ? _GEN4102 : _GEN4101;
wire  _GEN4104 = io_x[37] ? _GEN4102 : _GEN4101;
wire  _GEN4105 = io_x[41] ? _GEN4104 : _GEN4103;
assign io_y[1] = _GEN4105;
wire  _GEN4106 = 1'b0;
wire  _GEN4107 = 1'b1;
wire  _GEN4108 = io_x[34] ? _GEN4107 : _GEN4106;
wire  _GEN4109 = io_x[34] ? _GEN4107 : _GEN4106;
wire  _GEN4110 = io_x[45] ? _GEN4109 : _GEN4108;
assign io_y[0] = _GEN4110;
endmodule
